library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.fda_package.all;

package content_package is

-- 320x320 - 80fdas
constant c_PIXEL : t_MATRIX := (
0 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
1 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
2 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
3 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
4 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
5 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
6 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
7 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
8 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
9 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
10 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
11 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
12 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
13 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
14 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
15 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
16 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
17 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
18 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
19 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
20 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),21 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),22 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),23 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),24 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),25 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),26 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),27 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),28 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),29 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
30 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),31 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),32 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),33 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),34 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),35 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),36 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),37 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),38 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),39 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
40 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),41 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),42 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),43 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),44 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),45 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),46 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),47 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),48 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),49 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
50 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),51 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),52 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),53 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),54 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),55 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),56 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),57 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),58 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),59 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
60 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),61 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),62 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),63 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),64 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),65 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),66 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),67 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),68 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),69 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),
70 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),71 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),72 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),73 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),74 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),75 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),76 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),77 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),78 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",),79 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00", 1024=>x"8300",
1025=>x"8400", 1026=>x"8100", 1027=>x"8100", 1028=>x"8100",
1029=>x"8200", 1030=>x"8200", 1031=>x"7f00", 1032=>x"8300",
1033=>x"8300", 1034=>x"8200", 1035=>x"7e00", 1036=>x"8600",
1037=>x"8100", 1038=>x"8100", 1039=>x"7f00", 1040=>x"8900",
1041=>x"8000", 1042=>x"8100", 1043=>x"7e00", 1044=>x"8200",
1045=>x"8200", 1046=>x"8100", 1047=>x"8100", 1048=>x"8100",
1049=>x"8200", 1050=>x"8000", 1051=>x"7f00", 1052=>x"7f00",
1053=>x"7f00", 1054=>x"7f00", 1055=>x"7e00", 1056=>x"8100",
1057=>x"7e00", 1058=>x"7f00", 1059=>x"7f00", 1060=>x"7f00",
1061=>x"7d00", 1062=>x"8000", 1063=>x"7f00", 1064=>x"8000",
1065=>x"7d00", 1066=>x"7e00", 1067=>x"7e00", 1068=>x"7f00",
1069=>x"8100", 1070=>x"8000", 1071=>x"8000", 1072=>x"7f00",
1073=>x"8000", 1074=>x"8100", 1075=>x"8000", 1076=>x"7e00",
1077=>x"8100", 1078=>x"7f00", 1079=>x"7f00", 1080=>x"7d00",
1081=>x"8100", 1082=>x"7f00", 1083=>x"7c00", 1084=>x"8300",
1085=>x"8000", 1086=>x"7e00", 1087=>x"7f00", 1088=>x"7f00",
1089=>x"7f00", 1090=>x"7e00", 1091=>x"8000", 1092=>x"7d00",
1093=>x"7d00", 1094=>x"7c00", 1095=>x"7f00", 1096=>x"7c00",
1097=>x"7c00", 1098=>x"7d00", 1099=>x"7d00", 1100=>x"7900",
1101=>x"7a00", 1102=>x"7c00", 1103=>x"7a00", 1104=>x"7500",
1105=>x"7600", 1106=>x"7900", 1107=>x"7800", 1108=>x"7200",
1109=>x"7000", 1110=>x"7700", 1111=>x"7800", 1112=>x"a500",
1113=>x"7c00", 1114=>x"6f00", 1115=>x"7300", 1116=>x"c600",
1117=>x"bb00", 1118=>x"8e00", 1119=>x"9100", 1120=>x"c300",
1121=>x"cb00", 1122=>x"c400", 1123=>x"a200", 1124=>x"c600",
1125=>x"c500", 1126=>x"ca00", 1127=>x"c800", 1128=>x"c500",
1129=>x"c400", 1130=>x"c400", 1131=>x"c200", 1132=>x"c500",
1133=>x"c300", 1134=>x"c400", 1135=>x"c500", 1136=>x"c400",
1137=>x"c300", 1138=>x"c700", 1139=>x"c500", 1140=>x"c300",
1141=>x"c600", 1142=>x"c500", 1143=>x"c400", 1144=>x"c400",
1145=>x"c400", 1146=>x"c400", 1147=>x"c400", 1148=>x"c400",
1149=>x"c400", 1150=>x"c400", 1151=>x"c000", 1152=>x"c300",
1153=>x"c300", 1154=>x"c500", 1155=>x"c000", 1156=>x"c300",
1157=>x"c000", 1158=>x"c000", 1159=>x"bc00", 1160=>x"ba00",
1161=>x"b900", 1162=>x"b900", 1163=>x"b900", 1164=>x"b800",
1165=>x"bc00", 1166=>x"cb00", 1167=>x"d300", 1168=>x"ce00",
1169=>x"d400", 1170=>x"d300", 1171=>x"d500", 1172=>x"d500",
1173=>x"d200", 1174=>x"cd00", 1175=>x"cd00", 1176=>x"d200",
1177=>x"ce00", 1178=>x"c800", 1179=>x"3500", 1180=>x"cb00",
1181=>x"cd00", 1182=>x"d000", 1183=>x"c900", 1184=>x"d500",
1185=>x"d000", 1186=>x"cd00", 1187=>x"cb00", 1188=>x"d000",
1189=>x"d000", 1190=>x"cc00", 1191=>x"c900", 1192=>x"cc00",
1193=>x"c500", 1194=>x"c500", 1195=>x"c400", 1196=>x"c300",
1197=>x"c200", 1198=>x"c300", 1199=>x"c700", 1200=>x"c400",
1201=>x"cb00", 1202=>x"c600", 1203=>x"c200", 1204=>x"ca00",
1205=>x"c000", 1206=>x"c400", 1207=>x"c500", 1208=>x"c400",
1209=>x"c800", 1210=>x"cc00", 1211=>x"cb00", 1212=>x"cc00",
1213=>x"cd00", 1214=>x"ce00", 1215=>x"cc00", 1216=>x"c900",
1217=>x"cd00", 1218=>x"cc00", 1219=>x"ce00", 1220=>x"c500",
1221=>x"c900", 1222=>x"cc00", 1223=>x"cb00", 1224=>x"c700",
1225=>x"c600", 1226=>x"cd00", 1227=>x"ce00", 1228=>x"c300",
1229=>x"cc00", 1230=>x"c700", 1231=>x"3100", 1232=>x"c400",
1233=>x"c600", 1234=>x"c500", 1235=>x"c400", 1236=>x"c400",
1237=>x"c000", 1238=>x"c600", 1239=>x"c600", 1240=>x"c400",
1241=>x"c100", 1242=>x"c000", 1243=>x"c200", 1244=>x"be00",
1245=>x"be00", 1246=>x"bb00", 1247=>x"b700", 1248=>x"ba00",
1249=>x"b100", 1250=>x"c100", 1251=>x"c300", 1252=>x"b400",
1253=>x"c600", 1254=>x"c900", 1255=>x"ca00", 1256=>x"c000",
1257=>x"c400", 1258=>x"c800", 1259=>x"c700", 1260=>x"bc00",
1261=>x"be00", 1262=>x"c500", 1263=>x"c800", 1264=>x"b500",
1265=>x"bc00", 1266=>x"c100", 1267=>x"c300", 1268=>x"b800",
1269=>x"b400", 1270=>x"bc00", 1271=>x"bf00", 1272=>x"c100",
1273=>x"b900", 1274=>x"b800", 1275=>x"c000", 1276=>x"b200",
1277=>x"bd00", 1278=>x"bd00", 1279=>x"b500",)
);



---- 100x100 - 20 FDAs
---- constant c_PIXEL  : t_MATRIX := (
---- 0   => (0=>x"a200", 1=>x"a100", 2=>x"9f00", 3=>x"9d00", 4=>x"9b00", 5=>x"9e00", 6=>x"9f00", 7=>x"9c00", 8=>x"9a00", 9=>x"9a00",
---- 10=>x"9e00", 11=>x"9200", 12=>x"9c00", 13=>x"9c00", 14=>x"9c00", 15=>x"9000", 16=>x"9900", 17=>x"9c00", 18=>x"9c00",
---- 19=>x"9a00", 20=>x"9d00", 21=>x"9c00", 22=>x"9e00", 23=>x"9e00", 24=>x"9a00", 25=>x"9500", 26=>x"9b00", 27=>x"9a00",
---- 28=>x"9e00", 29=>x"9c00", 30=>x"9200", 31=>x"9c00", 32=>x"9700", 33=>x"a100", 34=>x"a300", 35=>x"a300", 36=>x"8300",
---- 37=>x"a600", 38=>x"9100", 39=>x"aa00", 40=>x"a000", 41=>x"a200", 42=>x"a200", 43=>x"ac00", 44=>x"a500", 45=>x"a200",
---- 46=>x"9f00", 47=>x"9a00", 48=>x"a400", 49=>x"8f00", 50=>x"a200", 51=>x"a100", 52=>x"ab00", 53=>x"a600", 54=>x"8900",
---- 55=>x"8400", 56=>x"aa00", 57=>x"a900", 58=>x"9900", 59=>x"7e00", 60=>x"a700", 61=>x"ad00", 62=>x"a000", 63=>x"8100",
---- 64=>x"5e00", 65=>x"ad00", 66=>x"a900", 67=>x"9700", 68=>x"7200", 69=>x"4300", 70=>x"ad00", 71=>x"a200", 72=>x"8600",
---- 73=>x"5400", 74=>x"7500", 75=>x"a000", 76=>x"9200", 77=>x"6900", 78=>x"4f00", 79=>x"4d00", 80=>x"9d00", 81=>x"8700",
---- 82=>x"4f00", 83=>x"5400", 84=>x"5300", 85=>x"8d00", 86=>x"5d00", 87=>x"5100", 88=>x"5700", 89=>x"6000", 90=>x"7200",
---- 91=>x"5100", 92=>x"6500", 93=>x"5700", 94=>x"5300", 95=>x"5700", 96=>x"5600", 97=>x"6000", 98=>x"5a00", 99=>x"5400",
---- 100=>x"5500", 101=>x"5c00", 102=>x"5c00", 103=>x"5a00", 104=>x"5800", 105=>x"5a00", 106=>x"5c00", 107=>x"5b00", 108=>x"5900",
---- 109=>x"5400", 110=>x"5a00", 111=>x"5900", 112=>x"5700", 113=>x"6400", 114=>x"5c00", 115=>x"6100", 116=>x"6000", 117=>x"5700",
---- 118=>x"5b00", 119=>x"5200", 120=>x"5700", 121=>x"5900", 122=>x"6c00", 123=>x"5d00", 124=>x"5500", 125=>x"6d00", 126=>x"5d00",
---- 127=>x"5f00", 128=>x"6e00", 129=>x"5c00", 130=>x"6100", 131=>x"6200", 132=>x"6c00", 133=>x"6400", 134=>x"5b00", 135=>x"6300",
---- 136=>x"6400", 137=>x"6200", 138=>x"6300", 139=>x"6100", 140=>x"6400", 141=>x"6400", 142=>x"6200", 143=>x"6300", 144=>x"6100",
---- 145=>x"6400", 146=>x"6200", 147=>x"6000", 148=>x"6000", 149=>x"6100", 150=>x"5f00", 151=>x"6f00", 152=>x"5e00", 153=>x"6f00",
---- 154=>x"5d00", 155=>x"6000", 156=>x"5d00", 157=>x"6900", 158=>x"5d00", 159=>x"5f00", 160=>x"6000", 161=>x"6400", 162=>x"5e00",
---- 163=>x"5d00", 164=>x"6000", 165=>x"5e00", 166=>x"6800", 167=>x"5e00", 168=>x"6100", 169=>x"6600", 170=>x"6900", 171=>x"6500",
---- 172=>x"6100", 173=>x"6200", 174=>x"6e00", 175=>x"6000", 176=>x"7200", 177=>x"6100", 178=>x"6400", 179=>x"6a00", 180=>x"6400",
---- 181=>x"6500", 182=>x"6000", 183=>x"6200", 184=>x"6b00", 185=>x"6800", 186=>x"7100", 187=>x"6f00", 188=>x"6300", 189=>x"7000",
---- 190=>x"6b00", 191=>x"6700", 192=>x"6d00", 193=>x"6200", 194=>x"6500", 195=>x"6a00", 196=>x"6a00", 197=>x"6500", 198=>x"6200",
---- 199=>x"6200", 200=>x"6b00", 201=>x"6a00", 202=>x"6e00", 203=>x"6500", 204=>x"6800", 205=>x"6b00", 206=>x"6900", 207=>x"7100",
---- 208=>x"6300", 209=>x"5800", 210=>x"7100", 211=>x"6800", 212=>x"6700", 213=>x"6200", 214=>x"5600", 215=>x"6600", 216=>x"6900",
---- 217=>x"6500", 218=>x"6400", 219=>x"5a00", 220=>x"6700", 221=>x"6600", 222=>x"6700", 223=>x"6200", 224=>x"5a00", 225=>x"6800",
---- 226=>x"7000", 227=>x"6100", 228=>x"6000", 229=>x"5800", 230=>x"6600", 231=>x"6800", 232=>x"6200", 233=>x"6100", 234=>x"5800",
---- 235=>x"6500", 236=>x"6400", 237=>x"6000", 238=>x"6000", 239=>x"5800", 240=>x"6600", 241=>x"6400", 242=>x"6d00", 243=>x"6700",
---- 244=>x"5900", 245=>x"7500", 246=>x"6500", 247=>x"6500", 248=>x"6d00", 249=>x"6100", 250=>x"6200", 251=>x"6600", 252=>x"6300",
---- 253=>x"6100", 254=>x"5200", 255=>x"5f00", 256=>x"5e00", 257=>x"5c00", 258=>x"5a00", 259=>x"4c00", 260=>x"6400", 261=>x"5f00",
---- 262=>x"6800", 263=>x"5800", 264=>x"4800", 265=>x"6300", 266=>x"6100", 267=>x"6400", 268=>x"5800", 269=>x"4800", 270=>x"6700",
---- 271=>x"6700", 272=>x"5e00", 273=>x"6600", 274=>x"4700", 275=>x"6400", 276=>x"6300", 277=>x"5800", 278=>x"5600", 279=>x"4100",
---- 280=>x"5c00", 281=>x"7500", 282=>x"4f00", 283=>x"4f00", 284=>x"3b00", 285=>x"5700", 286=>x"5600", 287=>x"6200", 288=>x"4a00",
---- 289=>x"3a00", 290=>x"5100", 291=>x"4b00", 292=>x"4800", 293=>x"4700", 294=>x"3800", 295=>x"4b00", 296=>x"4800", 297=>x"5a00",
---- 298=>x"5000", 299=>x"4a00", 300=>x"4e00", 301=>x"4c00", 302=>x"4a00", 303=>x"4000", 304=>x"3000", 305=>x"5000", 306=>x"4c00",
---- 307=>x"4a00", 308=>x"4000", 309=>x"2b00", 310=>x"5600", 311=>x"5000", 312=>x"4a00", 313=>x"4100", 314=>x"2700", 315=>x"5100",
---- 316=>x"4e00", 317=>x"4e00", 318=>x"4100", 319=>x"5600", 320=>x"4d00", 321=>x"4b00", 322=>x"4c00", 323=>x"4200", 324=>x"4400",
---- 325=>x"5a00", 326=>x"5300", 327=>x"4d00", 328=>x"4300", 329=>x"4300", 330=>x"4600", 331=>x"5300", 332=>x"4400", 333=>x"3d00",
---- 334=>x"4300", 335=>x"4100", 336=>x"4a00", 337=>x"4400", 338=>x"3f00", 339=>x"4400", 340=>x"4700", 341=>x"4500", 342=>x"3f00",
---- 343=>x"3b00", 344=>x"5c00", 345=>x"3600", 346=>x"3800", 347=>x"4000", 348=>x"3b00", 349=>x"4d00", 350=>x"3700", 351=>x"3700",
---- 352=>x"3b00", 353=>x"3400", 354=>x"6500", 355=>x"3400", 356=>x"3200", 357=>x"3500", 358=>x"3300", 359=>x"5700", 360=>x"3000",
---- 361=>x"3200", 362=>x"2d00", 363=>x"3a00", 364=>x"6900", 365=>x"5000", 366=>x"2d00", 367=>x"2e00", 368=>x"4300", 369=>x"6900",
---- 370=>x"2e00", 371=>x"3100", 372=>x"2c00", 373=>x"3c00", 374=>x"5c00", 375=>x"2700", 376=>x"2e00", 377=>x"2700", 378=>x"2e00",
---- 379=>x"6300", 380=>x"5000", 381=>x"3300", 382=>x"4700", 383=>x"2700", 384=>x"4a00", 385=>x"5500", 386=>x"4000", 387=>x"3f00",
---- 388=>x"2d00", 389=>x"3d00", 390=>x"8800", 391=>x"7600", 392=>x"5700", 393=>x"4300", 394=>x"3600", 395=>x"8700", 396=>x"9200",
---- 397=>x"8100", 398=>x"6500", 399=>x"4e00", 400=>x"8000", 401=>x"9400", 402=>x"9800", 403=>x"8400", 404=>x"4f00", 405=>x"4b00",
---- 406=>x"8300", 407=>x"9f00", 408=>x"a000", 409=>x"6900", 410=>x"1f00", 411=>x"6800", 412=>x"a700", 413=>x"a900", 414=>x"7f00",
---- 415=>x"1e00", 416=>x"4400", 417=>x"a800", 418=>x"af00", 419=>x"8400", 420=>x"1800", 421=>x"7700", 422=>x"9b00", 423=>x"b000",
---- 424=>x"7f00", 425=>x"1a00", 426=>x"3b00", 427=>x"9a00", 428=>x"b100", 429=>x"9400", 430=>x"1c00", 431=>x"2900", 432=>x"9a00",
---- 433=>x"9e00", 434=>x"9100", 435=>x"1a00", 436=>x"4900", 437=>x"8c00", 438=>x"b300", 439=>x"9900", 440=>x"2300", 441=>x"1e00",
---- 442=>x"8200", 443=>x"af00", 444=>x"9a00", 445=>x"2700", 446=>x"1e00", 447=>x"7300", 448=>x"aa00", 449=>x"9c00", 450=>x"2300",
---- 451=>x"1d00", 452=>x"6a00", 453=>x"ac00", 454=>x"a500", 455=>x"2100", 456=>x"1800", 457=>x"6100", 458=>x"b500", 459=>x"9800",
---- 460=>x"2e00", 461=>x"3000", 462=>x"5f00", 463=>x"b300", 464=>x"b800", 465=>x"5b00", 466=>x"5500", 467=>x"6a00", 468=>x"ad00",
---- 469=>x"bb00", 470=>x"5400", 471=>x"6500", 472=>x"7e00", 473=>x"ae00", 474=>x"b800", 475=>x"3d00", 476=>x"7600", 477=>x"6e00",
---- 478=>x"a400", 479=>x"b600", 480=>x"2e00", 481=>x"4a00", 482=>x"6500", 483=>x"9c00", 484=>x"b200", 485=>x"3400", 486=>x"5b00",
---- 487=>x"5400", 488=>x"9700", 489=>x"c300", 490=>x"3300", 491=>x"3100", 492=>x"3800", 493=>x"b100", 494=>x"d600", 495=>x"2f00",
---- 496=>x"3100", 497=>x"5000", 498=>x"af00", 499=>x"af00"),
---- 1   => (0=>x"9900", 1=>x"9b00", 2=>x"9400", 3=>x"ac00", 4=>x"9a00", 5=>x"9a00", 6=>x"9a00", 7=>x"a200", 8=>x"aa00", 9=>x"ae00",
---- 10=>x"8900", 11=>x"9500", 12=>x"a700", 13=>x"a900", 14=>x"a900", 15=>x"9b00", 16=>x"a400", 17=>x"a800", 18=>x"a600",
---- 19=>x"a500", 20=>x"9c00", 21=>x"a600", 22=>x"a000", 23=>x"9f00", 24=>x"a100", 25=>x"a300", 26=>x"a900", 27=>x"9200",
---- 28=>x"9e00", 29=>x"9f00", 30=>x"a900", 31=>x"a900", 32=>x"a600", 33=>x"9e00", 34=>x"a100", 35=>x"a000", 36=>x"a600",
---- 37=>x"a000", 38=>x"9f00", 39=>x"9200", 40=>x"9700", 41=>x"9f00", 42=>x"a000", 43=>x"a000", 44=>x"9300", 45=>x"9200",
---- 46=>x"9000", 47=>x"a300", 48=>x"a100", 49=>x"9c00", 50=>x"8500", 51=>x"8d00", 52=>x"a500", 53=>x"a200", 54=>x"9600",
---- 55=>x"7a00", 56=>x"9700", 57=>x"a600", 58=>x"a400", 59=>x"a600", 60=>x"7700", 61=>x"9900", 62=>x"a700", 63=>x"a500",
---- 64=>x"a500", 65=>x"7900", 66=>x"9a00", 67=>x"a800", 68=>x"a700", 69=>x"a400", 70=>x"7700", 71=>x"8b00", 72=>x"aa00",
---- 73=>x"9500", 74=>x"a500", 75=>x"7c00", 76=>x"9a00", 77=>x"a700", 78=>x"ab00", 79=>x"a500", 80=>x"7a00", 81=>x"9800",
---- 82=>x"a900", 83=>x"9500", 84=>x"a800", 85=>x"8000", 86=>x"9300", 87=>x"a600", 88=>x"a700", 89=>x"a700", 90=>x"7800",
---- 91=>x"9700", 92=>x"a400", 93=>x"a700", 94=>x"a500", 95=>x"7600", 96=>x"9400", 97=>x"a400", 98=>x"a600", 99=>x"a500",
---- 100=>x"7800", 101=>x"9500", 102=>x"a300", 103=>x"a500", 104=>x"a600", 105=>x"7700", 106=>x"9600", 107=>x"a200", 108=>x"a400",
---- 109=>x"a300", 110=>x"7600", 111=>x"9500", 112=>x"a300", 113=>x"a400", 114=>x"a300", 115=>x"7400", 116=>x"9400", 117=>x"a300",
---- 118=>x"a400", 119=>x"a300", 120=>x"7200", 121=>x"8800", 122=>x"a700", 123=>x"a700", 124=>x"a500", 125=>x"7400", 126=>x"9500",
---- 127=>x"9500", 128=>x"aa00", 129=>x"a700", 130=>x"7300", 131=>x"9400", 132=>x"a400", 133=>x"a600", 134=>x"a800", 135=>x"7800",
---- 136=>x"9400", 137=>x"a200", 138=>x"ab00", 139=>x"ac00", 140=>x"7800", 141=>x"9600", 142=>x"a800", 143=>x"9700", 144=>x"af00",
---- 145=>x"7500", 146=>x"8e00", 147=>x"a900", 148=>x"af00", 149=>x"b000", 150=>x"7400", 151=>x"9000", 152=>x"a900", 153=>x"af00",
---- 154=>x"9800", 155=>x"7800", 156=>x"9100", 157=>x"aa00", 158=>x"ab00", 159=>x"ad00", 160=>x"7a00", 161=>x"9400", 162=>x"9500",
---- 163=>x"ac00", 164=>x"ac00", 165=>x"7b00", 166=>x"9100", 167=>x"aa00", 168=>x"ac00", 169=>x"ac00", 170=>x"7d00", 171=>x"9800",
---- 172=>x"aa00", 173=>x"ad00", 174=>x"ae00", 175=>x"7e00", 176=>x"9900", 177=>x"ab00", 178=>x"ac00", 179=>x"ae00", 180=>x"7f00",
---- 181=>x"9800", 182=>x"ab00", 183=>x"ab00", 184=>x"ad00", 185=>x"7d00", 186=>x"9700", 187=>x"a900", 188=>x"a600", 189=>x"ab00",
---- 190=>x"7c00", 191=>x"9700", 192=>x"aa00", 193=>x"9f00", 194=>x"ad00", 195=>x"7800", 196=>x"9700", 197=>x"ac00", 198=>x"9800",
---- 199=>x"ad00", 200=>x"7600", 201=>x"9500", 202=>x"ab00", 203=>x"ae00", 204=>x"af00", 205=>x"7100", 206=>x"9800", 207=>x"9500",
---- 208=>x"b000", 209=>x"ae00", 210=>x"7000", 211=>x"8a00", 212=>x"ad00", 213=>x"9800", 214=>x"b000", 215=>x"6f00", 216=>x"9400",
---- 217=>x"a900", 218=>x"a200", 219=>x"af00", 220=>x"6d00", 221=>x"9500", 222=>x"a800", 223=>x"a700", 224=>x"ad00", 225=>x"7000",
---- 226=>x"9000", 227=>x"aa00", 228=>x"b000", 229=>x"9400", 230=>x"6e00", 231=>x"9300", 232=>x"9700", 233=>x"b200", 234=>x"9b00",
---- 235=>x"6b00", 236=>x"9600", 237=>x"9d00", 238=>x"af00", 239=>x"b100", 240=>x"6900", 241=>x"9600", 242=>x"9800", 243=>x"b100",
---- 244=>x"b100", 245=>x"6700", 246=>x"9200", 247=>x"aa00", 248=>x"ae00", 249=>x"b000", 250=>x"6700", 251=>x"9200", 252=>x"a900",
---- 253=>x"b100", 254=>x"b200", 255=>x"5f00", 256=>x"9000", 257=>x"aa00", 258=>x"af00", 259=>x"b300", 260=>x"7000", 261=>x"9000",
---- 262=>x"ab00", 263=>x"b200", 264=>x"a300", 265=>x"5a00", 266=>x"9100", 267=>x"aa00", 268=>x"b400", 269=>x"af00", 270=>x"5900",
---- 271=>x"8a00", 272=>x"aa00", 273=>x"b400", 274=>x"b800", 275=>x"5100", 276=>x"9000", 277=>x"ab00", 278=>x"9c00", 279=>x"b800",
---- 280=>x"4e00", 281=>x"8e00", 282=>x"a800", 283=>x"b500", 284=>x"b600", 285=>x"4f00", 286=>x"8d00", 287=>x"ab00", 288=>x"b200",
---- 289=>x"b700", 290=>x"4c00", 291=>x"8f00", 292=>x"9900", 293=>x"b300", 294=>x"9d00", 295=>x"4700", 296=>x"8e00", 297=>x"a700",
---- 298=>x"ae00", 299=>x"b000", 300=>x"4800", 301=>x"8d00", 302=>x"a500", 303=>x"ae00", 304=>x"ab00", 305=>x"3d00", 306=>x"8c00",
---- 307=>x"a600", 308=>x"af00", 309=>x"a000", 310=>x"6700", 311=>x"8400", 312=>x"a800", 313=>x"af00", 314=>x"9d00", 315=>x"5900",
---- 316=>x"8600", 317=>x"a700", 318=>x"af00", 319=>x"9b00", 320=>x"6900", 321=>x"9700", 322=>x"a600", 323=>x"aa00", 324=>x"af00",
---- 325=>x"7300", 326=>x"9900", 327=>x"a500", 328=>x"aa00", 329=>x"b000", 330=>x"7200", 331=>x"9800", 332=>x"a700", 333=>x"9f00",
---- 334=>x"b000", 335=>x"6c00", 336=>x"9700", 337=>x"a700", 338=>x"a200", 339=>x"b100", 340=>x"6b00", 341=>x"9a00", 342=>x"aa00",
---- 343=>x"b000", 344=>x"b300", 345=>x"7300", 346=>x"9900", 347=>x"aa00", 348=>x"b100", 349=>x"b300", 350=>x"6a00", 351=>x"9800",
---- 352=>x"a700", 353=>x"b100", 354=>x"b500", 355=>x"6400", 356=>x"9100", 357=>x"a600", 358=>x"b300", 359=>x"b300", 360=>x"6f00",
---- 361=>x"8b00", 362=>x"a300", 363=>x"b100", 364=>x"b300", 365=>x"6f00", 366=>x"8c00", 367=>x"a400", 368=>x"b200", 369=>x"9900",
---- 370=>x"7600", 371=>x"8d00", 372=>x"a500", 373=>x"ae00", 374=>x"b200", 375=>x"6c00", 376=>x"9000", 377=>x"a600", 378=>x"ad00",
---- 379=>x"b100", 380=>x"6800", 381=>x"8d00", 382=>x"a500", 383=>x"ad00", 384=>x"ad00", 385=>x"5100", 386=>x"7f00", 387=>x"a400",
---- 388=>x"ac00", 389=>x"a900", 390=>x"5600", 391=>x"6f00", 392=>x"a300", 393=>x"a800", 394=>x"ab00", 395=>x"2900", 396=>x"7500",
---- 397=>x"9f00", 398=>x"9500", 399=>x"ac00", 400=>x"2c00", 401=>x"7400", 402=>x"9800", 403=>x"b100", 404=>x"ad00", 405=>x"2900",
---- 406=>x"7400", 407=>x"a800", 408=>x"b200", 409=>x"b000", 410=>x"2300", 411=>x"7200", 412=>x"a700", 413=>x"b100", 414=>x"b100",
---- 415=>x"1a00", 416=>x"7000", 417=>x"a500", 418=>x"b500", 419=>x"af00", 420=>x"1800", 421=>x"6d00", 422=>x"a800", 423=>x"b200",
---- 424=>x"b300", 425=>x"1b00", 426=>x"6800", 427=>x"a800", 428=>x"b600", 429=>x"a400", 430=>x"2200", 431=>x"6200", 432=>x"a900",
---- 433=>x"b300", 434=>x"ad00", 435=>x"2400", 436=>x"7000", 437=>x"a800", 438=>x"9b00", 439=>x"b300", 440=>x"3100", 441=>x"5f00",
---- 442=>x"a400", 443=>x"b400", 444=>x"b100", 445=>x"4300", 446=>x"5c00", 447=>x"a300", 448=>x"b100", 449=>x"af00", 450=>x"4200",
---- 451=>x"5a00", 452=>x"a000", 453=>x"ae00", 454=>x"b000", 455=>x"7500", 456=>x"5100", 457=>x"9d00", 458=>x"ac00", 459=>x"b000",
---- 460=>x"5e00", 461=>x"5300", 462=>x"9e00", 463=>x"ae00", 464=>x"ae00", 465=>x"7200", 466=>x"5900", 467=>x"9b00", 468=>x"b000",
---- 469=>x"b000", 470=>x"8100", 471=>x"5600", 472=>x"9900", 473=>x"ae00", 474=>x"b200", 475=>x"8100", 476=>x"5800", 477=>x"9800",
---- 478=>x"ae00", 479=>x"b100", 480=>x"8d00", 481=>x"6300", 482=>x"9200", 483=>x"b000", 484=>x"b700", 485=>x"9f00", 486=>x"6200",
---- 487=>x"9500", 488=>x"9800", 489=>x"b600", 490=>x"ac00", 491=>x"7000", 492=>x"9100", 493=>x"b100", 494=>x"b300", 495=>x"ad00",
---- 496=>x"7400", 497=>x"9200", 498=>x"ae00", 499=>x"b300"),
---- 2   => (0=>x"a900", 1=>x"9300", 2=>x"6800", 3=>x"5c00", 4=>x"6c00", 5=>x"a500", 6=>x"8c00", 7=>x"6800", 8=>x"5700", 9=>x"6600",
---- 10=>x"a200", 11=>x"8800", 12=>x"6600", 13=>x"5700", 14=>x"5e00", 15=>x"9d00", 16=>x"8900", 17=>x"6700", 18=>x"5800",
---- 19=>x"6500", 20=>x"9e00", 21=>x"8c00", 22=>x"6d00", 23=>x"6000", 24=>x"5f00", 25=>x"a000", 26=>x"8a00", 27=>x"6300",
---- 28=>x"5100", 29=>x"5f00", 30=>x"a200", 31=>x"8c00", 32=>x"6500", 33=>x"5700", 34=>x"6000", 35=>x"a000", 36=>x"8900",
---- 37=>x"6300", 38=>x"5100", 39=>x"6000", 40=>x"a000", 41=>x"8a00", 42=>x"6000", 43=>x"5200", 44=>x"6000", 45=>x"9a00",
---- 46=>x"8d00", 47=>x"6400", 48=>x"5100", 49=>x"5e00", 50=>x"a300", 51=>x"8c00", 52=>x"6000", 53=>x"6700", 54=>x"5b00",
---- 55=>x"a000", 56=>x"8400", 57=>x"6c00", 58=>x"4800", 59=>x"6100", 60=>x"a200", 61=>x"8e00", 62=>x"6500", 63=>x"4a00",
---- 64=>x"5500", 65=>x"a000", 66=>x"8900", 67=>x"6000", 68=>x"4700", 69=>x"5600", 70=>x"9f00", 71=>x"8a00", 72=>x"5d00",
---- 73=>x"4600", 74=>x"5700", 75=>x"9100", 76=>x"8c00", 77=>x"5d00", 78=>x"4900", 79=>x"5700", 80=>x"9e00", 81=>x"8600",
---- 82=>x"5e00", 83=>x"4a00", 84=>x"5900", 85=>x"9d00", 86=>x"8600", 87=>x"5f00", 88=>x"4900", 89=>x"5900", 90=>x"9f00",
---- 91=>x"8500", 92=>x"7000", 93=>x"4800", 94=>x"5c00", 95=>x"9f00", 96=>x"8600", 97=>x"5e00", 98=>x"4b00", 99=>x"5800",
---- 100=>x"9200", 101=>x"8a00", 102=>x"5e00", 103=>x"5c00", 104=>x"5600", 105=>x"a100", 106=>x"8100", 107=>x"7200", 108=>x"4700",
---- 109=>x"5600", 110=>x"a100", 111=>x"8900", 112=>x"6200", 113=>x"4800", 114=>x"5700", 115=>x"a000", 116=>x"8700", 117=>x"5c00",
---- 118=>x"4300", 119=>x"5200", 120=>x"9f00", 121=>x"8800", 122=>x"5b00", 123=>x"4600", 124=>x"4f00", 125=>x"a200", 126=>x"8b00",
---- 127=>x"5f00", 128=>x"4900", 129=>x"5400", 130=>x"a500", 131=>x"8c00", 132=>x"6000", 133=>x"4a00", 134=>x"5600", 135=>x"a800",
---- 136=>x"8600", 137=>x"7000", 138=>x"4800", 139=>x"5900", 140=>x"ab00", 141=>x"8d00", 142=>x"6000", 143=>x"4800", 144=>x"6000",
---- 145=>x"aa00", 146=>x"8e00", 147=>x"6200", 148=>x"4800", 149=>x"5500", 150=>x"ab00", 151=>x"9000", 152=>x"6200", 153=>x"4900",
---- 154=>x"6c00", 155=>x"a700", 156=>x"9100", 157=>x"6000", 158=>x"4900", 159=>x"5700", 160=>x"aa00", 161=>x"9200", 162=>x"6400",
---- 163=>x"4b00", 164=>x"5900", 165=>x"a800", 166=>x"9500", 167=>x"6300", 168=>x"4600", 169=>x"5d00", 170=>x"aa00", 171=>x"9500",
---- 172=>x"6100", 173=>x"4500", 174=>x"5500", 175=>x"ab00", 176=>x"9500", 177=>x"6300", 178=>x"4600", 179=>x"5500", 180=>x"ab00",
---- 181=>x"9600", 182=>x"6100", 183=>x"4800", 184=>x"5600", 185=>x"aa00", 186=>x"9700", 187=>x"6300", 188=>x"4600", 189=>x"5600",
---- 190=>x"aa00", 191=>x"9500", 192=>x"7600", 193=>x"4000", 194=>x"9600", 195=>x"ac00", 196=>x"9000", 197=>x"6900", 198=>x"4200",
---- 199=>x"5600", 200=>x"ad00", 201=>x"8400", 202=>x"6600", 203=>x"4500", 204=>x"5300", 205=>x"ac00", 206=>x"9a00", 207=>x"6700",
---- 208=>x"4100", 209=>x"5200", 210=>x"ad00", 211=>x"9900", 212=>x"6700", 213=>x"4300", 214=>x"5500", 215=>x"ac00", 216=>x"9300",
---- 217=>x"6a00", 218=>x"4500", 219=>x"5300", 220=>x"af00", 221=>x"9500", 222=>x"6d00", 223=>x"4600", 224=>x"5200", 225=>x"a800",
---- 226=>x"9900", 227=>x"6c00", 228=>x"4a00", 229=>x"5900", 230=>x"af00", 231=>x"9a00", 232=>x"6900", 233=>x"4800", 234=>x"5700",
---- 235=>x"af00", 236=>x"9a00", 237=>x"6a00", 238=>x"4800", 239=>x"5500", 240=>x"b000", 241=>x"8e00", 242=>x"6a00", 243=>x"4800",
---- 244=>x"5500", 245=>x"b200", 246=>x"9c00", 247=>x"6b00", 248=>x"4a00", 249=>x"5900", 250=>x"ae00", 251=>x"9d00", 252=>x"6d00",
---- 253=>x"4700", 254=>x"5200", 255=>x"af00", 256=>x"9900", 257=>x"6c00", 258=>x"4300", 259=>x"5300", 260=>x"b700", 261=>x"9900",
---- 262=>x"6d00", 263=>x"4700", 264=>x"5900", 265=>x"9e00", 266=>x"9c00", 267=>x"6f00", 268=>x"4d00", 269=>x"5c00", 270=>x"b800",
---- 271=>x"9f00", 272=>x"7600", 273=>x"5b00", 274=>x"5e00", 275=>x"b700", 276=>x"9f00", 277=>x"7100", 278=>x"5a00", 279=>x"5e00",
---- 280=>x"b500", 281=>x"a000", 282=>x"7100", 283=>x"4b00", 284=>x"5c00", 285=>x"b500", 286=>x"9e00", 287=>x"7600", 288=>x"4a00",
---- 289=>x"5800", 290=>x"b400", 291=>x"9e00", 292=>x"7700", 293=>x"4a00", 294=>x"5a00", 295=>x"b000", 296=>x"9c00", 297=>x"7d00",
---- 298=>x"4400", 299=>x"6900", 300=>x"b000", 301=>x"9c00", 302=>x"7000", 303=>x"3e00", 304=>x"8500", 305=>x"b400", 306=>x"a000",
---- 307=>x"7200", 308=>x"4200", 309=>x"5200", 310=>x"b500", 311=>x"9f00", 312=>x"7300", 313=>x"5600", 314=>x"7b00", 315=>x"b500",
---- 316=>x"9f00", 317=>x"7900", 318=>x"4900", 319=>x"5300", 320=>x"b400", 321=>x"a100", 322=>x"7600", 323=>x"4700", 324=>x"5900",
---- 325=>x"b400", 326=>x"a300", 327=>x"7900", 328=>x"4800", 329=>x"5300", 330=>x"b500", 331=>x"9c00", 332=>x"7900", 333=>x"4100",
---- 334=>x"7900", 335=>x"b700", 336=>x"9f00", 337=>x"7a00", 338=>x"4000", 339=>x"6200", 340=>x"a600", 341=>x"a700", 342=>x"7300",
---- 343=>x"4b00", 344=>x"7b00", 345=>x"b200", 346=>x"9200", 347=>x"7900", 348=>x"8400", 349=>x"4700", 350=>x"a300", 351=>x"ad00",
---- 352=>x"8800", 353=>x"3d00", 354=>x"5b00", 355=>x"b200", 356=>x"a000", 357=>x"7700", 358=>x"4800", 359=>x"8000", 360=>x"b500",
---- 361=>x"9f00", 362=>x"7700", 363=>x"3b00", 364=>x"7400", 365=>x"b500", 366=>x"a300", 367=>x"7500", 368=>x"4000", 369=>x"5e00",
---- 370=>x"b600", 371=>x"a600", 372=>x"7800", 373=>x"3b00", 374=>x"5b00", 375=>x"9c00", 376=>x"a500", 377=>x"6d00", 378=>x"4400",
---- 379=>x"8e00", 380=>x"b200", 381=>x"9a00", 382=>x"7a00", 383=>x"af00", 384=>x"4600", 385=>x"ae00", 386=>x"a900", 387=>x"a200",
---- 388=>x"3300", 389=>x"6100", 390=>x"b300", 391=>x"ac00", 392=>x"6d00", 393=>x"6000", 394=>x"8600", 395=>x"af00", 396=>x"a000",
---- 397=>x"7500", 398=>x"8d00", 399=>x"4300", 400=>x"aa00", 401=>x"9900", 402=>x"be00", 403=>x"8100", 404=>x"2f00", 405=>x"a600",
---- 406=>x"9e00", 407=>x"a600", 408=>x"5a00", 409=>x"2300", 410=>x"b400", 411=>x"a000", 412=>x"9500", 413=>x"7400", 414=>x"2100",
---- 415=>x"b400", 416=>x"a700", 417=>x"7d00", 418=>x"7900", 419=>x"2500", 420=>x"b700", 421=>x"a600", 422=>x"9800", 423=>x"5300",
---- 424=>x"2a00", 425=>x"ae00", 426=>x"a800", 427=>x"8e00", 428=>x"3800", 429=>x"3a00", 430=>x"af00", 431=>x"a300", 432=>x"8b00",
---- 433=>x"5200", 434=>x"2c00", 435=>x"b400", 436=>x"a600", 437=>x"9300", 438=>x"4400", 439=>x"2d00", 440=>x"b300", 441=>x"a400",
---- 442=>x"9b00", 443=>x"4a00", 444=>x"3000", 445=>x"b300", 446=>x"a600", 447=>x"9800", 448=>x"5e00", 449=>x"3200", 450=>x"b500",
---- 451=>x"9800", 452=>x"8b00", 453=>x"5a00", 454=>x"4500", 455=>x"b300", 456=>x"ac00", 457=>x"7b00", 458=>x"6100", 459=>x"3b00",
---- 460=>x"b400", 461=>x"b100", 462=>x"6c00", 463=>x"6100", 464=>x"3000", 465=>x"b700", 466=>x"af00", 467=>x"6f00", 468=>x"6b00",
---- 469=>x"2600", 470=>x"b800", 471=>x"b100", 472=>x"6b00", 473=>x"6000", 474=>x"2a00", 475=>x"ba00", 476=>x"b400", 477=>x"6800",
---- 478=>x"5200", 479=>x"2500", 480=>x"9d00", 481=>x"9e00", 482=>x"6b00", 483=>x"5400", 484=>x"2e00", 485=>x"be00", 486=>x"aa00",
---- 487=>x"4d00", 488=>x"3800", 489=>x"2e00", 490=>x"b700", 491=>x"ac00", 492=>x"6100", 493=>x"2c00", 494=>x"3500", 495=>x"b700",
---- 496=>x"a800", 497=>x"4e00", 498=>x"2f00", 499=>x"2d00"),
---- 3   => (0=>x"6a00", 1=>x"6900", 2=>x"6b00", 3=>x"6d00", 4=>x"6a00", 5=>x"7300", 6=>x"6600", 7=>x"6800", 8=>x"6800", 9=>x"6900",
---- 10=>x"6f00", 11=>x"6900", 12=>x"6900", 13=>x"6600", 14=>x"6400", 15=>x"6a00", 16=>x"6900", 17=>x"7300", 18=>x"6700",
---- 19=>x"6400", 20=>x"6900", 21=>x"6700", 22=>x"7000", 23=>x"6400", 24=>x"6600", 25=>x"6700", 26=>x"6900", 27=>x"6800",
---- 28=>x"6600", 29=>x"6600", 30=>x"6600", 31=>x"6c00", 32=>x"6a00", 33=>x"6500", 34=>x"6500", 35=>x"6700", 36=>x"6400",
---- 37=>x"6600", 38=>x"6400", 39=>x"6700", 40=>x"6600", 41=>x"7200", 42=>x"6500", 43=>x"7200", 44=>x"6400", 45=>x"6500",
---- 46=>x"6900", 47=>x"6600", 48=>x"6500", 49=>x"6500", 50=>x"6300", 51=>x"6700", 52=>x"6700", 53=>x"6600", 54=>x"6800",
---- 55=>x"6800", 56=>x"6800", 57=>x"6800", 58=>x"6c00", 59=>x"6900", 60=>x"5d00", 61=>x"6100", 62=>x"6200", 63=>x"6900",
---- 64=>x"6900", 65=>x"5e00", 66=>x"6300", 67=>x"6300", 68=>x"6100", 69=>x"6500", 70=>x"6000", 71=>x"6200", 72=>x"6300",
---- 73=>x"7b00", 74=>x"5f00", 75=>x"6300", 76=>x"5f00", 77=>x"6f00", 78=>x"5f00", 79=>x"7100", 80=>x"5f00", 81=>x"6400",
---- 82=>x"6100", 83=>x"6500", 84=>x"6300", 85=>x"5e00", 86=>x"6200", 87=>x"6600", 88=>x"6700", 89=>x"6200", 90=>x"6300",
---- 91=>x"6000", 92=>x"6000", 93=>x"7e00", 94=>x"6100", 95=>x"6100", 96=>x"6400", 97=>x"6200", 98=>x"6000", 99=>x"6400",
---- 100=>x"6000", 101=>x"6000", 102=>x"6600", 103=>x"6100", 104=>x"6300", 105=>x"5d00", 106=>x"6300", 107=>x"6300", 108=>x"6c00",
---- 109=>x"6700", 110=>x"5c00", 111=>x"5f00", 112=>x"6200", 113=>x"6200", 114=>x"6400", 115=>x"5b00", 116=>x"6000", 117=>x"6100",
---- 118=>x"5f00", 119=>x"6100", 120=>x"5d00", 121=>x"6300", 122=>x"6300", 123=>x"6300", 124=>x"6300", 125=>x"6e00", 126=>x"6200",
---- 127=>x"6400", 128=>x"6600", 129=>x"6500", 130=>x"6000", 131=>x"6400", 132=>x"6600", 133=>x"6800", 134=>x"6100", 135=>x"5f00",
---- 136=>x"6200", 137=>x"6600", 138=>x"6400", 139=>x"6300", 140=>x"6600", 141=>x"6300", 142=>x"6300", 143=>x"6200", 144=>x"6200",
---- 145=>x"5d00", 146=>x"6100", 147=>x"6100", 148=>x"6200", 149=>x"6100", 150=>x"6000", 151=>x"6a00", 152=>x"7600", 153=>x"6100",
---- 154=>x"6100", 155=>x"6800", 156=>x"6300", 157=>x"6000", 158=>x"6200", 159=>x"6000", 160=>x"5f00", 161=>x"6100", 162=>x"6100",
---- 163=>x"6100", 164=>x"6800", 165=>x"6900", 166=>x"6100", 167=>x"5d00", 168=>x"6000", 169=>x"6700", 170=>x"5f00", 171=>x"6100",
---- 172=>x"6300", 173=>x"6900", 174=>x"6800", 175=>x"5f00", 176=>x"6100", 177=>x"6200", 178=>x"6300", 179=>x"6100", 180=>x"5f00",
---- 181=>x"6200", 182=>x"6200", 183=>x"6400", 184=>x"6100", 185=>x"5e00", 186=>x"5f00", 187=>x"6000", 188=>x"6700", 189=>x"6000",
---- 190=>x"5900", 191=>x"5e00", 192=>x"6300", 193=>x"6c00", 194=>x"6100", 195=>x"5a00", 196=>x"6f00", 197=>x"5e00", 198=>x"6000",
---- 199=>x"5d00", 200=>x"5b00", 201=>x"6000", 202=>x"5f00", 203=>x"6700", 204=>x"7500", 205=>x"5a00", 206=>x"5f00", 207=>x"6500",
---- 208=>x"5e00", 209=>x"6000", 210=>x"5d00", 211=>x"5f00", 212=>x"7500", 213=>x"6100", 214=>x"6100", 215=>x"5d00", 216=>x"6f00",
---- 217=>x"6000", 218=>x"6400", 219=>x"6300", 220=>x"5e00", 221=>x"6400", 222=>x"6700", 223=>x"6600", 224=>x"6300", 225=>x"5f00",
---- 226=>x"6400", 227=>x"6500", 228=>x"6500", 229=>x"6400", 230=>x"6d00", 231=>x"6400", 232=>x"6500", 233=>x"6900", 234=>x"6400",
---- 235=>x"6000", 236=>x"6400", 237=>x"7100", 238=>x"6200", 239=>x"7000", 240=>x"5e00", 241=>x"6a00", 242=>x"6500", 243=>x"7000",
---- 244=>x"6500", 245=>x"5f00", 246=>x"7800", 247=>x"6300", 248=>x"6100", 249=>x"6200", 250=>x"5c00", 251=>x"7000", 252=>x"6400",
---- 253=>x"6200", 254=>x"7000", 255=>x"6c00", 256=>x"6d00", 257=>x"5f00", 258=>x"5f00", 259=>x"5a00", 260=>x"6100", 261=>x"6300",
---- 262=>x"6300", 263=>x"6a00", 264=>x"6200", 265=>x"6500", 266=>x"7300", 267=>x"7700", 268=>x"4900", 269=>x"3900", 270=>x"7200",
---- 271=>x"7100", 272=>x"8500", 273=>x"3200", 274=>x"8a00", 275=>x"6900", 276=>x"6c00", 277=>x"6a00", 278=>x"a400", 279=>x"9500",
---- 280=>x"6600", 281=>x"6b00", 282=>x"7500", 283=>x"7a00", 284=>x"9300", 285=>x"6e00", 286=>x"8700", 287=>x"8f00", 288=>x"8800",
---- 289=>x"4600", 290=>x"6900", 291=>x"6c00", 292=>x"7100", 293=>x"4f00", 294=>x"7400", 295=>x"5d00", 296=>x"7e00", 297=>x"8100",
---- 298=>x"6800", 299=>x"5b00", 300=>x"7e00", 301=>x"8500", 302=>x"7200", 303=>x"3800", 304=>x"7a00", 305=>x"7a00", 306=>x"7700",
---- 307=>x"6d00", 308=>x"4800", 309=>x"5d00", 310=>x"6600", 311=>x"7600", 312=>x"5200", 313=>x"5d00", 314=>x"7000", 315=>x"6300",
---- 316=>x"7300", 317=>x"5600", 318=>x"4e00", 319=>x"7800", 320=>x"6300", 321=>x"7a00", 322=>x"4100", 323=>x"4e00", 324=>x"3a00",
---- 325=>x"5d00", 326=>x"9200", 327=>x"4700", 328=>x"4100", 329=>x"6100", 330=>x"8600", 331=>x"7800", 332=>x"5100", 333=>x"6100",
---- 334=>x"5800", 335=>x"6e00", 336=>x"7200", 337=>x"4d00", 338=>x"5b00", 339=>x"3e00", 340=>x"5500", 341=>x"9100", 342=>x"5000",
---- 343=>x"3b00", 344=>x"5700", 345=>x"8000", 346=>x"7500", 347=>x"3d00", 348=>x"3f00", 349=>x"3700", 350=>x"8400", 351=>x"6200",
---- 352=>x"4300", 353=>x"6100", 354=>x"2300", 355=>x"6800", 356=>x"4a00", 357=>x"5600", 358=>x"4b00", 359=>x"2a00", 360=>x"6500",
---- 361=>x"4400", 362=>x"5800", 363=>x"2e00", 364=>x"2f00", 365=>x"6600", 366=>x"4000", 367=>x"5b00", 368=>x"4700", 369=>x"4400",
---- 370=>x"4100", 371=>x"3000", 372=>x"6400", 373=>x"3000", 374=>x"3b00", 375=>x"5f00", 376=>x"3000", 377=>x"4a00", 378=>x"3a00",
---- 379=>x"4100", 380=>x"5c00", 381=>x"2700", 382=>x"5200", 383=>x"3f00", 384=>x"3a00", 385=>x"4000", 386=>x"2100", 387=>x"5200",
---- 388=>x"3400", 389=>x"3000", 390=>x"1e00", 391=>x"2600", 392=>x"2b00", 393=>x"5d00", 394=>x"1500", 395=>x"2400", 396=>x"3200",
---- 397=>x"7700", 398=>x"6c00", 399=>x"5b00", 400=>x"2f00", 401=>x"3b00", 402=>x"3b00", 403=>x"2b00", 404=>x"4a00", 405=>x"2800",
---- 406=>x"4200", 407=>x"3e00", 408=>x"3900", 409=>x"2600", 410=>x"2a00", 411=>x"3a00", 412=>x"3400", 413=>x"3100", 414=>x"2900",
---- 415=>x"2c00", 416=>x"3500", 417=>x"5300", 418=>x"2d00", 419=>x"2400", 420=>x"3700", 421=>x"5200", 422=>x"2500", 423=>x"2900",
---- 424=>x"5500", 425=>x"2d00", 426=>x"2800", 427=>x"2d00", 428=>x"2700", 429=>x"6500", 430=>x"2c00", 431=>x"2e00", 432=>x"3200",
---- 433=>x"4500", 434=>x"2a00", 435=>x"2f00", 436=>x"2f00", 437=>x"2a00", 438=>x"5500", 439=>x"2e00", 440=>x"2600", 441=>x"2f00",
---- 442=>x"4700", 443=>x"3700", 444=>x"2d00", 445=>x"2500", 446=>x"4700", 447=>x"3400", 448=>x"2a00", 449=>x"3600", 450=>x"4200",
---- 451=>x"3000", 452=>x"2d00", 453=>x"3100", 454=>x"3a00", 455=>x"2e00", 456=>x"2a00", 457=>x"2b00", 458=>x"5800", 459=>x"5700",
---- 460=>x"2c00", 461=>x"2d00", 462=>x"3900", 463=>x"3300", 464=>x"3100", 465=>x"3300", 466=>x"3c00", 467=>x"2b00", 468=>x"3300",
---- 469=>x"3000", 470=>x"2f00", 471=>x"2d00", 472=>x"2c00", 473=>x"3700", 474=>x"2e00", 475=>x"3300", 476=>x"3100", 477=>x"5c00",
---- 478=>x"3200", 479=>x"5000", 480=>x"3000", 481=>x"3500", 482=>x"3400", 483=>x"3900", 484=>x"4000", 485=>x"2f00", 486=>x"3400",
---- 487=>x"5900", 488=>x"4800", 489=>x"5300", 490=>x"3000", 491=>x"3a00", 492=>x"3500", 493=>x"4200", 494=>x"4300", 495=>x"3500",
---- 496=>x"3c00", 497=>x"4000", 498=>x"4d00", 499=>x"3700"),
---- 4   => (0=>x"7400", 1=>x"7300", 2=>x"7b00", 3=>x"7c00", 4=>x"7e00", 5=>x"6a00", 6=>x"7300", 7=>x"7c00", 8=>x"7c00", 9=>x"7b00",
---- 10=>x"7100", 11=>x"7400", 12=>x"7600", 13=>x"7b00", 14=>x"7e00", 15=>x"7300", 16=>x"7200", 17=>x"7700", 18=>x"7c00",
---- 19=>x"7e00", 20=>x"6b00", 21=>x"7100", 22=>x"7700", 23=>x"7800", 24=>x"7c00", 25=>x"6b00", 26=>x"7100", 27=>x"7800",
---- 28=>x"7900", 29=>x"7c00", 30=>x"6b00", 31=>x"7000", 32=>x"7700", 33=>x"7a00", 34=>x"7c00", 35=>x"6a00", 36=>x"7100",
---- 37=>x"7500", 38=>x"7600", 39=>x"7900", 40=>x"6900", 41=>x"7100", 42=>x"7800", 43=>x"7700", 44=>x"7d00", 45=>x"6e00",
---- 46=>x"7000", 47=>x"7600", 48=>x"7d00", 49=>x"7c00", 50=>x"6c00", 51=>x"7400", 52=>x"7800", 53=>x"7a00", 54=>x"7b00",
---- 55=>x"7300", 56=>x"7200", 57=>x"7500", 58=>x"7800", 59=>x"7a00", 60=>x"6900", 61=>x"6e00", 62=>x"7500", 63=>x"7500",
---- 64=>x"7600", 65=>x"6800", 66=>x"6b00", 67=>x"7100", 68=>x"7a00", 69=>x"7600", 70=>x"6800", 71=>x"6d00", 72=>x"7000",
---- 73=>x"7900", 74=>x"7300", 75=>x"6700", 76=>x"6e00", 77=>x"7300", 78=>x"7500", 79=>x"7400", 80=>x"6700", 81=>x"6e00",
---- 82=>x"7100", 83=>x"7200", 84=>x"7500", 85=>x"6800", 86=>x"7400", 87=>x"7000", 88=>x"7300", 89=>x"7700", 90=>x"6700",
---- 91=>x"6b00", 92=>x"7200", 93=>x"7400", 94=>x"7600", 95=>x"7200", 96=>x"6b00", 97=>x"7300", 98=>x"7300", 99=>x"7500",
---- 100=>x"6500", 101=>x"6d00", 102=>x"7100", 103=>x"7700", 104=>x"7400", 105=>x"6700", 106=>x"6d00", 107=>x"7300", 108=>x"7200",
---- 109=>x"6a00", 110=>x"6900", 111=>x"6c00", 112=>x"6f00", 113=>x"7500", 114=>x"5f00", 115=>x"6f00", 116=>x"6a00", 117=>x"6e00",
---- 118=>x"6600", 119=>x"8600", 120=>x"6500", 121=>x"6b00", 122=>x"7100", 123=>x"6600", 124=>x"b000", 125=>x"6900", 126=>x"6d00",
---- 127=>x"7100", 128=>x"5e00", 129=>x"ce00", 130=>x"7300", 131=>x"6d00", 132=>x"7100", 133=>x"6700", 134=>x"b000", 135=>x"6500",
---- 136=>x"6c00", 137=>x"6900", 138=>x"6b00", 139=>x"d400", 140=>x"6500", 141=>x"6900", 142=>x"6000", 143=>x"8400", 144=>x"ce00",
---- 145=>x"6400", 146=>x"6a00", 147=>x"5a00", 148=>x"a100", 149=>x"c900", 150=>x"6300", 151=>x"6700", 152=>x"5c00", 153=>x"7f00",
---- 154=>x"c500", 155=>x"6d00", 156=>x"6800", 157=>x"5300", 158=>x"ab00", 159=>x"bc00", 160=>x"6200", 161=>x"6400", 162=>x"4b00",
---- 163=>x"b900", 164=>x"bc00", 165=>x"6100", 166=>x"6200", 167=>x"4400", 168=>x"c900", 169=>x"c600", 170=>x"6c00", 171=>x"5f00",
---- 172=>x"4900", 173=>x"8800", 174=>x"be00", 175=>x"6300", 176=>x"6100", 177=>x"4d00", 178=>x"a500", 179=>x"ba00", 180=>x"6200",
---- 181=>x"6a00", 182=>x"5100", 183=>x"8700", 184=>x"db00", 185=>x"6300", 186=>x"6500", 187=>x"5d00", 188=>x"5c00", 189=>x"da00",
---- 190=>x"5f00", 191=>x"6d00", 192=>x"6100", 193=>x"4800", 194=>x"cb00", 195=>x"5f00", 196=>x"6900", 197=>x"7800", 198=>x"5800",
---- 199=>x"8300", 200=>x"6100", 201=>x"6700", 202=>x"6800", 203=>x"6800", 204=>x"4700", 205=>x"6300", 206=>x"6900", 207=>x"6f00",
---- 208=>x"6f00", 209=>x"5f00", 210=>x"6200", 211=>x"6800", 212=>x"7100", 213=>x"7000", 214=>x"6400", 215=>x"6600", 216=>x"6f00",
---- 217=>x"6e00", 218=>x"7200", 219=>x"6900", 220=>x"6000", 221=>x"7d00", 222=>x"7c00", 223=>x"7100", 224=>x"7000", 225=>x"6500",
---- 226=>x"7300", 227=>x"7000", 228=>x"7800", 229=>x"7600", 230=>x"6700", 231=>x"7000", 232=>x"7800", 233=>x"7100", 234=>x"7000",
---- 235=>x"6700", 236=>x"7200", 237=>x"7a00", 238=>x"7600", 239=>x"7400", 240=>x"6500", 241=>x"6f00", 242=>x"7400", 243=>x"7900",
---- 244=>x"9300", 245=>x"6600", 246=>x"6900", 247=>x"7100", 248=>x"8a00", 249=>x"9200", 250=>x"5d00", 251=>x"6d00", 252=>x"8f00",
---- 253=>x"9400", 254=>x"9800", 255=>x"5900", 256=>x"cd00", 257=>x"9600", 258=>x"8f00", 259=>x"9200", 260=>x"3500", 261=>x"9100",
---- 262=>x"a400", 263=>x"ab00", 264=>x"7300", 265=>x"5d00", 266=>x"a500", 267=>x"d400", 268=>x"9a00", 269=>x"3200", 270=>x"9b00",
---- 271=>x"8500", 272=>x"6000", 273=>x"1d00", 274=>x"4700", 275=>x"4b00", 276=>x"4600", 277=>x"3600", 278=>x"3300", 279=>x"2f00",
---- 280=>x"7c00", 281=>x"5000", 282=>x"6f00", 283=>x"5a00", 284=>x"6a00", 285=>x"5800", 286=>x"3300", 287=>x"3c00", 288=>x"5500",
---- 289=>x"6c00", 290=>x"5500", 291=>x"4200", 292=>x"6200", 293=>x"4200", 294=>x"8100", 295=>x"6500", 296=>x"5900", 297=>x"3d00",
---- 298=>x"3700", 299=>x"7700", 300=>x"5a00", 301=>x"5400", 302=>x"6100", 303=>x"5c00", 304=>x"8300", 305=>x"5400", 306=>x"4b00",
---- 307=>x"6600", 308=>x"4e00", 309=>x"8000", 310=>x"4800", 311=>x"4500", 312=>x"5700", 313=>x"5300", 314=>x"6c00", 315=>x"2b00",
---- 316=>x"7300", 317=>x"4e00", 318=>x"4700", 319=>x"6900", 320=>x"4e00", 321=>x"5200", 322=>x"4e00", 323=>x"5500", 324=>x"6600",
---- 325=>x"5d00", 326=>x"2700", 327=>x"4600", 328=>x"5a00", 329=>x"6b00", 330=>x"3600", 331=>x"4b00", 332=>x"4300", 333=>x"4300",
---- 334=>x"5800", 335=>x"3b00", 336=>x"4d00", 337=>x"4e00", 338=>x"4f00", 339=>x"5e00", 340=>x"4f00", 341=>x"3100", 342=>x"5a00",
---- 343=>x"7100", 344=>x"5d00", 345=>x"4600", 346=>x"4200", 347=>x"5900", 348=>x"6800", 349=>x"5b00", 350=>x"5000", 351=>x"4800",
---- 352=>x"7700", 353=>x"7600", 354=>x"4c00", 355=>x"5000", 356=>x"3400", 357=>x"9b00", 358=>x"5a00", 359=>x"8300", 360=>x"4500",
---- 361=>x"3000", 362=>x"9300", 363=>x"6f00", 364=>x"8a00", 365=>x"3c00", 366=>x"3a00", 367=>x"7300", 368=>x"4c00", 369=>x"7000",
---- 370=>x"3900", 371=>x"2c00", 372=>x"8800", 373=>x"3c00", 374=>x"5900", 375=>x"2f00", 376=>x"2400", 377=>x"8100", 378=>x"7200",
---- 379=>x"4300", 380=>x"3900", 381=>x"2800", 382=>x"7600", 383=>x"8800", 384=>x"5200", 385=>x"7300", 386=>x"3c00", 387=>x"3b00",
---- 388=>x"8a00", 389=>x"7800", 390=>x"6200", 391=>x"5500", 392=>x"2e00", 393=>x"4b00", 394=>x"7900", 395=>x"6800", 396=>x"4500",
---- 397=>x"3800", 398=>x"5d00", 399=>x"3e00", 400=>x"4f00", 401=>x"6600", 402=>x"5500", 403=>x"2900", 404=>x"7a00", 405=>x"5700",
---- 406=>x"4200", 407=>x"2200", 408=>x"4d00", 409=>x"2600", 410=>x"6600", 411=>x"3900", 412=>x"3100", 413=>x"3900", 414=>x"3c00",
---- 415=>x"7800", 416=>x"2b00", 417=>x"3d00", 418=>x"2600", 419=>x"4100", 420=>x"8600", 421=>x"4c00", 422=>x"3200", 423=>x"3d00",
---- 424=>x"3500", 425=>x"6000", 426=>x"2200", 427=>x"3300", 428=>x"3c00", 429=>x"2500", 430=>x"6200", 431=>x"3000", 432=>x"3a00",
---- 433=>x"3500", 434=>x"2a00", 435=>x"4c00", 436=>x"3400", 437=>x"3000", 438=>x"3c00", 439=>x"2900", 440=>x"3e00", 441=>x"3e00",
---- 442=>x"4100", 443=>x"3b00", 444=>x"2c00", 445=>x"4000", 446=>x"3600", 447=>x"4200", 448=>x"3500", 449=>x"3a00", 450=>x"3500",
---- 451=>x"4400", 452=>x"3300", 453=>x"2f00", 454=>x"2900", 455=>x"4800", 456=>x"4600", 457=>x"3d00", 458=>x"2d00", 459=>x"3100",
---- 460=>x"3000", 461=>x"4000", 462=>x"3b00", 463=>x"3700", 464=>x"2f00", 465=>x"3900", 466=>x"3900", 467=>x"4000", 468=>x"3400",
---- 469=>x"2900", 470=>x"2b00", 471=>x"4000", 472=>x"3100", 473=>x"4b00", 474=>x"2c00", 475=>x"2c00", 476=>x"5300", 477=>x"5700",
---- 478=>x"5e00", 479=>x"3700", 480=>x"3100", 481=>x"4e00", 482=>x"2b00", 483=>x"6400", 484=>x"6e00", 485=>x"2300", 486=>x"5900",
---- 487=>x"2000", 488=>x"5400", 489=>x"8000", 490=>x"2800", 491=>x"6e00", 492=>x"2300", 493=>x"6400", 494=>x"5400", 495=>x"5500",
---- 496=>x"5800", 497=>x"3000", 498=>x"6200", 499=>x"3b00"),
---- 5   => (0=>x"8100", 1=>x"8300", 2=>x"8400", 3=>x"8000", 4=>x"8200", 5=>x"8000", 6=>x"8100", 7=>x"8200", 8=>x"8100", 9=>x"8000",
---- 10=>x"7e00", 11=>x"7f00", 12=>x"8100", 13=>x"8200", 14=>x"8200", 15=>x"7f00", 16=>x"8000", 17=>x"8200", 18=>x"8200",
---- 19=>x"8400", 20=>x"7e00", 21=>x"8100", 22=>x"8100", 23=>x"8100", 24=>x"8100", 25=>x"8000", 26=>x"7e00", 27=>x"8000",
---- 28=>x"7f00", 29=>x"8100", 30=>x"7e00", 31=>x"7f00", 32=>x"8000", 33=>x"7d00", 34=>x"7f00", 35=>x"7c00", 36=>x"7d00",
---- 37=>x"7f00", 38=>x"7e00", 39=>x"7b00", 40=>x"7b00", 41=>x"7c00", 42=>x"7d00", 43=>x"7b00", 44=>x"7d00", 45=>x"7b00",
---- 46=>x"7e00", 47=>x"7d00", 48=>x"7e00", 49=>x"8100", 50=>x"8000", 51=>x"7c00", 52=>x"7d00", 53=>x"8200", 54=>x"7e00",
---- 55=>x"7a00", 56=>x"7a00", 57=>x"7d00", 58=>x"7e00", 59=>x"7f00", 60=>x"7a00", 61=>x"7c00", 62=>x"7b00", 63=>x"7d00",
---- 64=>x"7b00", 65=>x"7900", 66=>x"7900", 67=>x"7b00", 68=>x"7d00", 69=>x"7b00", 70=>x"7800", 71=>x"7600", 72=>x"7b00",
---- 73=>x"7900", 74=>x"8500", 75=>x"7b00", 76=>x"7900", 77=>x"7800", 78=>x"7a00", 79=>x"8c00", 80=>x"7800", 81=>x"7900",
---- 82=>x"7900", 83=>x"8000", 84=>x"7100", 85=>x"7900", 86=>x"7800", 87=>x"7f00", 88=>x"7500", 89=>x"6800", 90=>x"7700",
---- 91=>x"7d00", 92=>x"7a00", 93=>x"6a00", 94=>x"7000", 95=>x"7900", 96=>x"8300", 97=>x"6e00", 98=>x"7100", 99=>x"7600",
---- 100=>x"7c00", 101=>x"8000", 102=>x"6400", 103=>x"6a00", 104=>x"7300", 105=>x"a000", 106=>x"7000", 107=>x"6800", 108=>x"6c00",
---- 109=>x"6d00", 110=>x"c900", 111=>x"5f00", 112=>x"6700", 113=>x"6b00", 114=>x"7000", 115=>x"b900", 116=>x"6600", 117=>x"6600",
---- 118=>x"6c00", 119=>x"7100", 120=>x"a400", 121=>x"6100", 122=>x"6500", 123=>x"6b00", 124=>x"7300", 125=>x"8a00", 126=>x"5f00",
---- 127=>x"6600", 128=>x"6e00", 129=>x"6900", 130=>x"8200", 131=>x"5f00", 132=>x"6900", 133=>x"7600", 134=>x"6e00", 135=>x"8000",
---- 136=>x"6800", 137=>x"6800", 138=>x"6400", 139=>x"6200", 140=>x"8b00", 141=>x"7600", 142=>x"6400", 143=>x"6a00", 144=>x"6b00",
---- 145=>x"8f00", 146=>x"7a00", 147=>x"7400", 148=>x"6700", 149=>x"6c00", 150=>x"9d00", 151=>x"8c00", 152=>x"7c00", 153=>x"6b00",
---- 154=>x"6300", 155=>x"9f00", 156=>x"9100", 157=>x"8a00", 158=>x"6b00", 159=>x"5d00", 160=>x"a200", 161=>x"9600", 162=>x"8900",
---- 163=>x"7700", 164=>x"7000", 165=>x"ae00", 166=>x"9000", 167=>x"9700", 168=>x"8600", 169=>x"7b00", 170=>x"b400", 171=>x"9f00",
---- 172=>x"9200", 173=>x"9600", 174=>x"7200", 175=>x"c600", 176=>x"9b00", 177=>x"7800", 178=>x"8500", 179=>x"6900", 180=>x"bf00",
---- 181=>x"9200", 182=>x"7900", 183=>x"8e00", 184=>x"8000", 185=>x"c700", 186=>x"a600", 187=>x"7f00", 188=>x"9500", 189=>x"7400",
---- 190=>x"c600", 191=>x"bd00", 192=>x"9c00", 193=>x"9000", 194=>x"6500", 195=>x"e100", 196=>x"ae00", 197=>x"b500", 198=>x"7600",
---- 199=>x"7d00", 200=>x"c800", 201=>x"c500", 202=>x"ba00", 203=>x"7c00", 204=>x"7e00", 205=>x"8100", 206=>x"df00", 207=>x"c300",
---- 208=>x"8800", 209=>x"7600", 210=>x"8300", 211=>x"bd00", 212=>x"c000", 213=>x"6a00", 214=>x"7900", 215=>x"6f00", 216=>x"f000",
---- 217=>x"8a00", 218=>x"6400", 219=>x"7000", 220=>x"5f00", 221=>x"dc00", 222=>x"7900", 223=>x"7500", 224=>x"6a00", 225=>x"6e00",
---- 226=>x"9500", 227=>x"a000", 228=>x"6700", 229=>x"8000", 230=>x"7000", 231=>x"7500", 232=>x"7800", 233=>x"7b00", 234=>x"8400",
---- 235=>x"9400", 236=>x"6e00", 237=>x"8f00", 238=>x"7600", 239=>x"8100", 240=>x"8500", 241=>x"1500", 242=>x"3600", 243=>x"b300",
---- 244=>x"6300", 245=>x"8200", 246=>x"4800", 247=>x"5700", 248=>x"8100", 249=>x"5100", 250=>x"a300", 251=>x"9b00", 252=>x"5100",
---- 253=>x"2b00", 254=>x"5800", 255=>x"8200", 256=>x"3800", 257=>x"1d00", 258=>x"5e00", 259=>x"4b00", 260=>x"5000", 261=>x"1f00",
---- 262=>x"5900", 263=>x"3700", 264=>x"5500", 265=>x"2000", 266=>x"5f00", 267=>x"4600", 268=>x"3400", 269=>x"5f00", 270=>x"7000",
---- 271=>x"6200", 272=>x"3600", 273=>x"4000", 274=>x"5400", 275=>x"6e00", 276=>x"7700", 277=>x"4800", 278=>x"2c00", 279=>x"4500",
---- 280=>x"5c00", 281=>x"6000", 282=>x"2000", 283=>x"2b00", 284=>x"6500", 285=>x"7b00", 286=>x"3700", 287=>x"2700", 288=>x"5f00",
---- 289=>x"2c00", 290=>x"4400", 291=>x"3200", 292=>x"2c00", 293=>x"4500", 294=>x"4800", 295=>x"5300", 296=>x"3200", 297=>x"3500",
---- 298=>x"4100", 299=>x"2500", 300=>x"6500", 301=>x"5600", 302=>x"5000", 303=>x"2e00", 304=>x"2600", 305=>x"5a00", 306=>x"2800",
---- 307=>x"2d00", 308=>x"2f00", 309=>x"2a00", 310=>x"5400", 311=>x"4d00", 312=>x"3700", 313=>x"3600", 314=>x"2400", 315=>x"8600",
---- 316=>x"6200", 317=>x"2300", 318=>x"4800", 319=>x"2600", 320=>x"7b00", 321=>x"8100", 322=>x"1800", 323=>x"4b00", 324=>x"8900",
---- 325=>x"7200", 326=>x"8700", 327=>x"4d00", 328=>x"4900", 329=>x"6100", 330=>x"4400", 331=>x"8200", 332=>x"7a00", 333=>x"7000",
---- 334=>x"2400", 335=>x"4e00", 336=>x"4900", 337=>x"8700", 338=>x"4f00", 339=>x"3000", 340=>x"5f00", 341=>x"6300", 342=>x"5a00",
---- 343=>x"5500", 344=>x"8b00", 345=>x"6800", 346=>x"5300", 347=>x"5000", 348=>x"6300", 349=>x"9200", 350=>x"5900", 351=>x"6800",
---- 352=>x"5a00", 353=>x"9600", 354=>x"8a00", 355=>x"4800", 356=>x"6900", 357=>x"8000", 358=>x"6c00", 359=>x"7c00", 360=>x"6d00",
---- 361=>x"6400", 362=>x"7a00", 363=>x"5600", 364=>x"6b00", 365=>x"8400", 366=>x"6800", 367=>x"6800", 368=>x"8400", 369=>x"4f00",
---- 370=>x"7500", 371=>x"8900", 372=>x"7900", 373=>x"8e00", 374=>x"5f00", 375=>x"6600", 376=>x"6000", 377=>x"7a00", 378=>x"9700",
---- 379=>x"8800", 380=>x"3000", 381=>x"6400", 382=>x"7c00", 383=>x"7400", 384=>x"8300", 385=>x"6000", 386=>x"9c00", 387=>x"4f00",
---- 388=>x"5b00", 389=>x"7300", 390=>x"5d00", 391=>x"6700", 392=>x"6500", 393=>x"6600", 394=>x"7400", 395=>x"7300", 396=>x"3b00",
---- 397=>x"4e00", 398=>x"7400", 399=>x"8500", 400=>x"3200", 401=>x"4400", 402=>x"5e00", 403=>x"5e00", 404=>x"7c00", 405=>x"6000",
---- 406=>x"3600", 407=>x"5400", 408=>x"6800", 409=>x"7000", 410=>x"5a00", 411=>x"5000", 412=>x"6000", 413=>x"4c00", 414=>x"6000",
---- 415=>x"5c00", 416=>x"4d00", 417=>x"6100", 418=>x"6700", 419=>x"4a00", 420=>x"3200", 421=>x"6600", 422=>x"4f00", 423=>x"6f00",
---- 424=>x"3b00", 425=>x"5400", 426=>x"2b00", 427=>x"3a00", 428=>x"7900", 429=>x"4400", 430=>x"3600", 431=>x"3200", 432=>x"4900",
---- 433=>x"2b00", 434=>x"7b00", 435=>x"3200", 436=>x"4300", 437=>x"3f00", 438=>x"3300", 439=>x"6500", 440=>x"3300", 441=>x"4800",
---- 442=>x"4e00", 443=>x"4200", 444=>x"7000", 445=>x"3c00", 446=>x"3900", 447=>x"4200", 448=>x"4900", 449=>x"3e00", 450=>x"3900",
---- 451=>x"3600", 452=>x"4f00", 453=>x"8300", 454=>x"3000", 455=>x"3000", 456=>x"3300", 457=>x"5000", 458=>x"8400", 459=>x"7c00",
---- 460=>x"3100", 461=>x"3200", 462=>x"4500", 463=>x"5800", 464=>x"9400", 465=>x"2e00", 466=>x"3100", 467=>x"3d00", 468=>x"2300",
---- 469=>x"5900", 470=>x"3300", 471=>x"6300", 472=>x"3e00", 473=>x"3c00", 474=>x"4400", 475=>x"3300", 476=>x"4200", 477=>x"4100",
---- 478=>x"4800", 479=>x"4000", 480=>x"2300", 481=>x"5d00", 482=>x"2200", 483=>x"5e00", 484=>x"3900", 485=>x"2300", 486=>x"6800",
---- 487=>x"3b00", 488=>x"6000", 489=>x"5000", 490=>x"6a00", 491=>x"2a00", 492=>x"5900", 493=>x"2900", 494=>x"6100", 495=>x"6b00",
---- 496=>x"3b00", 497=>x"6f00", 498=>x"2800", 499=>x"4900"),
---- 6   => (0=>x"8300", 1=>x"8200", 2=>x"8500", 3=>x"8500", 4=>x"8600", 5=>x"8300", 6=>x"8200", 7=>x"8600", 8=>x"8400", 9=>x"8100",
---- 10=>x"8000", 11=>x"8200", 12=>x"8100", 13=>x"8400", 14=>x"8200", 15=>x"8100", 16=>x"8300", 17=>x"8400", 18=>x"8500",
---- 19=>x"8600", 20=>x"8100", 21=>x"8100", 22=>x"8200", 23=>x"8300", 24=>x"8300", 25=>x"8200", 26=>x"8100", 27=>x"8100",
---- 28=>x"8000", 29=>x"8300", 30=>x"8100", 31=>x"8300", 32=>x"8100", 33=>x"8200", 34=>x"8000", 35=>x"7e00", 36=>x"7f00",
---- 37=>x"8000", 38=>x"7e00", 39=>x"8000", 40=>x"8100", 41=>x"7f00", 42=>x"7d00", 43=>x"8000", 44=>x"8000", 45=>x"8000",
---- 46=>x"8000", 47=>x"7d00", 48=>x"8200", 49=>x"8200", 50=>x"8000", 51=>x"8000", 52=>x"7d00", 53=>x"7d00", 54=>x"7f00",
---- 55=>x"7f00", 56=>x"7a00", 57=>x"8400", 58=>x"8e00", 59=>x"8e00", 60=>x"8000", 61=>x"8600", 62=>x"8700", 63=>x"8200",
---- 64=>x"7a00", 65=>x"7d00", 66=>x"6c00", 67=>x"7600", 68=>x"7700", 69=>x"7a00", 70=>x"7d00", 71=>x"7000", 72=>x"6f00",
---- 73=>x"7100", 74=>x"7a00", 75=>x"6e00", 76=>x"7100", 77=>x"6e00", 78=>x"7600", 79=>x"7500", 80=>x"6a00", 81=>x"7400",
---- 82=>x"7700", 83=>x"7700", 84=>x"7900", 85=>x"6e00", 86=>x"7100", 87=>x"7700", 88=>x"7500", 89=>x"7600", 90=>x"7100",
---- 91=>x"7500", 92=>x"7900", 93=>x"6f00", 94=>x"6e00", 95=>x"6f00", 96=>x"7500", 97=>x"7100", 98=>x"7700", 99=>x"7800",
---- 100=>x"6f00", 101=>x"7100", 102=>x"7600", 103=>x"7600", 104=>x"8000", 105=>x"7200", 106=>x"7200", 107=>x"7500", 108=>x"7d00",
---- 109=>x"7b00", 110=>x"7200", 111=>x"7000", 112=>x"7700", 113=>x"7f00", 114=>x"8600", 115=>x"7300", 116=>x"7600", 117=>x"7c00",
---- 118=>x"8200", 119=>x"8300", 120=>x"6f00", 121=>x"7500", 122=>x"8200", 123=>x"7d00", 124=>x"7300", 125=>x"7800", 126=>x"7d00",
---- 127=>x"7600", 128=>x"7400", 129=>x"8500", 130=>x"6d00", 131=>x"7500", 132=>x"7900", 133=>x"8100", 134=>x"7c00", 135=>x"7000",
---- 136=>x"6f00", 137=>x"7c00", 138=>x"7300", 139=>x"7600", 140=>x"7000", 141=>x"7600", 142=>x"7200", 143=>x"7e00", 144=>x"7300",
---- 145=>x"6b00", 146=>x"7700", 147=>x"7b00", 148=>x"6f00", 149=>x"9100", 150=>x"6f00", 151=>x"7600", 152=>x"6800", 153=>x"9100",
---- 154=>x"8c00", 155=>x"6c00", 156=>x"6b00", 157=>x"9000", 158=>x"8700", 159=>x"8a00", 160=>x"6c00", 161=>x"8f00", 162=>x"8600",
---- 163=>x"8400", 164=>x"7b00", 165=>x"8800", 166=>x"8000", 167=>x"8800", 168=>x"7500", 169=>x"7d00", 170=>x"7600", 171=>x"8300",
---- 172=>x"6f00", 173=>x"8300", 174=>x"8800", 175=>x"7d00", 176=>x"6900", 177=>x"7f00", 178=>x"8a00", 179=>x"8900", 180=>x"6800",
---- 181=>x"7500", 182=>x"8a00", 183=>x"8500", 184=>x"7700", 185=>x"6f00", 186=>x"8700", 187=>x"8700", 188=>x"7400", 189=>x"8000",
---- 190=>x"8a00", 191=>x"8b00", 192=>x"6a00", 193=>x"7c00", 194=>x"7f00", 195=>x"8100", 196=>x"7100", 197=>x"7d00", 198=>x"7d00",
---- 199=>x"7700", 200=>x"7d00", 201=>x"7600", 202=>x"8500", 203=>x"7f00", 204=>x"7b00", 205=>x"6b00", 206=>x"8100", 207=>x"7300",
---- 208=>x"7600", 209=>x"8200", 210=>x"8000", 211=>x"6900", 212=>x"8600", 213=>x"8a00", 214=>x"7900", 215=>x"7000", 216=>x"7e00",
---- 217=>x"7800", 218=>x"7200", 219=>x"7000", 220=>x"7e00", 221=>x"8500", 222=>x"6600", 223=>x"4e00", 224=>x"3200", 225=>x"8200",
---- 226=>x"8000", 227=>x"5200", 228=>x"3a00", 229=>x"3900", 230=>x"8100", 231=>x"5400", 232=>x"3600", 233=>x"3500", 234=>x"4100",
---- 235=>x"7b00", 236=>x"3500", 237=>x"4c00", 238=>x"3200", 239=>x"4b00", 240=>x"4000", 241=>x"5600", 242=>x"3a00", 243=>x"6000",
---- 244=>x"3700", 245=>x"3b00", 246=>x"5400", 247=>x"5500", 248=>x"4000", 249=>x"5000", 250=>x"6d00", 251=>x"4500", 252=>x"6200",
---- 253=>x"2000", 254=>x"4b00", 255=>x"3f00", 256=>x"5800", 257=>x"6b00", 258=>x"4e00", 259=>x"3400", 260=>x"4c00", 261=>x"6500",
---- 262=>x"6600", 263=>x"2300", 264=>x"2b00", 265=>x"5300", 266=>x"6600", 267=>x"7a00", 268=>x"3000", 269=>x"2f00", 270=>x"3f00",
---- 271=>x"7600", 272=>x"7e00", 273=>x"5b00", 274=>x"2400", 275=>x"6800", 276=>x"5a00", 277=>x"6f00", 278=>x"5000", 279=>x"2e00",
---- 280=>x"5300", 281=>x"7d00", 282=>x"8200", 283=>x"4e00", 284=>x"3300", 285=>x"5b00", 286=>x"5f00", 287=>x"2100", 288=>x"8400",
---- 289=>x"5700", 290=>x"3000", 291=>x"5a00", 292=>x"2000", 293=>x"7900", 294=>x"7900", 295=>x"4000", 296=>x"3200", 297=>x"2e00",
---- 298=>x"7500", 299=>x"7a00", 300=>x"6000", 301=>x"4200", 302=>x"5800", 303=>x"bd00", 304=>x"4e00", 305=>x"6000", 306=>x"6a00",
---- 307=>x"7800", 308=>x"5b00", 309=>x"3400", 310=>x"5800", 311=>x"3700", 312=>x"6d00", 313=>x"3500", 314=>x"1d00", 315=>x"2400",
---- 316=>x"5300", 317=>x"5a00", 318=>x"3d00", 319=>x"1500", 320=>x"1300", 321=>x"5700", 322=>x"2f00", 323=>x"5900", 324=>x"8b00",
---- 325=>x"3400", 326=>x"2800", 327=>x"8f00", 328=>x"a300", 329=>x"9500", 330=>x"3700", 331=>x"7100", 332=>x"9100", 333=>x"c500",
---- 334=>x"5700", 335=>x"9700", 336=>x"9e00", 337=>x"c800", 338=>x"6b00", 339=>x"6f00", 340=>x"9700", 341=>x"b400", 342=>x"8300",
---- 343=>x"5900", 344=>x"9600", 345=>x"8a00", 346=>x"c000", 347=>x"5700", 348=>x"af00", 349=>x"2e00", 350=>x"a500", 351=>x"7200",
---- 352=>x"b700", 353=>x"6900", 354=>x"2900", 355=>x"ac00", 356=>x"b600", 357=>x"6d00", 358=>x"2f00", 359=>x"3300", 360=>x"cd00",
---- 361=>x"9900", 362=>x"1e00", 363=>x"3300", 364=>x"2f00", 365=>x"9700", 366=>x"3a00", 367=>x"2c00", 368=>x"2f00", 369=>x"3100",
---- 370=>x"4900", 371=>x"3600", 372=>x"3d00", 373=>x"6600", 374=>x"2a00", 375=>x"9b00", 376=>x"3a00", 377=>x"2800", 378=>x"2f00",
---- 379=>x"3500", 380=>x"4700", 381=>x"ae00", 382=>x"3e00", 383=>x"2700", 384=>x"3500", 385=>x"5400", 386=>x"8c00", 387=>x"8900",
---- 388=>x"3400", 389=>x"5600", 390=>x"7b00", 391=>x"9300", 392=>x"3f00", 393=>x"7800", 394=>x"3900", 395=>x"8c00", 396=>x"5200",
---- 397=>x"6a00", 398=>x"5000", 399=>x"5700", 400=>x"8e00", 401=>x"7500", 402=>x"5c00", 403=>x"7200", 404=>x"7200", 405=>x"8500",
---- 406=>x"8d00", 407=>x"6a00", 408=>x"7f00", 409=>x"6c00", 410=>x"7400", 411=>x"8e00", 412=>x"8300", 413=>x"1b00", 414=>x"a100",
---- 415=>x"7600", 416=>x"9300", 417=>x"6500", 418=>x"2100", 419=>x"bd00", 420=>x"7800", 421=>x"8900", 422=>x"8000", 423=>x"2e00",
---- 424=>x"9d00", 425=>x"7b00", 426=>x"9500", 427=>x"7b00", 428=>x"8a00", 429=>x"8400", 430=>x"8600", 431=>x"7a00", 432=>x"5200",
---- 433=>x"8400", 434=>x"8000", 435=>x"7600", 436=>x"7700", 437=>x"6100", 438=>x"3400", 439=>x"2700", 440=>x"7900", 441=>x"5a00",
---- 442=>x"7900", 443=>x"6100", 444=>x"3a00", 445=>x"6400", 446=>x"6000", 447=>x"3e00", 448=>x"9d00", 449=>x"6800", 450=>x"2700",
---- 451=>x"4800", 452=>x"6800", 453=>x"6800", 454=>x"3e00", 455=>x"4000", 456=>x"5d00", 457=>x"6b00", 458=>x"4000", 459=>x"3300",
---- 460=>x"7d00", 461=>x"5900", 462=>x"5800", 463=>x"2200", 464=>x"2f00", 465=>x"8a00", 466=>x"6c00", 467=>x"6c00", 468=>x"2b00",
---- 469=>x"4000", 470=>x"6200", 471=>x"6a00", 472=>x"4200", 473=>x"2a00", 474=>x"3f00", 475=>x"7b00", 476=>x"4c00", 477=>x"5700",
---- 478=>x"2200", 479=>x"4a00", 480=>x"7700", 481=>x"6e00", 482=>x"4000", 483=>x"2a00", 484=>x"2a00", 485=>x"5300", 486=>x"6600",
---- 487=>x"3800", 488=>x"2800", 489=>x"2e00", 490=>x"3300", 491=>x"6600", 492=>x"5600", 493=>x"2100", 494=>x"2800", 495=>x"3a00",
---- 496=>x"4000", 497=>x"5700", 498=>x"5f00", 499=>x"3700"),
---- 7   => (0=>x"8300", 1=>x"8600", 2=>x"8200", 3=>x"8500", 4=>x"8500", 5=>x"8400", 6=>x"8200", 7=>x"8500", 8=>x"8400", 9=>x"8400",
---- 10=>x"8300", 11=>x"8400", 12=>x"8300", 13=>x"8300", 14=>x"8100", 15=>x"8400", 16=>x"8400", 17=>x"8300", 18=>x"8400",
---- 19=>x"8400", 20=>x"8100", 21=>x"8200", 22=>x"8300", 23=>x"8100", 24=>x"8100", 25=>x"7f00", 26=>x"8100", 27=>x"8600",
---- 28=>x"8600", 29=>x"7e00", 30=>x"8100", 31=>x"7f00", 32=>x"8300", 33=>x"8200", 34=>x"8000", 35=>x"8300", 36=>x"8000",
---- 37=>x"8000", 38=>x"8000", 39=>x"7d00", 40=>x"8000", 41=>x"7f00", 42=>x"8000", 43=>x"7e00", 44=>x"7d00", 45=>x"8000",
---- 46=>x"7f00", 47=>x"7c00", 48=>x"8400", 49=>x"8500", 50=>x"7e00", 51=>x"7f00", 52=>x"8c00", 53=>x"9800", 54=>x"9100",
---- 55=>x"7c00", 56=>x"8400", 57=>x"8c00", 58=>x"8d00", 59=>x"9100", 60=>x"7900", 61=>x"8000", 62=>x"8500", 63=>x"7f00",
---- 64=>x"8400", 65=>x"7600", 66=>x"8100", 67=>x"8200", 68=>x"8000", 69=>x"8800", 70=>x"7d00", 71=>x"7f00", 72=>x"8300",
---- 73=>x"8800", 74=>x"8500", 75=>x"7e00", 76=>x"7c00", 77=>x"8100", 78=>x"8000", 79=>x"8800", 80=>x"7800", 81=>x"7700",
---- 82=>x"7d00", 83=>x"8400", 84=>x"8500", 85=>x"7200", 86=>x"7b00", 87=>x"7e00", 88=>x"8a00", 89=>x"8100", 90=>x"7b00",
---- 91=>x"8000", 92=>x"8300", 93=>x"8300", 94=>x"8f00", 95=>x"8100", 96=>x"7c00", 97=>x"8600", 98=>x"8900", 99=>x"8400",
---- 100=>x"8300", 101=>x"8b00", 102=>x"8d00", 103=>x"8b00", 104=>x"8c00", 105=>x"8800", 106=>x"8c00", 107=>x"8100", 108=>x"8900",
---- 109=>x"8d00", 110=>x"8700", 111=>x"8a00", 112=>x"8300", 113=>x"8c00", 114=>x"7e00", 115=>x"7d00", 116=>x"8100", 117=>x"8800",
---- 118=>x"7e00", 119=>x"6600", 120=>x"8200", 121=>x"8200", 122=>x"7b00", 123=>x"6400", 124=>x"9900", 125=>x"8600", 126=>x"7f00",
---- 127=>x"6800", 128=>x"9b00", 129=>x"ac00", 130=>x"7600", 131=>x"6900", 132=>x"9a00", 133=>x"a100", 134=>x"9400", 135=>x"7500",
---- 136=>x"9400", 137=>x"9b00", 138=>x"9100", 139=>x"9000", 140=>x"9600", 141=>x"9800", 142=>x"8b00", 143=>x"8900", 144=>x"9000",
---- 145=>x"9100", 146=>x"9000", 147=>x"8300", 148=>x"8f00", 149=>x"9200", 150=>x"9200", 151=>x"7900", 152=>x"8d00", 153=>x"9700",
---- 154=>x"9700", 155=>x"7600", 156=>x"8600", 157=>x"9600", 158=>x"8700", 159=>x"8f00", 160=>x"8a00", 161=>x"9400", 162=>x"8b00",
---- 163=>x"8800", 164=>x"8800", 165=>x"8d00", 166=>x"9000", 167=>x"7f00", 168=>x"8100", 169=>x"9700", 170=>x"8800", 171=>x"7a00",
---- 172=>x"8100", 173=>x"8e00", 174=>x"8100", 175=>x"7a00", 176=>x"8100", 177=>x"8700", 178=>x"7d00", 179=>x"9200", 180=>x"7f00",
---- 181=>x"8800", 182=>x"7c00", 183=>x"8b00", 184=>x"8300", 185=>x"8300", 186=>x"7a00", 187=>x"8a00", 188=>x"8c00", 189=>x"7200",
---- 190=>x"7a00", 191=>x"7f00", 192=>x"7700", 193=>x"7c00", 194=>x"8c00", 195=>x"7e00", 196=>x"8800", 197=>x"7800", 198=>x"4600",
---- 199=>x"4800", 200=>x"7c00", 201=>x"7c00", 202=>x"5d00", 203=>x"6900", 204=>x"4f00", 205=>x"7f00", 206=>x"6500", 207=>x"4b00",
---- 208=>x"3d00", 209=>x"5800", 210=>x"4d00", 211=>x"4400", 212=>x"4c00", 213=>x"2700", 214=>x"4100", 215=>x"2900", 216=>x"4a00",
---- 217=>x"2300", 218=>x"2f00", 219=>x"3100", 220=>x"3400", 221=>x"6400", 222=>x"4800", 223=>x"3a00", 224=>x"2c00", 225=>x"4000",
---- 226=>x"4c00", 227=>x"2f00", 228=>x"3700", 229=>x"5600", 230=>x"2f00", 231=>x"3000", 232=>x"4e00", 233=>x"3600", 234=>x"2b00",
---- 235=>x"2800", 236=>x"5000", 237=>x"4800", 238=>x"2600", 239=>x"3200", 240=>x"2c00", 241=>x"3a00", 242=>x"3500", 243=>x"2f00",
---- 244=>x"2f00", 245=>x"3600", 246=>x"3100", 247=>x"5300", 248=>x"2b00", 249=>x"2000", 250=>x"4000", 251=>x"2600", 252=>x"3200",
---- 253=>x"5800", 254=>x"4b00", 255=>x"4b00", 256=>x"3500", 257=>x"4800", 258=>x"4600", 259=>x"4c00", 260=>x"2d00", 261=>x"5800",
---- 262=>x"2200", 263=>x"2c00", 264=>x"2500", 265=>x"2900", 266=>x"3500", 267=>x"2f00", 268=>x"4f00", 269=>x"2400", 270=>x"2c00",
---- 271=>x"2e00", 272=>x"2f00", 273=>x"2c00", 274=>x"1500", 275=>x"2d00", 276=>x"2e00", 277=>x"3000", 278=>x"2400", 279=>x"3f00",
---- 280=>x"2f00", 281=>x"2a00", 282=>x"3200", 283=>x"2200", 284=>x"7e00", 285=>x"2a00", 286=>x"2f00", 287=>x"2700", 288=>x"4d00",
---- 289=>x"7c00", 290=>x"1d00", 291=>x"2600", 292=>x"1b00", 293=>x"7f00", 294=>x"9000", 295=>x"6e00", 296=>x"1800", 297=>x"4100",
---- 298=>x"7200", 299=>x"c600", 300=>x"6200", 301=>x"700", 302=>x"7800", 303=>x"8600", 304=>x"d600", 305=>x"1c00", 306=>x"4000",
---- 307=>x"7300", 308=>x"b700", 309=>x"8500", 310=>x"2b00", 311=>x"b700", 312=>x"9600", 313=>x"b300", 314=>x"3f00", 315=>x"6500",
---- 316=>x"c000", 317=>x"d100", 318=>x"4a00", 319=>x"2500", 320=>x"7000", 321=>x"7a00", 322=>x"7600", 323=>x"1600", 324=>x"4100",
---- 325=>x"5800", 326=>x"ba00", 327=>x"2300", 328=>x"3400", 329=>x"3700", 330=>x"9700", 331=>x"2e00", 332=>x"2f00", 333=>x"3100",
---- 334=>x"3200", 335=>x"5500", 336=>x"1f00", 337=>x"4d00", 338=>x"2b00", 339=>x"3500", 340=>x"1900", 341=>x"5200", 342=>x"3b00",
---- 343=>x"2600", 344=>x"3d00", 345=>x"3300", 346=>x"2100", 347=>x"5800", 348=>x"4500", 349=>x"4700", 350=>x"3900", 351=>x"4000",
---- 352=>x"2e00", 353=>x"2e00", 354=>x"3300", 355=>x"3700", 356=>x"5c00", 357=>x"2f00", 358=>x"5100", 359=>x"3e00", 360=>x"3700",
---- 361=>x"2e00", 362=>x"3400", 363=>x"2d00", 364=>x"3e00", 365=>x"4800", 366=>x"2c00", 367=>x"3f00", 368=>x"4d00", 369=>x"2700",
---- 370=>x"6c00", 371=>x"2b00", 372=>x"3900", 373=>x"3200", 374=>x"3200", 375=>x"6200", 376=>x"2700", 377=>x"3e00", 378=>x"2d00",
---- 379=>x"3400", 380=>x"4b00", 381=>x"2900", 382=>x"3a00", 383=>x"4b00", 384=>x"4100", 385=>x"5300", 386=>x"2a00", 387=>x"4300",
---- 388=>x"2d00", 389=>x"5200", 390=>x"5200", 391=>x"2700", 392=>x"4100", 393=>x"3500", 394=>x"2a00", 395=>x"3000", 396=>x"3f00",
---- 397=>x"4a00", 398=>x"4d00", 399=>x"2d00", 400=>x"3300", 401=>x"3300", 402=>x"4500", 403=>x"3300", 404=>x"3500", 405=>x"4c00",
---- 406=>x"2900", 407=>x"4400", 408=>x"3600", 409=>x"2f00", 410=>x"4700", 411=>x"2200", 412=>x"4200", 413=>x"3800", 414=>x"2800",
---- 415=>x"4200", 416=>x"2700", 417=>x"4300", 418=>x"4200", 419=>x"2d00", 420=>x"4b00", 421=>x"2c00", 422=>x"4700", 423=>x"3c00",
---- 424=>x"3300", 425=>x"4f00", 426=>x"3200", 427=>x"3700", 428=>x"3a00", 429=>x"3800", 430=>x"6900", 431=>x"5500", 432=>x"4300",
---- 433=>x"4400", 434=>x"3600", 435=>x"2c00", 436=>x"4d00", 437=>x"6400", 438=>x"6100", 439=>x"3a00", 440=>x"3000", 441=>x"2e00",
---- 442=>x"3a00", 443=>x"3000", 444=>x"3900", 445=>x"2a00", 446=>x"7200", 447=>x"2f00", 448=>x"3d00", 449=>x"2b00", 450=>x"3100",
---- 451=>x"2700", 452=>x"2f00", 453=>x"3b00", 454=>x"2c00", 455=>x"2a00", 456=>x"2f00", 457=>x"2b00", 458=>x"2600", 459=>x"3700",
---- 460=>x"2e00", 461=>x"2c00", 462=>x"2600", 463=>x"2800", 464=>x"4500", 465=>x"2800", 466=>x"2500", 467=>x"2900", 468=>x"3b00",
---- 469=>x"5500", 470=>x"2800", 471=>x"2500", 472=>x"3200", 473=>x"4d00", 474=>x"6c00", 475=>x"2600", 476=>x"2700", 477=>x"4700",
---- 478=>x"5d00", 479=>x"3b00", 480=>x"2b00", 481=>x"2a00", 482=>x"3000", 483=>x"3f00", 484=>x"5100", 485=>x"2a00", 486=>x"3b00",
---- 487=>x"5a00", 488=>x"7100", 489=>x"7100", 490=>x"3b00", 491=>x"5800", 492=>x"7400", 493=>x"7000", 494=>x"7700", 495=>x"5300",
---- 496=>x"5f00", 497=>x"6c00", 498=>x"7500", 499=>x"7800"),
---- 8   => (0=>x"8600", 1=>x"8500", 2=>x"8000", 3=>x"8000", 4=>x"8500", 5=>x"8400", 6=>x"8400", 7=>x"8100", 8=>x"8100", 9=>x"8400",
---- 10=>x"8200", 11=>x"8300", 12=>x"8100", 13=>x"8200", 14=>x"8100", 15=>x"8400", 16=>x"8400", 17=>x"8500", 18=>x"8000",
---- 19=>x"8400", 20=>x"8200", 21=>x"8000", 22=>x"8000", 23=>x"8100", 24=>x"8100", 25=>x"7c00", 26=>x"7a00", 27=>x"7e00",
---- 28=>x"7f00", 29=>x"7d00", 30=>x"7a00", 31=>x"7a00", 32=>x"7900", 33=>x"7d00", 34=>x"7d00", 35=>x"7c00", 36=>x"7a00",
---- 37=>x"7b00", 38=>x"7b00", 39=>x"7900", 40=>x"8000", 41=>x"7a00", 42=>x"7800", 43=>x"7900", 44=>x"7900", 45=>x"8800",
---- 46=>x"8d00", 47=>x"8b00", 48=>x"9e00", 49=>x"b500", 50=>x"9300", 51=>x"a100", 52=>x"a200", 53=>x"af00", 54=>x"b600",
---- 55=>x"9600", 56=>x"9400", 57=>x"9c00", 58=>x"9e00", 59=>x"a700", 60=>x"8e00", 61=>x"9600", 62=>x"a000", 63=>x"9c00",
---- 64=>x"a700", 65=>x"8500", 66=>x"8a00", 67=>x"9500", 68=>x"a100", 69=>x"a000", 70=>x"8700", 71=>x"8b00", 72=>x"8d00",
---- 73=>x"9b00", 74=>x"a100", 75=>x"8100", 76=>x"8500", 77=>x"8d00", 78=>x"9700", 79=>x"a200", 80=>x"8300", 81=>x"8900",
---- 82=>x"8700", 83=>x"9600", 84=>x"9400", 85=>x"8900", 86=>x"8d00", 87=>x"9100", 88=>x"9500", 89=>x"9f00", 90=>x"9100",
---- 91=>x"8f00", 92=>x"8b00", 93=>x"8b00", 94=>x"9d00", 95=>x"8e00", 96=>x"8800", 97=>x"8900", 98=>x"8e00", 99=>x"a000",
---- 100=>x"8900", 101=>x"8600", 102=>x"8700", 103=>x"7f00", 104=>x"8500", 105=>x"8500", 106=>x"7700", 107=>x"7400", 108=>x"a200",
---- 109=>x"bc00", 110=>x"7300", 111=>x"7900", 112=>x"ac00", 113=>x"c500", 114=>x"a000", 115=>x"8b00", 116=>x"b500", 117=>x"b300",
---- 118=>x"b400", 119=>x"b300", 120=>x"b600", 121=>x"ad00", 122=>x"a800", 123=>x"aa00", 124=>x"aa00", 125=>x"a300", 126=>x"a600",
---- 127=>x"8200", 128=>x"b600", 129=>x"b600", 130=>x"9900", 131=>x"a200", 132=>x"a700", 133=>x"b300", 134=>x"b500", 135=>x"9400",
---- 136=>x"a300", 137=>x"b300", 138=>x"9000", 139=>x"a200", 140=>x"a200", 141=>x"a500", 142=>x"9c00", 143=>x"a900", 144=>x"af00",
---- 145=>x"8b00", 146=>x"9500", 147=>x"ab00", 148=>x"ae00", 149=>x"a100", 150=>x"8e00", 151=>x"9300", 152=>x"9f00", 153=>x"9c00",
---- 154=>x"a500", 155=>x"9300", 156=>x"9b00", 157=>x"8e00", 158=>x"9900", 159=>x"9e00", 160=>x"9700", 161=>x"8900", 162=>x"9300",
---- 163=>x"9300", 164=>x"a200", 165=>x"8500", 166=>x"9800", 167=>x"9a00", 168=>x"7e00", 169=>x"7b00", 170=>x"9900", 171=>x"8e00",
---- 172=>x"7100", 173=>x"8a00", 174=>x"7000", 175=>x"8000", 176=>x"7e00", 177=>x"8c00", 178=>x"6900", 179=>x"7300", 180=>x"7300",
---- 181=>x"8b00", 182=>x"7100", 183=>x"7400", 184=>x"5a00", 185=>x"8800", 186=>x"6400", 187=>x"4600", 188=>x"5100", 189=>x"3e00",
---- 190=>x"5500", 191=>x"4000", 192=>x"4d00", 193=>x"2a00", 194=>x"3200", 195=>x"4800", 196=>x"4f00", 197=>x"2e00", 198=>x"5800",
---- 199=>x"1e00", 200=>x"5500", 201=>x"2400", 202=>x"3700", 203=>x"5900", 204=>x"2d00", 205=>x"4600", 206=>x"2e00", 207=>x"4000",
---- 208=>x"6800", 209=>x"3c00", 210=>x"4a00", 211=>x"4600", 212=>x"3900", 213=>x"5800", 214=>x"5200", 215=>x"4b00", 216=>x"4500",
---- 217=>x"4700", 218=>x"2200", 219=>x"7900", 220=>x"3100", 221=>x"3800", 222=>x"5200", 223=>x"6300", 224=>x"6c00", 225=>x"3600",
---- 226=>x"2d00", 227=>x"4e00", 228=>x"4600", 229=>x"6000", 230=>x"3f00", 231=>x"3b00", 232=>x"2b00", 233=>x"4a00", 234=>x"1200",
---- 235=>x"3800", 236=>x"4900", 237=>x"3e00", 238=>x"4e00", 239=>x"4400", 240=>x"4500", 241=>x"4a00", 242=>x"3d00", 243=>x"2600",
---- 244=>x"8100", 245=>x"3600", 246=>x"5300", 247=>x"1800", 248=>x"7500", 249=>x"9600", 250=>x"2800", 251=>x"1e00", 252=>x"4700",
---- 253=>x"8b00", 254=>x"b400", 255=>x"2f00", 256=>x"1b00", 257=>x"7d00", 258=>x"ae00", 259=>x"ad00", 260=>x"2200", 261=>x"5900",
---- 262=>x"8800", 263=>x"a900", 264=>x"b800", 265=>x"2f00", 266=>x"7e00", 267=>x"aa00", 268=>x"b200", 269=>x"d000", 270=>x"7100",
---- 271=>x"7b00", 272=>x"b100", 273=>x"cd00", 274=>x"aa00", 275=>x"7d00", 276=>x"9d00", 277=>x"c200", 278=>x"b800", 279=>x"5600",
---- 280=>x"8c00", 281=>x"b300", 282=>x"c600", 283=>x"3b00", 284=>x"6800", 285=>x"b400", 286=>x"cf00", 287=>x"4800", 288=>x"4200",
---- 289=>x"7600", 290=>x"d400", 291=>x"6500", 292=>x"1d00", 293=>x"5500", 294=>x"7800", 295=>x"d600", 296=>x"1400", 297=>x"3500",
---- 298=>x"5000", 299=>x"7400", 300=>x"3000", 301=>x"1d00", 302=>x"4300", 303=>x"4c00", 304=>x"7000", 305=>x"1400", 306=>x"2400",
---- 307=>x"5300", 308=>x"4b00", 309=>x"6d00", 310=>x"2000", 311=>x"2600", 312=>x"5d00", 313=>x"4800", 314=>x"7100", 315=>x"3d00",
---- 316=>x"2500", 317=>x"6200", 318=>x"5400", 319=>x"6f00", 320=>x"3300", 321=>x"2600", 322=>x"6d00", 323=>x"5600", 324=>x"7300",
---- 325=>x"3a00", 326=>x"2a00", 327=>x"6a00", 328=>x"5e00", 329=>x"7600", 330=>x"3f00", 331=>x"2500", 332=>x"5e00", 333=>x"6100",
---- 334=>x"7100", 335=>x"4b00", 336=>x"2400", 337=>x"5600", 338=>x"5c00", 339=>x"6a00", 340=>x"5800", 341=>x"2400", 342=>x"5100",
---- 343=>x"5300", 344=>x"6000", 345=>x"4f00", 346=>x"2e00", 347=>x"4d00", 348=>x"4f00", 349=>x"5700", 350=>x"5200", 351=>x"3500",
---- 352=>x"5900", 353=>x"4800", 354=>x"4a00", 355=>x"3f00", 356=>x"3c00", 357=>x"3b00", 358=>x"4b00", 359=>x"4000", 360=>x"4700",
---- 361=>x"3e00", 362=>x"3000", 363=>x"4100", 364=>x"3a00", 365=>x"5700", 366=>x"3700", 367=>x"3400", 368=>x"3c00", 369=>x"3800",
---- 370=>x"2d00", 371=>x"3900", 372=>x"3800", 373=>x"3800", 374=>x"3b00", 375=>x"2f00", 376=>x"3000", 377=>x"3c00", 378=>x"3d00",
---- 379=>x"3b00", 380=>x"4400", 381=>x"2d00", 382=>x"3700", 383=>x"3900", 384=>x"3800", 385=>x"2f00", 386=>x"3100", 387=>x"3000",
---- 388=>x"3e00", 389=>x"3700", 390=>x"3700", 391=>x"4300", 392=>x"4200", 393=>x"3800", 394=>x"4400", 395=>x"3800", 396=>x"3b00",
---- 397=>x"2f00", 398=>x"3b00", 399=>x"4900", 400=>x"3900", 401=>x"3d00", 402=>x"3400", 403=>x"4400", 404=>x"5300", 405=>x"3300",
---- 406=>x"3f00", 407=>x"2c00", 408=>x"4000", 409=>x"5f00", 410=>x"5a00", 411=>x"3c00", 412=>x"3100", 413=>x"3400", 414=>x"6c00",
---- 415=>x"3400", 416=>x"3500", 417=>x"3000", 418=>x"3c00", 419=>x"6b00", 420=>x"3400", 421=>x"3800", 422=>x"2f00", 423=>x"5900",
---- 424=>x"6e00", 425=>x"3500", 426=>x"2f00", 427=>x"3a00", 428=>x"7400", 429=>x"7f00", 430=>x"3600", 431=>x"2f00", 432=>x"4900",
---- 433=>x"7700", 434=>x"7f00", 435=>x"2f00", 436=>x"3a00", 437=>x"5900", 438=>x"7d00", 439=>x"8400", 440=>x"2800", 441=>x"4a00",
---- 442=>x"6600", 443=>x"7d00", 444=>x"8500", 445=>x"3000", 446=>x"5600", 447=>x"7300", 448=>x"7d00", 449=>x"7e00", 450=>x"4100",
---- 451=>x"6500", 452=>x"7400", 453=>x"8000", 454=>x"6500", 455=>x"5300", 456=>x"7700", 457=>x"7700", 458=>x"7a00", 459=>x"2a00",
---- 460=>x"6600", 461=>x"7500", 462=>x"8400", 463=>x"4000", 464=>x"3500", 465=>x"7600", 466=>x"7e00", 467=>x"4f00", 468=>x"3300",
---- 469=>x"6f00", 470=>x"7800", 471=>x"3f00", 472=>x"2600", 473=>x"6c00", 474=>x"7f00", 475=>x"2900", 476=>x"4700", 477=>x"7000",
---- 478=>x"7e00", 479=>x"7e00", 480=>x"6a00", 481=>x"7900", 482=>x"7c00", 483=>x"7e00", 484=>x"7f00", 485=>x"7a00", 486=>x"7d00",
---- 487=>x"7e00", 488=>x"8000", 489=>x"7f00", 490=>x"7600", 491=>x"7e00", 492=>x"8000", 493=>x"7c00", 494=>x"8200", 495=>x"7a00",
---- 496=>x"7d00", 497=>x"7e00", 498=>x"8000", 499=>x"8000"),
---- 9   => (0=>x"8300", 1=>x"8300", 2=>x"8500", 3=>x"8600", 4=>x"8200", 5=>x"8100", 6=>x"8100", 7=>x"8400", 8=>x"8200", 9=>x"8200",
---- 10=>x"8000", 11=>x"8200", 12=>x"8500", 13=>x"8300", 14=>x"8000", 15=>x"8100", 16=>x"8200", 17=>x"8600", 18=>x"8800",
---- 19=>x"8300", 20=>x"7f00", 21=>x"7f00", 22=>x"8400", 23=>x"8700", 24=>x"8300", 25=>x"7e00", 26=>x"7d00", 27=>x"8000",
---- 28=>x"8100", 29=>x"8300", 30=>x"7d00", 31=>x"7b00", 32=>x"7f00", 33=>x"8100", 34=>x"7f00", 35=>x"7600", 36=>x"7900",
---- 37=>x"7d00", 38=>x"7f00", 39=>x"8100", 40=>x"7300", 41=>x"6e00", 42=>x"7200", 43=>x"7900", 44=>x"8000", 45=>x"b700",
---- 46=>x"b800", 47=>x"a300", 48=>x"8a00", 49=>x"7200", 50=>x"b200", 51=>x"a700", 52=>x"aa00", 53=>x"c100", 54=>x"c300",
---- 55=>x"af00", 56=>x"9500", 57=>x"ac00", 58=>x"bd00", 59=>x"aa00", 60=>x"b000", 61=>x"b800", 62=>x"b800", 63=>x"a000",
---- 64=>x"ba00", 65=>x"9b00", 66=>x"b600", 67=>x"b700", 68=>x"bc00", 69=>x"a500", 70=>x"ad00", 71=>x"b400", 72=>x"b600",
---- 73=>x"be00", 74=>x"c000", 75=>x"9e00", 76=>x"b500", 77=>x"bd00", 78=>x"ba00", 79=>x"be00", 80=>x"b500", 81=>x"b700",
---- 82=>x"9800", 83=>x"bf00", 84=>x"b600", 85=>x"ac00", 86=>x"b200", 87=>x"b100", 88=>x"a400", 89=>x"b600", 90=>x"9700",
---- 91=>x"9c00", 92=>x"a200", 93=>x"d000", 94=>x"cd00", 95=>x"8900", 96=>x"ad00", 97=>x"c800", 98=>x"c900", 99=>x"d000",
---- 100=>x"bf00", 101=>x"b200", 102=>x"c300", 103=>x"c000", 104=>x"c300", 105=>x"b600", 106=>x"c000", 107=>x"c100", 108=>x"b900",
---- 109=>x"bf00", 110=>x"af00", 111=>x"ba00", 112=>x"af00", 113=>x"be00", 114=>x"ab00", 115=>x"ac00", 116=>x"b600", 117=>x"bc00",
---- 118=>x"bb00", 119=>x"c200", 120=>x"a500", 121=>x"ae00", 122=>x"c000", 123=>x"bf00", 124=>x"a200", 125=>x"b100", 126=>x"be00",
---- 127=>x"b600", 128=>x"ba00", 129=>x"b700", 130=>x"b300", 131=>x"af00", 132=>x"b900", 133=>x"a900", 134=>x"af00", 135=>x"af00",
---- 136=>x"bb00", 137=>x"a000", 138=>x"b100", 139=>x"b100", 140=>x"a800", 141=>x"9300", 142=>x"b000", 143=>x"af00", 144=>x"ad00",
---- 145=>x"a400", 146=>x"af00", 147=>x"ac00", 148=>x"a900", 149=>x"9100", 150=>x"ae00", 151=>x"aa00", 152=>x"9100", 153=>x"ae00",
---- 154=>x"ae00", 155=>x"a700", 156=>x"a700", 157=>x"aa00", 158=>x"9f00", 159=>x"a600", 160=>x"9f00", 161=>x"9900", 162=>x"8c00",
---- 163=>x"a900", 164=>x"9e00", 165=>x"8c00", 166=>x"8d00", 167=>x"8a00", 168=>x"6100", 169=>x"9e00", 170=>x"5500", 171=>x"4c00",
---- 172=>x"b000", 173=>x"9e00", 174=>x"7300", 175=>x"6a00", 176=>x"5600", 177=>x"7f00", 178=>x"7f00", 179=>x"5000", 180=>x"4000",
---- 181=>x"3600", 182=>x"5a00", 183=>x"6d00", 184=>x"5c00", 185=>x"2b00", 186=>x"5200", 187=>x"7c00", 188=>x"3000", 189=>x"4e00",
---- 190=>x"2c00", 191=>x"7400", 192=>x"3800", 193=>x"4800", 194=>x"7000", 195=>x"4e00", 196=>x"3a00", 197=>x"3100", 198=>x"4f00",
---- 199=>x"5800", 200=>x"6200", 201=>x"3300", 202=>x"4400", 203=>x"3700", 204=>x"4800", 205=>x"2800", 206=>x"3200", 207=>x"3800",
---- 208=>x"3c00", 209=>x"5c00", 210=>x"2900", 211=>x"2d00", 212=>x"2000", 213=>x"2e00", 214=>x"7300", 215=>x"4100", 216=>x"1a00",
---- 217=>x"5200", 218=>x"9b00", 219=>x"8400", 220=>x"1800", 221=>x"1e00", 222=>x"8a00", 223=>x"7200", 224=>x"b800", 225=>x"2a00",
---- 226=>x"7e00", 227=>x"8500", 228=>x"ab00", 229=>x"bd00", 230=>x"7d00", 231=>x"8800", 232=>x"a700", 233=>x"9800", 234=>x"b200",
---- 235=>x"6d00", 236=>x"ac00", 237=>x"ac00", 238=>x"9700", 239=>x"b500", 240=>x"ab00", 241=>x"a700", 242=>x"bc00", 243=>x"8b00",
---- 244=>x"c500", 245=>x"af00", 246=>x"b400", 247=>x"a600", 248=>x"bd00", 249=>x"b000", 250=>x"b800", 251=>x"c900", 252=>x"c000",
---- 253=>x"9300", 254=>x"5300", 255=>x"c300", 256=>x"cc00", 257=>x"9900", 258=>x"3600", 259=>x"3700", 260=>x"d200", 261=>x"ab00",
---- 262=>x"5f00", 263=>x"4b00", 264=>x"2800", 265=>x"a100", 266=>x"6d00", 267=>x"7f00", 268=>x"9100", 269=>x"5e00", 270=>x"5d00",
---- 271=>x"8400", 272=>x"8b00", 273=>x"9200", 274=>x"9000", 275=>x"7600", 276=>x"8a00", 277=>x"8e00", 278=>x"9a00", 279=>x"9d00",
---- 280=>x"7c00", 281=>x"8900", 282=>x"9700", 283=>x"a200", 284=>x"a600", 285=>x"7e00", 286=>x"8700", 287=>x"9400", 288=>x"9f00",
---- 289=>x"aa00", 290=>x"7e00", 291=>x"8400", 292=>x"9100", 293=>x"8b00", 294=>x"a600", 295=>x"7f00", 296=>x"8400", 297=>x"8e00",
---- 298=>x"9900", 299=>x"9c00", 300=>x"7e00", 301=>x"8200", 302=>x"8a00", 303=>x"8c00", 304=>x"9c00", 305=>x"7c00", 306=>x"8300",
---- 307=>x"8800", 308=>x"9000", 309=>x"9800", 310=>x"7e00", 311=>x"8000", 312=>x"8700", 313=>x"8f00", 314=>x"8a00", 315=>x"7a00",
---- 316=>x"8000", 317=>x"8700", 318=>x"8700", 319=>x"9500", 320=>x"7b00", 321=>x"7f00", 322=>x"8300", 323=>x"8b00", 324=>x"9200",
---- 325=>x"7d00", 326=>x"7e00", 327=>x"8500", 328=>x"8c00", 329=>x"8c00", 330=>x"7d00", 331=>x"8100", 332=>x"8400", 333=>x"8800",
---- 334=>x"8b00", 335=>x"7d00", 336=>x"8000", 337=>x"8400", 338=>x"8700", 339=>x"8c00", 340=>x"7a00", 341=>x"8200", 342=>x"7d00",
---- 343=>x"8500", 344=>x"8c00", 345=>x"7500", 346=>x"7a00", 347=>x"7d00", 348=>x"8100", 349=>x"8600", 350=>x"6b00", 351=>x"7700",
---- 352=>x"7600", 353=>x"7d00", 354=>x"8100", 355=>x"6600", 356=>x"6a00", 357=>x"6f00", 358=>x"7800", 359=>x"8100", 360=>x"4900",
---- 361=>x"5f00", 362=>x"6b00", 363=>x"7500", 364=>x"7e00", 365=>x"4200", 366=>x"3800", 367=>x"5800", 368=>x"6a00", 369=>x"7d00",
---- 370=>x"4400", 371=>x"2e00", 372=>x"2e00", 373=>x"4d00", 374=>x"6f00", 375=>x"5600", 376=>x"5700", 377=>x"3600", 378=>x"4100",
---- 379=>x"4600", 380=>x"2b00", 381=>x"5500", 382=>x"5e00", 383=>x"8000", 384=>x"8400", 385=>x"3200", 386=>x"4a00", 387=>x"6c00",
---- 388=>x"7d00", 389=>x"7d00", 390=>x"3100", 391=>x"4000", 392=>x"6a00", 393=>x"7500", 394=>x"7b00", 395=>x"3700", 396=>x"4100",
---- 397=>x"6700", 398=>x"7a00", 399=>x"7d00", 400=>x"4d00", 401=>x"3200", 402=>x"6d00", 403=>x"7900", 404=>x"7400", 405=>x"6500",
---- 406=>x"2b00", 407=>x"6c00", 408=>x"7200", 409=>x"8300", 410=>x"7200", 411=>x"2400", 412=>x"6300", 413=>x"7e00", 414=>x"8500",
---- 415=>x"7800", 416=>x"2b00", 417=>x"6600", 418=>x"8000", 419=>x"7e00", 420=>x"7a00", 421=>x"2f00", 422=>x"6800", 423=>x"8400",
---- 424=>x"8300", 425=>x"7400", 426=>x"3600", 427=>x"6c00", 428=>x"8000", 429=>x"8700", 430=>x"6f00", 431=>x"3900", 432=>x"7100",
---- 433=>x"8400", 434=>x"8300", 435=>x"6500", 436=>x"4700", 437=>x"7a00", 438=>x"8400", 439=>x"8700", 440=>x"4e00", 441=>x"5600",
---- 442=>x"8100", 443=>x"8500", 444=>x"8900", 445=>x"3a00", 446=>x"6900", 447=>x"8700", 448=>x"8a00", 449=>x"8b00", 450=>x"3800",
---- 451=>x"7e00", 452=>x"8700", 453=>x"8900", 454=>x"8c00", 455=>x"6000", 456=>x"8700", 457=>x"8600", 458=>x"8700", 459=>x"8c00",
---- 460=>x"7f00", 461=>x"8800", 462=>x"8800", 463=>x"8a00", 464=>x"8b00", 465=>x"8400", 466=>x"8700", 467=>x"8800", 468=>x"8b00",
---- 469=>x"8a00", 470=>x"8200", 471=>x"8600", 472=>x"8a00", 473=>x"8c00", 474=>x"8500", 475=>x"8300", 476=>x"8700", 477=>x"8800",
---- 478=>x"8900", 479=>x"8d00", 480=>x"8000", 481=>x"8400", 482=>x"8500", 483=>x"8a00", 484=>x"8800", 485=>x"7e00", 486=>x"8500",
---- 487=>x"8800", 488=>x"8600", 489=>x"8900", 490=>x"8400", 491=>x"8200", 492=>x"8500", 493=>x"8800", 494=>x"8700", 495=>x"8400",
---- 496=>x"8100", 497=>x"8600", 498=>x"8a00", 499=>x"8500"),
---- 10  => (0=>x"8900", 1=>x"8000", 2=>x"8300", 3=>x"8000", 4=>x"8300", 5=>x"8500", 6=>x"8000", 7=>x"8000", 8=>x"7f00", 9=>x"7f00",
---- 10=>x"8100", 11=>x"8300", 12=>x"8000", 13=>x"8000", 14=>x"8000", 15=>x"8200", 16=>x"8300", 17=>x"8000", 18=>x"8000",
---- 19=>x"8000", 20=>x"8100", 21=>x"8200", 22=>x"8000", 23=>x"8000", 24=>x"7e00", 25=>x"8200", 26=>x"8200", 27=>x"7e00",
---- 28=>x"7e00", 29=>x"7f00", 30=>x"8400", 31=>x"8000", 32=>x"7e00", 33=>x"7f00", 34=>x"7f00", 35=>x"8400", 36=>x"7f00",
---- 37=>x"7f00", 38=>x"8000", 39=>x"7e00", 40=>x"8000", 41=>x"7f00", 42=>x"7f00", 43=>x"7e00", 44=>x"7f00", 45=>x"7000",
---- 46=>x"7a00", 47=>x"7c00", 48=>x"8000", 49=>x"8300", 50=>x"a400", 51=>x"7400", 52=>x"7000", 53=>x"7c00", 54=>x"7e00",
---- 55=>x"ca00", 56=>x"c900", 57=>x"9700", 58=>x"6a00", 59=>x"7a00", 60=>x"be00", 61=>x"c300", 62=>x"cc00", 63=>x"b500",
---- 64=>x"6f00", 65=>x"c100", 66=>x"c200", 67=>x"c500", 68=>x"c500", 69=>x"cb00", 70=>x"a200", 71=>x"c700", 72=>x"c400",
---- 73=>x"c200", 74=>x"c600", 75=>x"c300", 76=>x"c100", 77=>x"ba00", 78=>x"bf00", 79=>x"ca00", 80=>x"b000", 81=>x"be00",
---- 82=>x"d300", 83=>x"d600", 84=>x"d400", 85=>x"d500", 86=>x"d500", 87=>x"b500", 88=>x"c800", 89=>x"b400", 90=>x"cb00",
---- 91=>x"d300", 92=>x"cd00", 93=>x"c900", 94=>x"cd00", 95=>x"b400", 96=>x"bb00", 97=>x"c700", 98=>x"a500", 99=>x"cb00",
---- 100=>x"9800", 101=>x"be00", 102=>x"c900", 103=>x"ce00", 104=>x"ce00", 105=>x"c700", 106=>x"a800", 107=>x"d200", 108=>x"cd00",
---- 109=>x"c200", 110=>x"c700", 111=>x"ca00", 112=>x"b200", 113=>x"c500", 114=>x"b200", 115=>x"c600", 116=>x"a600", 117=>x"c400",
---- 118=>x"c200", 119=>x"c600", 120=>x"c200", 121=>x"bb00", 122=>x"c000", 123=>x"c500", 124=>x"c900", 125=>x"ae00", 126=>x"bc00",
---- 127=>x"c500", 128=>x"c600", 129=>x"c300", 130=>x"b600", 131=>x"be00", 132=>x"b900", 133=>x"c200", 134=>x"c100", 135=>x"b800",
---- 136=>x"b000", 137=>x"b500", 138=>x"b400", 139=>x"c400", 140=>x"ae00", 141=>x"ad00", 142=>x"b100", 143=>x"bf00", 144=>x"af00",
---- 145=>x"b400", 146=>x"9c00", 147=>x"9f00", 148=>x"b600", 149=>x"b800", 150=>x"a100", 151=>x"aa00", 152=>x"a800", 153=>x"a900",
---- 154=>x"aa00", 155=>x"a600", 156=>x"a100", 157=>x"a000", 158=>x"a600", 159=>x"ae00", 160=>x"8f00", 161=>x"a300", 162=>x"9400",
---- 163=>x"a600", 164=>x"a700", 165=>x"ac00", 166=>x"a000", 167=>x"9d00", 168=>x"a700", 169=>x"a600", 170=>x"7500", 171=>x"7700",
---- 172=>x"7d00", 173=>x"7300", 174=>x"6f00", 175=>x"4400", 176=>x"5b00", 177=>x"5c00", 178=>x"3000", 179=>x"2400", 180=>x"6b00",
---- 181=>x"4600", 182=>x"4a00", 183=>x"2e00", 184=>x"1400", 185=>x"5800", 186=>x"4600", 187=>x"4200", 188=>x"2000", 189=>x"8c00",
---- 190=>x"4200", 191=>x"2900", 192=>x"4600", 193=>x"8f00", 194=>x"8900", 195=>x"4800", 196=>x"4b00", 197=>x"8500", 198=>x"8300",
---- 199=>x"c300", 200=>x"6500", 201=>x"7f00", 202=>x"6900", 203=>x"c300", 204=>x"c500", 205=>x"4c00", 206=>x"7300", 207=>x"a500",
---- 208=>x"b000", 209=>x"a400", 210=>x"8000", 211=>x"9d00", 212=>x"b800", 213=>x"b800", 214=>x"bb00", 215=>x"a400", 216=>x"9a00",
---- 217=>x"b400", 218=>x"c000", 219=>x"9e00", 220=>x"a200", 221=>x"9200", 222=>x"b200", 223=>x"bb00", 224=>x"a900", 225=>x"b200",
---- 226=>x"8a00", 227=>x"c100", 228=>x"b600", 229=>x"a300", 230=>x"ab00", 231=>x"9000", 232=>x"9900", 233=>x"9900", 234=>x"9e00",
---- 235=>x"ae00", 236=>x"bb00", 237=>x"8300", 238=>x"9100", 239=>x"a600", 240=>x"bd00", 241=>x"7500", 242=>x"7700", 243=>x"6a00",
---- 244=>x"4f00", 245=>x"7300", 246=>x"9100", 247=>x"8100", 248=>x"a500", 249=>x"7200", 250=>x"4000", 251=>x"3600", 252=>x"2900",
---- 253=>x"3500", 254=>x"3b00", 255=>x"2f00", 256=>x"2a00", 257=>x"3100", 258=>x"9e00", 259=>x"5100", 260=>x"6a00", 261=>x"4500",
---- 262=>x"3b00", 263=>x"c500", 264=>x"d900", 265=>x"6800", 266=>x"7800", 267=>x"a000", 268=>x"d100", 269=>x"b100", 270=>x"8b00",
---- 271=>x"7200", 272=>x"7f00", 273=>x"7600", 274=>x"9a00", 275=>x"8d00", 276=>x"9500", 277=>x"9600", 278=>x"a100", 279=>x"a400",
---- 280=>x"af00", 281=>x"aa00", 282=>x"ac00", 283=>x"aa00", 284=>x"ac00", 285=>x"b100", 286=>x"b100", 287=>x"b100", 288=>x"b000",
---- 289=>x"ac00", 290=>x"af00", 291=>x"b400", 292=>x"b200", 293=>x"ae00", 294=>x"a600", 295=>x"a700", 296=>x"b000", 297=>x"a200",
---- 298=>x"a500", 299=>x"a400", 300=>x"a100", 301=>x"a500", 302=>x"a900", 303=>x"a500", 304=>x"9500", 305=>x"8e00", 306=>x"9c00",
---- 307=>x"a300", 308=>x"9300", 309=>x"9100", 310=>x"9900", 311=>x"9a00", 312=>x"9e00", 313=>x"a100", 314=>x"9100", 315=>x"9600",
---- 316=>x"9800", 317=>x"9d00", 318=>x"9f00", 319=>x"9a00", 320=>x"9100", 321=>x"9700", 322=>x"9200", 323=>x"8c00", 324=>x"9e00",
---- 325=>x"8d00", 326=>x"9800", 327=>x"9300", 328=>x"9b00", 329=>x"9c00", 330=>x"8c00", 331=>x"8c00", 332=>x"9500", 333=>x"9400",
---- 334=>x"9700", 335=>x"8700", 336=>x"8c00", 337=>x"8c00", 338=>x"8e00", 339=>x"9000", 340=>x"9000", 341=>x"8c00", 342=>x"5b00",
---- 343=>x"6000", 344=>x"7400", 345=>x"9300", 346=>x"9200", 347=>x"8600", 348=>x"7a00", 349=>x"7700", 350=>x"8a00", 351=>x"9100",
---- 352=>x"8e00", 353=>x"8300", 354=>x"7d00", 355=>x"8400", 356=>x"8b00", 357=>x"8d00", 358=>x"8700", 359=>x"8200", 360=>x"8700",
---- 361=>x"8400", 362=>x"8600", 363=>x"8800", 364=>x"8d00", 365=>x"8300", 366=>x"8800", 367=>x"8e00", 368=>x"9100", 369=>x"9b00",
---- 370=>x"7900", 371=>x"8400", 372=>x"8c00", 373=>x"9300", 374=>x"9100", 375=>x"5800", 376=>x"6600", 377=>x"7700", 378=>x"7f00",
---- 379=>x"9400", 380=>x"8700", 381=>x"8c00", 382=>x"8800", 383=>x"8d00", 384=>x"9800", 385=>x"7e00", 386=>x"8400", 387=>x"8900",
---- 388=>x"8700", 389=>x"8800", 390=>x"7f00", 391=>x"8100", 392=>x"8700", 393=>x"8800", 394=>x"8c00", 395=>x"7b00", 396=>x"8300",
---- 397=>x"8c00", 398=>x"8e00", 399=>x"8500", 400=>x"7f00", 401=>x"8b00", 402=>x"8800", 403=>x"8c00", 404=>x"8900", 405=>x"8500",
---- 406=>x"8a00", 407=>x"8b00", 408=>x"8900", 409=>x"8a00", 410=>x"8400", 411=>x"8700", 412=>x"8d00", 413=>x"8900", 414=>x"8d00",
---- 415=>x"8700", 416=>x"8900", 417=>x"8500", 418=>x"8900", 419=>x"8e00", 420=>x"8800", 421=>x"8400", 422=>x"8800", 423=>x"8900",
---- 424=>x"8b00", 425=>x"8900", 426=>x"8900", 427=>x"8700", 428=>x"8a00", 429=>x"8600", 430=>x"8b00", 431=>x"8d00", 432=>x"8800",
---- 433=>x"8500", 434=>x"8a00", 435=>x"8b00", 436=>x"8b00", 437=>x"8b00", 438=>x"8500", 439=>x"8700", 440=>x"8b00", 441=>x"8d00",
---- 442=>x"8800", 443=>x"8700", 444=>x"8800", 445=>x"9000", 446=>x"8d00", 447=>x"8900", 448=>x"8400", 449=>x"8700", 450=>x"8f00",
---- 451=>x"8e00", 452=>x"8b00", 453=>x"8c00", 454=>x"8700", 455=>x"8f00", 456=>x"8b00", 457=>x"8e00", 458=>x"8500", 459=>x"8a00",
---- 460=>x"8a00", 461=>x"8f00", 462=>x"8e00", 463=>x"8d00", 464=>x"8700", 465=>x"8b00", 466=>x"8f00", 467=>x"8f00", 468=>x"8f00",
---- 469=>x"8700", 470=>x"8b00", 471=>x"8d00", 472=>x"8d00", 473=>x"8e00", 474=>x"8f00", 475=>x"8b00", 476=>x"8e00", 477=>x"8f00",
---- 478=>x"9000", 479=>x"8b00", 480=>x"8c00", 481=>x"8c00", 482=>x"8e00", 483=>x"8f00", 484=>x"9300", 485=>x"8c00", 486=>x"8d00",
---- 487=>x"8c00", 488=>x"8b00", 489=>x"8a00", 490=>x"8500", 491=>x"8900", 492=>x"8b00", 493=>x"8f00", 494=>x"9000", 495=>x"8900",
---- 496=>x"8800", 497=>x"8b00", 498=>x"8f00", 499=>x"9100"),
---- 11  => (0=>x"8000", 1=>x"8100", 2=>x"8000", 3=>x"7f00", 4=>x"7f00", 5=>x"7e00", 6=>x"8100", 7=>x"8000", 8=>x"7f00", 9=>x"7b00",
---- 10=>x"8000", 11=>x"7e00", 12=>x"8000", 13=>x"8000", 14=>x"7d00", 15=>x"7e00", 16=>x"8000", 17=>x"8100", 18=>x"7f00",
---- 19=>x"8000", 20=>x"7d00", 21=>x"7e00", 22=>x"7f00", 23=>x"7e00", 24=>x"7e00", 25=>x"7e00", 26=>x"7d00", 27=>x"7d00",
---- 28=>x"8000", 29=>x"7e00", 30=>x"7d00", 31=>x"7e00", 32=>x"7d00", 33=>x"7f00", 34=>x"7f00", 35=>x"7d00", 36=>x"7d00",
---- 37=>x"7e00", 38=>x"7d00", 39=>x"7e00", 40=>x"7e00", 41=>x"7f00", 42=>x"7e00", 43=>x"7e00", 44=>x"7c00", 45=>x"8000",
---- 46=>x"7d00", 47=>x"7e00", 48=>x"7f00", 49=>x"7e00", 50=>x"7f00", 51=>x"7f00", 52=>x"7d00", 53=>x"7c00", 54=>x"7a00",
---- 55=>x"7d00", 56=>x"7900", 57=>x"7c00", 58=>x"7a00", 59=>x"7700", 60=>x"6c00", 61=>x"7600", 62=>x"7900", 63=>x"7700",
---- 64=>x"7600", 65=>x"8d00", 66=>x"5e00", 67=>x"6a00", 68=>x"6f00", 69=>x"7300", 70=>x"cf00", 71=>x"9500", 72=>x"6800",
---- 73=>x"6500", 74=>x"6d00", 75=>x"d500", 76=>x"e400", 77=>x"ee00", 78=>x"6500", 79=>x"5f00", 80=>x"d400", 81=>x"d300",
---- 82=>x"e300", 83=>x"d600", 84=>x"5800", 85=>x"bd00", 86=>x"ba00", 87=>x"d400", 88=>x"e900", 89=>x"ab00", 90=>x"d000",
---- 91=>x"d700", 92=>x"ae00", 93=>x"dd00", 94=>x"ed00", 95=>x"c900", 96=>x"ca00", 97=>x"d400", 98=>x"d100", 99=>x"d600",
---- 100=>x"cf00", 101=>x"d000", 102=>x"ce00", 103=>x"d100", 104=>x"d000", 105=>x"ce00", 106=>x"cd00", 107=>x"cc00", 108=>x"cc00",
---- 109=>x"cb00", 110=>x"c900", 111=>x"ca00", 112=>x"c700", 113=>x"d000", 114=>x"d100", 115=>x"ce00", 116=>x"cc00", 117=>x"cf00",
---- 118=>x"ca00", 119=>x"c200", 120=>x"a500", 121=>x"ce00", 122=>x"a400", 123=>x"cb00", 124=>x"bf00", 125=>x"c300", 126=>x"c800",
---- 127=>x"cb00", 128=>x"c400", 129=>x"b400", 130=>x"c700", 131=>x"cb00", 132=>x"b100", 133=>x"b100", 134=>x"c900", 135=>x"9f00",
---- 136=>x"b400", 137=>x"b800", 138=>x"ba00", 139=>x"c000", 140=>x"b200", 141=>x"be00", 142=>x"b500", 143=>x"be00", 144=>x"c000",
---- 145=>x"b500", 146=>x"b300", 147=>x"a500", 148=>x"be00", 149=>x"b900", 150=>x"b300", 151=>x"b800", 152=>x"b900", 153=>x"b700",
---- 154=>x"af00", 155=>x"a800", 156=>x"b200", 157=>x"a800", 158=>x"a400", 159=>x"9500", 160=>x"a700", 161=>x"a300", 162=>x"a400",
---- 163=>x"9400", 164=>x"a200", 165=>x"9b00", 166=>x"a300", 167=>x"9e00", 168=>x"9000", 169=>x"af00", 170=>x"5d00", 171=>x"2d00",
---- 172=>x"9d00", 173=>x"b100", 174=>x"a600", 175=>x"1e00", 176=>x"4d00", 177=>x"aa00", 178=>x"a800", 179=>x"ce00", 180=>x"6f00",
---- 181=>x"9b00", 182=>x"ae00", 183=>x"c600", 184=>x"8900", 185=>x"9200", 186=>x"ac00", 187=>x"c100", 188=>x"b300", 189=>x"be00",
---- 190=>x"bb00", 191=>x"c200", 192=>x"b300", 193=>x"b800", 194=>x"ac00", 195=>x"c400", 196=>x"bc00", 197=>x"ab00", 198=>x"b600",
---- 199=>x"b200", 200=>x"be00", 201=>x"b600", 202=>x"a400", 203=>x"b600", 204=>x"9e00", 205=>x"b400", 206=>x"a900", 207=>x"b000",
---- 208=>x"af00", 209=>x"af00", 210=>x"9300", 211=>x"a800", 212=>x"b500", 213=>x"a100", 214=>x"ab00", 215=>x"9d00", 216=>x"b100",
---- 217=>x"a300", 218=>x"a100", 219=>x"b800", 220=>x"ab00", 221=>x"9c00", 222=>x"9f00", 223=>x"9700", 224=>x"c100", 225=>x"9900",
---- 226=>x"9f00", 227=>x"ab00", 228=>x"b400", 229=>x"a800", 230=>x"9f00", 231=>x"aa00", 232=>x"ad00", 233=>x"b200", 234=>x"be00",
---- 235=>x"ac00", 236=>x"b200", 237=>x"b300", 238=>x"b000", 239=>x"b600", 240=>x"6200", 241=>x"9700", 242=>x"b000", 243=>x"b300",
---- 244=>x"ad00", 245=>x"5a00", 246=>x"4400", 247=>x"7200", 248=>x"a800", 249=>x"a900", 250=>x"6000", 251=>x"8800", 252=>x"7b00",
---- 253=>x"8c00", 254=>x"9300", 255=>x"1f00", 256=>x"6e00", 257=>x"8000", 258=>x"8800", 259=>x"9800", 260=>x"5f00", 261=>x"6900",
---- 262=>x"7300", 263=>x"8300", 264=>x"8c00", 265=>x"8600", 266=>x"7b00", 267=>x"7900", 268=>x"7e00", 269=>x"9600", 270=>x"a300",
---- 271=>x"7d00", 272=>x"7f00", 273=>x"7d00", 274=>x"8f00", 275=>x"a200", 276=>x"8400", 277=>x"8800", 278=>x"7d00", 279=>x"8900",
---- 280=>x"9c00", 281=>x"8b00", 282=>x"8900", 283=>x"7f00", 284=>x"8400", 285=>x"9c00", 286=>x"9300", 287=>x"8b00", 288=>x"8200",
---- 289=>x"7b00", 290=>x"9800", 291=>x"9100", 292=>x"8d00", 293=>x"7e00", 294=>x"8400", 295=>x"9300", 296=>x"8500", 297=>x"8200",
---- 298=>x"7b00", 299=>x"8000", 300=>x"9100", 301=>x"8300", 302=>x"8100", 303=>x"7800", 304=>x"7b00", 305=>x"8a00", 306=>x"7500",
---- 307=>x"8600", 308=>x"7f00", 309=>x"7b00", 310=>x"8100", 311=>x"7500", 312=>x"8a00", 313=>x"8a00", 314=>x"7a00", 315=>x"8c00",
---- 316=>x"7c00", 317=>x"6400", 318=>x"5600", 319=>x"7400", 320=>x"9800", 321=>x"8c00", 322=>x"7f00", 323=>x"8b00", 324=>x"7f00",
---- 325=>x"9800", 326=>x"9400", 327=>x"8e00", 328=>x"aa00", 329=>x"b600", 330=>x"9200", 331=>x"9600", 332=>x"9900", 333=>x"c100",
---- 334=>x"c400", 335=>x"8f00", 336=>x"9200", 337=>x"9c00", 338=>x"a100", 339=>x"b700", 340=>x"7200", 341=>x"6800", 342=>x"5b00",
---- 343=>x"6800", 344=>x"7600", 345=>x"7c00", 346=>x"8900", 347=>x"a200", 348=>x"a600", 349=>x"c100", 350=>x"7e00", 351=>x"8200",
---- 352=>x"9100", 353=>x"9700", 354=>x"8d00", 355=>x"7e00", 356=>x"7800", 357=>x"7400", 358=>x"7600", 359=>x"8400", 360=>x"8f00",
---- 361=>x"9c00", 362=>x"a500", 363=>x"9500", 364=>x"9e00", 365=>x"a200", 366=>x"a700", 367=>x"a800", 368=>x"aa00", 369=>x"9c00",
---- 370=>x"a500", 371=>x"ab00", 372=>x"a900", 373=>x"aa00", 374=>x"9900", 375=>x"8e00", 376=>x"a700", 377=>x"7f00", 378=>x"9c00",
---- 379=>x"8c00", 380=>x"9d00", 381=>x"9900", 382=>x"9f00", 383=>x"a400", 384=>x"9c00", 385=>x"8e00", 386=>x"8c00", 387=>x"8b00",
---- 388=>x"9f00", 389=>x"ba00", 390=>x"8a00", 391=>x"8e00", 392=>x"9800", 393=>x"a900", 394=>x"bb00", 395=>x"8900", 396=>x"9300",
---- 397=>x"9f00", 398=>x"a900", 399=>x"ba00", 400=>x"8c00", 401=>x"9a00", 402=>x"a100", 403=>x"a600", 404=>x"9a00", 405=>x"8c00",
---- 406=>x"8d00", 407=>x"a100", 408=>x"a200", 409=>x"ac00", 410=>x"9200", 411=>x"9700", 412=>x"9c00", 413=>x"a000", 414=>x"a600",
---- 415=>x"9300", 416=>x"9200", 417=>x"9a00", 418=>x"9e00", 419=>x"a300", 420=>x"9100", 421=>x"9200", 422=>x"8c00", 423=>x"9b00",
---- 424=>x"a300", 425=>x"8f00", 426=>x"9100", 427=>x"9700", 428=>x"9c00", 429=>x"a100", 430=>x"8c00", 431=>x"8e00", 432=>x"9300",
---- 433=>x"9900", 434=>x"9e00", 435=>x"8b00", 436=>x"8e00", 437=>x"9200", 438=>x"9600", 439=>x"9a00", 440=>x"8900", 441=>x"8c00",
---- 442=>x"9200", 443=>x"8d00", 444=>x"9200", 445=>x"8900", 446=>x"8d00", 447=>x"9000", 448=>x"9400", 449=>x"9900", 450=>x"8700",
---- 451=>x"8c00", 452=>x"9000", 453=>x"9400", 454=>x"8e00", 455=>x"8600", 456=>x"8000", 457=>x"8d00", 458=>x"9000", 459=>x"9400",
---- 460=>x"8900", 461=>x"8700", 462=>x"8900", 463=>x"8700", 464=>x"9300", 465=>x"8600", 466=>x"8900", 467=>x"8b00", 468=>x"8a00",
---- 469=>x"8f00", 470=>x"8700", 471=>x"8600", 472=>x"8600", 473=>x"8500", 474=>x"8f00", 475=>x"9000", 476=>x"8e00", 477=>x"8b00",
---- 478=>x"8c00", 479=>x"8a00", 480=>x"9000", 481=>x"8f00", 482=>x"8b00", 483=>x"8d00", 484=>x"8d00", 485=>x"9200", 486=>x"8a00",
---- 487=>x"9300", 488=>x"8e00", 489=>x"8e00", 490=>x"9300", 491=>x"9200", 492=>x"8f00", 493=>x"8a00", 494=>x"9500", 495=>x"8f00",
---- 496=>x"9100", 497=>x"9200", 498=>x"9100", 499=>x"9500"),
---- 12  => (0=>x"7900", 1=>x"7100", 2=>x"6600", 3=>x"7d00", 4=>x"9200", 5=>x"7800", 6=>x"7000", 7=>x"6600", 8=>x"7600", 9=>x"8d00",
---- 10=>x"7900", 11=>x"7100", 12=>x"6c00", 13=>x"6c00", 14=>x"8200", 15=>x"7a00", 16=>x"7200", 17=>x"7100", 18=>x"6600",
---- 19=>x"7400", 20=>x"7a00", 21=>x"7800", 22=>x"6e00", 23=>x"6900", 24=>x"6d00", 25=>x"7a00", 26=>x"7a00", 27=>x"6f00",
---- 28=>x"6a00", 29=>x"7100", 30=>x"7b00", 31=>x"7500", 32=>x"7700", 33=>x"6b00", 34=>x"7100", 35=>x"7a00", 36=>x"7900",
---- 37=>x"7300", 38=>x"6c00", 39=>x"6f00", 40=>x"7a00", 41=>x"7500", 42=>x"7800", 43=>x"6d00", 44=>x"6f00", 45=>x"7900",
---- 46=>x"7400", 47=>x"7200", 48=>x"6f00", 49=>x"6d00", 50=>x"7900", 51=>x"7800", 52=>x"7100", 53=>x"6d00", 54=>x"6c00",
---- 55=>x"7300", 56=>x"7000", 57=>x"6e00", 58=>x"6900", 59=>x"6e00", 60=>x"7300", 61=>x"7600", 62=>x"6d00", 63=>x"6500",
---- 64=>x"6a00", 65=>x"7600", 66=>x"6c00", 67=>x"7200", 68=>x"6400", 69=>x"6800", 70=>x"6d00", 71=>x"6a00", 72=>x"6900",
---- 73=>x"7900", 74=>x"6f00", 75=>x"7700", 76=>x"6300", 77=>x"6900", 78=>x"6a00", 79=>x"6500", 80=>x"5b00", 81=>x"6400",
---- 82=>x"6300", 83=>x"5e00", 84=>x"6200", 85=>x"4100", 86=>x"5b00", 87=>x"6400", 88=>x"6700", 89=>x"6d00", 90=>x"7e00",
---- 91=>x"3e00", 92=>x"5100", 93=>x"5700", 94=>x"5f00", 95=>x"e800", 96=>x"ad00", 97=>x"3f00", 98=>x"4e00", 99=>x"5c00",
---- 100=>x"d500", 101=>x"ea00", 102=>x"a100", 103=>x"2d00", 104=>x"5700", 105=>x"d500", 106=>x"db00", 107=>x"ef00", 108=>x"6500",
---- 109=>x"4500", 110=>x"cf00", 111=>x"d700", 112=>x"af00", 113=>x"b000", 114=>x"3000", 115=>x"cf00", 116=>x"cc00", 117=>x"d900",
---- 118=>x"f000", 119=>x"6800", 120=>x"d000", 121=>x"ce00", 122=>x"cd00", 123=>x"dc00", 124=>x"c400", 125=>x"ba00", 126=>x"cc00",
---- 127=>x"cc00", 128=>x"ce00", 129=>x"dd00", 130=>x"cb00", 131=>x"c900", 132=>x"c900", 133=>x"c400", 134=>x"ca00", 135=>x"c300",
---- 136=>x"c400", 137=>x"c200", 138=>x"c700", 139=>x"be00", 140=>x"c000", 141=>x"ba00", 142=>x"bd00", 143=>x"a200", 144=>x"b600",
---- 145=>x"b200", 146=>x"ac00", 147=>x"bb00", 148=>x"a600", 149=>x"a500", 150=>x"b800", 151=>x"ac00", 152=>x"a700", 153=>x"a400",
---- 154=>x"b800", 155=>x"b200", 156=>x"9900", 157=>x"a800", 158=>x"ba00", 159=>x"b700", 160=>x"7f00", 161=>x"bb00", 162=>x"b300",
---- 163=>x"bf00", 164=>x"c800", 165=>x"b800", 166=>x"b500", 167=>x"c700", 168=>x"c700", 169=>x"ba00", 170=>x"ba00", 171=>x"cf00",
---- 172=>x"a300", 173=>x"c500", 174=>x"c100", 175=>x"c600", 176=>x"c300", 177=>x"c600", 178=>x"c400", 179=>x"be00", 180=>x"c900",
---- 181=>x"ae00", 182=>x"a000", 183=>x"b500", 184=>x"c100", 185=>x"bb00", 186=>x"b500", 187=>x"b700", 188=>x"ba00", 189=>x"bf00",
---- 190=>x"ae00", 191=>x"b800", 192=>x"a800", 193=>x"c000", 194=>x"c200", 195=>x"b100", 196=>x"b200", 197=>x"c100", 198=>x"c000",
---- 199=>x"b800", 200=>x"ac00", 201=>x"a200", 202=>x"ba00", 203=>x"b900", 204=>x"c500", 205=>x"ac00", 206=>x"be00", 207=>x"b700",
---- 208=>x"a500", 209=>x"ca00", 210=>x"bd00", 211=>x"c800", 212=>x"c500", 213=>x"be00", 214=>x"c800", 215=>x"c400", 216=>x"aa00",
---- 217=>x"c400", 218=>x"b300", 219=>x"d500", 220=>x"c500", 221=>x"ca00", 222=>x"c900", 223=>x"d300", 224=>x"ac00", 225=>x"af00",
---- 226=>x"ca00", 227=>x"cc00", 228=>x"ce00", 229=>x"d500", 230=>x"bf00", 231=>x"c700", 232=>x"c800", 233=>x"cc00", 234=>x"d100",
---- 235=>x"c100", 236=>x"c400", 237=>x"c600", 238=>x"c800", 239=>x"cc00", 240=>x"bb00", 241=>x"c300", 242=>x"a100", 243=>x"c600",
---- 244=>x"cd00", 245=>x"b700", 246=>x"c000", 247=>x"c000", 248=>x"be00", 249=>x"9800", 250=>x"b000", 251=>x"c600", 252=>x"ca00",
---- 253=>x"9a00", 254=>x"5400", 255=>x"b700", 256=>x"dc00", 257=>x"a000", 258=>x"2300", 259=>x"2e00", 260=>x"c200", 261=>x"da00",
---- 262=>x"5700", 263=>x"4500", 264=>x"4000", 265=>x"d300", 266=>x"c200", 267=>x"6400", 268=>x"7e00", 269=>x"7800", 270=>x"cc00",
---- 271=>x"d000", 272=>x"9a00", 273=>x"8800", 274=>x"8400", 275=>x"ba00", 276=>x"d900", 277=>x"ac00", 278=>x"9700", 279=>x"8800",
---- 280=>x"a900", 281=>x"de00", 282=>x"af00", 283=>x"9300", 284=>x"9100", 285=>x"b400", 286=>x"e200", 287=>x"b100", 288=>x"a400",
---- 289=>x"9100", 290=>x"ae00", 291=>x"e500", 292=>x"b100", 293=>x"a100", 294=>x"9500", 295=>x"9f00", 296=>x"e100", 297=>x"b400",
---- 298=>x"9c00", 299=>x"9400", 300=>x"9b00", 301=>x"da00", 302=>x"c500", 303=>x"9900", 304=>x"9200", 305=>x"9400", 306=>x"d500",
---- 307=>x"a500", 308=>x"8900", 309=>x"9400", 310=>x"8a00", 311=>x"cc00", 312=>x"cb00", 313=>x"8600", 314=>x"8e00", 315=>x"6d00",
---- 316=>x"b000", 317=>x"a800", 318=>x"9200", 319=>x"8c00", 320=>x"ab00", 321=>x"be00", 322=>x"a000", 323=>x"9300", 324=>x"8700",
---- 325=>x"c300", 326=>x"c100", 327=>x"9c00", 328=>x"8f00", 329=>x"8a00", 330=>x"c600", 331=>x"c400", 332=>x"9600", 333=>x"8f00",
---- 334=>x"7c00", 335=>x"b500", 336=>x"af00", 337=>x"8300", 338=>x"9100", 339=>x"4c00", 340=>x"5d00", 341=>x"6800", 342=>x"7900",
---- 343=>x"8c00", 344=>x"2100", 345=>x"9800", 346=>x"8d00", 347=>x"9700", 348=>x"5c00", 349=>x"2600", 350=>x"8b00", 351=>x"9900",
---- 352=>x"7a00", 353=>x"2100", 354=>x"2f00", 355=>x"9600", 356=>x"8b00", 357=>x"3c00", 358=>x"2700", 359=>x"2c00", 360=>x"9400",
---- 361=>x"7500", 362=>x"3d00", 363=>x"2900", 364=>x"3100", 365=>x"9200", 366=>x"2c00", 367=>x"3500", 368=>x"2e00", 369=>x"3a00",
---- 370=>x"8500", 371=>x"2700", 372=>x"3700", 373=>x"3800", 374=>x"3b00", 375=>x"6d00", 376=>x"1f00", 377=>x"3300", 378=>x"3700",
---- 379=>x"3700", 380=>x"c400", 381=>x"aa00", 382=>x"5700", 383=>x"2900", 384=>x"2d00", 385=>x"c500", 386=>x"ce00", 387=>x"da00",
---- 388=>x"bc00", 389=>x"5f00", 390=>x"c000", 391=>x"c500", 392=>x"cb00", 393=>x"ad00", 394=>x"e000", 395=>x"b900", 396=>x"a700",
---- 397=>x"c300", 398=>x"ce00", 399=>x"cf00", 400=>x"b600", 401=>x"bb00", 402=>x"c200", 403=>x"a700", 404=>x"aa00", 405=>x"ae00",
---- 406=>x"b400", 407=>x"b800", 408=>x"c500", 409=>x"cd00", 410=>x"ab00", 411=>x"b200", 412=>x"b700", 413=>x"bf00", 414=>x"c500",
---- 415=>x"ab00", 416=>x"b100", 417=>x"b800", 418=>x"bb00", 419=>x"c400", 420=>x"a900", 421=>x"9e00", 422=>x"af00", 423=>x"bc00",
---- 424=>x"c300", 425=>x"9300", 426=>x"af00", 427=>x"b300", 428=>x"b900", 429=>x"c300", 430=>x"9800", 431=>x"aa00", 432=>x"ac00",
---- 433=>x"ae00", 434=>x"ad00", 435=>x"9b00", 436=>x"a900", 437=>x"9700", 438=>x"b800", 439=>x"b800", 440=>x"a000", 441=>x"a500",
---- 442=>x"a900", 443=>x"b200", 444=>x"bd00", 445=>x"9a00", 446=>x"9e00", 447=>x"a600", 448=>x"af00", 449=>x"b700", 450=>x"9a00",
---- 451=>x"a200", 452=>x"a500", 453=>x"a900", 454=>x"b300", 455=>x"9700", 456=>x"8900", 457=>x"a100", 458=>x"a900", 459=>x"ad00",
---- 460=>x"9800", 461=>x"9100", 462=>x"a000", 463=>x"a300", 464=>x"af00", 465=>x"9300", 466=>x"9000", 467=>x"9400", 468=>x"a200",
---- 469=>x"a900", 470=>x"9100", 471=>x"9600", 472=>x"9600", 473=>x"a300", 474=>x"a400", 475=>x"9000", 476=>x"9300", 477=>x"9a00",
---- 478=>x"8f00", 479=>x"a500", 480=>x"8d00", 481=>x"9300", 482=>x"9700", 483=>x"9e00", 484=>x"a000", 485=>x"9100", 486=>x"9300",
---- 487=>x"8b00", 488=>x"9a00", 489=>x"9f00", 490=>x"9100", 491=>x"9500", 492=>x"9700", 493=>x"9900", 494=>x"a200", 495=>x"9300",
---- 496=>x"9600", 497=>x"9600", 498=>x"9400", 499=>x"9200"),
---- 13  => (0=>x"9b00", 1=>x"a100", 2=>x"9600", 3=>x"9800", 4=>x"9b00", 5=>x"9900", 6=>x"a100", 7=>x"9900", 8=>x"9700", 9=>x"9900",
---- 10=>x"9400", 11=>x"a000", 12=>x"9e00", 13=>x"9a00", 14=>x"9e00", 15=>x"9100", 16=>x"8a00", 17=>x"a400", 18=>x"a200",
---- 19=>x"a000", 20=>x"8a00", 21=>x"8d00", 22=>x"9100", 23=>x"a400", 24=>x"a100", 25=>x"8500", 26=>x"9900", 27=>x"9e00",
---- 28=>x"a200", 29=>x"a100", 30=>x"8400", 31=>x"9300", 32=>x"9c00", 33=>x"a000", 34=>x"a000", 35=>x"8200", 36=>x"8e00",
---- 37=>x"9800", 38=>x"9300", 39=>x"9900", 40=>x"7e00", 41=>x"8d00", 42=>x"9300", 43=>x"9900", 44=>x"9a00", 45=>x"7d00",
---- 46=>x"8e00", 47=>x"8b00", 48=>x"9200", 49=>x"9600", 50=>x"7f00", 51=>x"8e00", 52=>x"8e00", 53=>x"9000", 54=>x"9300",
---- 55=>x"7f00", 56=>x"8f00", 57=>x"9200", 58=>x"8f00", 59=>x"9300", 60=>x"8000", 61=>x"8a00", 62=>x"9500", 63=>x"9000",
---- 64=>x"9100", 65=>x"7f00", 66=>x"9300", 67=>x"9800", 68=>x"9400", 69=>x"9000", 70=>x"7e00", 71=>x"9600", 72=>x"9a00",
---- 73=>x"9a00", 74=>x"9400", 75=>x"7f00", 76=>x"9600", 77=>x"9c00", 78=>x"9c00", 79=>x"9900", 80=>x"7d00", 81=>x"9300",
---- 82=>x"9b00", 83=>x"9100", 84=>x"9600", 85=>x"7a00", 86=>x"9400", 87=>x"9c00", 88=>x"9a00", 89=>x"9900", 90=>x"7e00",
---- 91=>x"9400", 92=>x"9c00", 93=>x"9a00", 94=>x"9b00", 95=>x"7d00", 96=>x"9400", 97=>x"9b00", 98=>x"9900", 99=>x"9a00",
---- 100=>x"7b00", 101=>x"9300", 102=>x"9a00", 103=>x"9900", 104=>x"9b00", 105=>x"7600", 106=>x"9200", 107=>x"9a00", 108=>x"9800",
---- 109=>x"9900", 110=>x"7600", 111=>x"9300", 112=>x"8e00", 113=>x"9500", 114=>x"9800", 115=>x"6400", 116=>x"9300", 117=>x"9a00",
---- 118=>x"9a00", 119=>x"9b00", 120=>x"5200", 121=>x"9000", 122=>x"9d00", 123=>x"9d00", 124=>x"9c00", 125=>x"ac00", 126=>x"8200",
---- 127=>x"9800", 128=>x"9b00", 129=>x"9a00", 130=>x"de00", 131=>x"b000", 132=>x"9400", 133=>x"9600", 134=>x"8e00", 135=>x"c000",
---- 136=>x"cd00", 137=>x"9000", 138=>x"9000", 139=>x"b300", 140=>x"b800", 141=>x"be00", 142=>x"b300", 143=>x"cd00", 144=>x"bf00",
---- 145=>x"aa00", 146=>x"c100", 147=>x"bb00", 148=>x"c100", 149=>x"cb00", 150=>x"c000", 151=>x"ba00", 152=>x"c700", 153=>x"cd00",
---- 154=>x"c600", 155=>x"c600", 156=>x"ce00", 157=>x"c700", 158=>x"bf00", 159=>x"bf00", 160=>x"c300", 161=>x"bc00", 162=>x"be00",
---- 163=>x"c600", 164=>x"a500", 165=>x"ba00", 166=>x"c100", 167=>x"c400", 168=>x"c600", 169=>x"cc00", 170=>x"c000", 171=>x"c500",
---- 172=>x"c800", 173=>x"c900", 174=>x"cd00", 175=>x"c200", 176=>x"c600", 177=>x"c800", 178=>x"c400", 179=>x"ce00", 180=>x"c100",
---- 181=>x"c300", 182=>x"c800", 183=>x"d300", 184=>x"d000", 185=>x"c200", 186=>x"ce00", 187=>x"cb00", 188=>x"8400", 189=>x"6e00",
---- 190=>x"d400", 191=>x"8600", 192=>x"5b00", 193=>x"6700", 194=>x"6900", 195=>x"6d00", 196=>x"3600", 197=>x"5c00", 198=>x"7400",
---- 199=>x"7700", 200=>x"a700", 201=>x"5900", 202=>x"6700", 203=>x"6200", 204=>x"8400", 205=>x"c800", 206=>x"6900", 207=>x"4100",
---- 208=>x"5800", 209=>x"5800", 210=>x"c600", 211=>x"8d00", 212=>x"4700", 213=>x"3e00", 214=>x"8a00", 215=>x"d100", 216=>x"a300",
---- 217=>x"5600", 218=>x"1d00", 219=>x"3a00", 220=>x"d800", 221=>x"ba00", 222=>x"6700", 223=>x"2a00", 224=>x"2800", 225=>x"d700",
---- 226=>x"c800", 227=>x"7700", 228=>x"3200", 229=>x"2100", 230=>x"d600", 231=>x"d500", 232=>x"8d00", 233=>x"5d00", 234=>x"2000",
---- 235=>x"d800", 236=>x"b300", 237=>x"a300", 238=>x"5e00", 239=>x"2600", 240=>x"ca00", 241=>x"9c00", 242=>x"6400", 243=>x"3100",
---- 244=>x"2300", 245=>x"6400", 246=>x"6a00", 247=>x"7600", 248=>x"5800", 249=>x"3100", 250=>x"3600", 251=>x"2800", 252=>x"3700",
---- 253=>x"3f00", 254=>x"3000", 255=>x"7400", 256=>x"4900", 257=>x"2b00", 258=>x"5200", 259=>x"2b00", 260=>x"8600", 261=>x"8400",
---- 262=>x"2600", 263=>x"4800", 264=>x"2700", 265=>x"a700", 266=>x"6800", 267=>x"5200", 268=>x"6100", 269=>x"3700", 270=>x"6000",
---- 271=>x"4200", 272=>x"5200", 273=>x"2f00", 274=>x"2b00", 275=>x"7a00", 276=>x"6d00", 277=>x"6700", 278=>x"3800", 279=>x"2900",
---- 280=>x"8400", 281=>x"7b00", 282=>x"7000", 283=>x"3600", 284=>x"5600", 285=>x"8400", 286=>x"8100", 287=>x"7700", 288=>x"3500",
---- 289=>x"3500", 290=>x"8900", 291=>x"8100", 292=>x"6f00", 293=>x"3100", 294=>x"3300", 295=>x"8a00", 296=>x"8200", 297=>x"6200",
---- 298=>x"2900", 299=>x"3400", 300=>x"8700", 301=>x"8200", 302=>x"4f00", 303=>x"2700", 304=>x"3d00", 305=>x"8300", 306=>x"7d00",
---- 307=>x"3600", 308=>x"2800", 309=>x"4000", 310=>x"8400", 311=>x"6300", 312=>x"2100", 313=>x"5000", 314=>x"3a00", 315=>x"8400",
---- 316=>x"7000", 317=>x"2400", 318=>x"3e00", 319=>x"6500", 320=>x"7200", 321=>x"2c00", 322=>x"2d00", 323=>x"3600", 324=>x"4f00",
---- 325=>x"4500", 326=>x"2b00", 327=>x"2d00", 328=>x"3d00", 329=>x"5000", 330=>x"2400", 331=>x"4100", 332=>x"2c00", 333=>x"4d00",
---- 334=>x"4c00", 335=>x"2300", 336=>x"4400", 337=>x"2e00", 338=>x"5f00", 339=>x"5500", 340=>x"5600", 341=>x"2900", 342=>x"3600",
---- 343=>x"4100", 344=>x"4a00", 345=>x"3100", 346=>x"2b00", 347=>x"3a00", 348=>x"4000", 349=>x"4e00", 350=>x"3200", 351=>x"2d00",
---- 352=>x"3600", 353=>x"4200", 354=>x"4e00", 355=>x"3500", 356=>x"3900", 357=>x"3300", 358=>x"4900", 359=>x"4e00", 360=>x"3a00",
---- 361=>x"3700", 362=>x"2d00", 363=>x"4c00", 364=>x"4f00", 365=>x"4300", 366=>x"4100", 367=>x"3c00", 368=>x"5600", 369=>x"5400",
---- 370=>x"4600", 371=>x"4200", 372=>x"4000", 373=>x"5b00", 374=>x"5300", 375=>x"3d00", 376=>x"3000", 377=>x"3000", 378=>x"5c00",
---- 379=>x"5800", 380=>x"3400", 381=>x"5500", 382=>x"3200", 383=>x"5a00", 384=>x"5700", 385=>x"2500", 386=>x"2200", 387=>x"2f00",
---- 388=>x"6000", 389=>x"5200", 390=>x"b700", 391=>x"3000", 392=>x"2100", 393=>x"5b00", 394=>x"5300", 395=>x"db00", 396=>x"b200",
---- 397=>x"4f00", 398=>x"5200", 399=>x"4400", 400=>x"d500", 401=>x"da00", 402=>x"e700", 403=>x"5300", 404=>x"3b00", 405=>x"ae00",
---- 406=>x"d800", 407=>x"b800", 408=>x"d900", 409=>x"2800", 410=>x"cb00", 411=>x"cf00", 412=>x"d600", 413=>x"d700", 414=>x"9d00",
---- 415=>x"cc00", 416=>x"d100", 417=>x"d600", 418=>x"c700", 419=>x"eb00", 420=>x"cb00", 421=>x"d000", 422=>x"d300", 423=>x"d800",
---- 424=>x"e900", 425=>x"c800", 426=>x"d000", 427=>x"d100", 428=>x"d800", 429=>x"de00", 430=>x"c900", 431=>x"ce00", 432=>x"d000",
---- 433=>x"b000", 434=>x"db00", 435=>x"c500", 436=>x"cb00", 437=>x"d000", 438=>x"d600", 439=>x"d500", 440=>x"c400", 441=>x"cb00",
---- 442=>x"d000", 443=>x"d300", 444=>x"d400", 445=>x"c300", 446=>x"ab00", 447=>x"ac00", 448=>x"b300", 449=>x"da00", 450=>x"bf00",
---- 451=>x"b500", 452=>x"c000", 453=>x"d900", 454=>x"af00", 455=>x"ba00", 456=>x"c500", 457=>x"cd00", 458=>x"cf00", 459=>x"d400",
---- 460=>x"b600", 461=>x"b200", 462=>x"b900", 463=>x"cf00", 464=>x"d000", 465=>x"b300", 466=>x"a200", 467=>x"ca00", 468=>x"b600",
---- 469=>x"c600", 470=>x"ad00", 471=>x"b800", 472=>x"bf00", 473=>x"c900", 474=>x"cf00", 475=>x"a900", 476=>x"b100", 477=>x"bb00",
---- 478=>x"c400", 479=>x"ca00", 480=>x"a900", 481=>x"b200", 482=>x"b900", 483=>x"bf00", 484=>x"c800", 485=>x"a600", 486=>x"ac00",
---- 487=>x"b300", 488=>x"bb00", 489=>x"c200", 490=>x"a600", 491=>x"ab00", 492=>x"b500", 493=>x"ae00", 494=>x"c000", 495=>x"a500",
---- 496=>x"a800", 497=>x"9b00", 498=>x"ab00", 499=>x"c000"),
---- 14  => (0=>x"9d00", 1=>x"9900", 2=>x"9900", 3=>x"9800", 4=>x"9a00", 5=>x"9900", 6=>x"9a00", 7=>x"8e00", 8=>x"9900", 9=>x"9900",
---- 10=>x"a000", 11=>x"9200", 12=>x"9d00", 13=>x"9c00", 14=>x"9000", 15=>x"a300", 16=>x"a200", 17=>x"9d00", 18=>x"9e00",
---- 19=>x"9b00", 20=>x"a100", 21=>x"a100", 22=>x"9e00", 23=>x"9b00", 24=>x"9b00", 25=>x"9d00", 26=>x"9e00", 27=>x"9f00",
---- 28=>x"9b00", 29=>x"9c00", 30=>x"9d00", 31=>x"9f00", 32=>x"9e00", 33=>x"9c00", 34=>x"9c00", 35=>x"9e00", 36=>x"9c00",
---- 37=>x"9c00", 38=>x"9c00", 39=>x"9a00", 40=>x"9c00", 41=>x"9a00", 42=>x"9a00", 43=>x"9b00", 44=>x"9900", 45=>x"9a00",
---- 46=>x"9a00", 47=>x"9900", 48=>x"8900", 49=>x"9500", 50=>x"9800", 51=>x"9900", 52=>x"9800", 53=>x"9a00", 54=>x"9600",
---- 55=>x"9400", 56=>x"9800", 57=>x"9900", 58=>x"8900", 59=>x"9300", 60=>x"9200", 61=>x"9300", 62=>x"9700", 63=>x"9700",
---- 64=>x"8d00", 65=>x"8e00", 66=>x"8c00", 67=>x"8c00", 68=>x"9700", 69=>x"9000", 70=>x"8700", 71=>x"8000", 72=>x"8000",
---- 73=>x"9200", 74=>x"8900", 75=>x"8900", 76=>x"6d00", 77=>x"6b00", 78=>x"8700", 79=>x"9100", 80=>x"8e00", 81=>x"6500",
---- 82=>x"4100", 83=>x"6d00", 84=>x"8f00", 85=>x"9100", 86=>x"6e00", 87=>x"2900", 88=>x"5e00", 89=>x"7d00", 90=>x"9300",
---- 91=>x"7200", 92=>x"2b00", 93=>x"3300", 94=>x"6c00", 95=>x"9500", 96=>x"6f00", 97=>x"3000", 98=>x"2900", 99=>x"4800",
---- 100=>x"9200", 101=>x"7100", 102=>x"3500", 103=>x"2600", 104=>x"2700", 105=>x"8f00", 106=>x"7100", 107=>x"4000", 108=>x"2b00",
---- 109=>x"2400", 110=>x"9000", 111=>x"7200", 112=>x"4c00", 113=>x"2a00", 114=>x"2700", 115=>x"9400", 116=>x"7000", 117=>x"3000",
---- 118=>x"1d00", 119=>x"1800", 120=>x"9300", 121=>x"6700", 122=>x"3b00", 123=>x"4e00", 124=>x"c200", 125=>x"8800", 126=>x"4500",
---- 127=>x"6300", 128=>x"da00", 129=>x"bc00", 130=>x"7600", 131=>x"bc00", 132=>x"d200", 133=>x"bb00", 134=>x"d500", 135=>x"d600",
---- 136=>x"bc00", 137=>x"c500", 138=>x"d300", 139=>x"cb00", 140=>x"c100", 141=>x"d100", 142=>x"cf00", 143=>x"c900", 144=>x"c900",
---- 145=>x"d500", 146=>x"a700", 147=>x"ca00", 148=>x"c800", 149=>x"a900", 150=>x"c600", 151=>x"a900", 152=>x"c900", 153=>x"cc00",
---- 154=>x"ac00", 155=>x"c300", 156=>x"cb00", 157=>x"ca00", 158=>x"bc00", 159=>x"c100", 160=>x"cc00", 161=>x"cc00", 162=>x"bc00",
---- 163=>x"cd00", 164=>x"d900", 165=>x"cd00", 166=>x"cc00", 167=>x"bc00", 168=>x"d500", 169=>x"c800", 170=>x"b300", 171=>x"c700",
---- 172=>x"db00", 173=>x"d200", 174=>x"9300", 175=>x"da00", 176=>x"c600", 177=>x"8a00", 178=>x"5e00", 179=>x"4d00", 180=>x"7b00",
---- 181=>x"4b00", 182=>x"4800", 183=>x"6300", 184=>x"6e00", 185=>x"7b00", 186=>x"6800", 187=>x"7f00", 188=>x"9d00", 189=>x"aa00",
---- 190=>x"9e00", 191=>x"ab00", 192=>x"ab00", 193=>x"aa00", 194=>x"d300", 195=>x"8400", 196=>x"a300", 197=>x"b100", 198=>x"ce00",
---- 199=>x"6a00", 200=>x"7b00", 201=>x"b200", 202=>x"a800", 203=>x"4400", 204=>x"1e00", 205=>x"8d00", 206=>x"9b00", 207=>x"4400",
---- 208=>x"2000", 209=>x"2c00", 210=>x"8100", 211=>x"9a00", 212=>x"3f00", 213=>x"2800", 214=>x"2900", 215=>x"7e00", 216=>x"a500",
---- 217=>x"2900", 218=>x"2d00", 219=>x"3100", 220=>x"5e00", 221=>x"ab00", 222=>x"3500", 223=>x"3100", 224=>x"3400", 225=>x"4f00",
---- 226=>x"a500", 227=>x"5600", 228=>x"2e00", 229=>x"3800", 230=>x"3400", 231=>x"a800", 232=>x"6300", 233=>x"2b00", 234=>x"3900",
---- 235=>x"4b00", 236=>x"9a00", 237=>x"5a00", 238=>x"3900", 239=>x"3c00", 240=>x"2b00", 241=>x"8400", 242=>x"7500", 243=>x"3300",
---- 244=>x"3c00", 245=>x"2800", 246=>x"7600", 247=>x"8700", 248=>x"3500", 249=>x"4d00", 250=>x"2900", 251=>x"6f00", 252=>x"8f00",
---- 253=>x"3f00", 254=>x"5100", 255=>x"2a00", 256=>x"6400", 257=>x"9000", 258=>x"3d00", 259=>x"4200", 260=>x"3700", 261=>x"5b00",
---- 262=>x"9500", 263=>x"5b00", 264=>x"3e00", 265=>x"3c00", 266=>x"5000", 267=>x"a200", 268=>x"5500", 269=>x"3d00", 270=>x"5100",
---- 271=>x"4a00", 272=>x"ad00", 273=>x"4e00", 274=>x"3900", 275=>x"4100", 276=>x"4300", 277=>x"b800", 278=>x"4b00", 279=>x"3500",
---- 280=>x"3c00", 281=>x"3500", 282=>x"c000", 283=>x"5200", 284=>x"2f00", 285=>x"4e00", 286=>x"2d00", 287=>x"b400", 288=>x"5e00",
---- 289=>x"2600", 290=>x"5300", 291=>x"2500", 292=>x"a900", 293=>x"7600", 294=>x"1d00", 295=>x"4800", 296=>x"2000", 297=>x"8c00",
---- 298=>x"8800", 299=>x"2100", 300=>x"4b00", 301=>x"1b00", 302=>x"9900", 303=>x"9200", 304=>x"2300", 305=>x"4700", 306=>x"1a00",
---- 307=>x"8600", 308=>x"9c00", 309=>x"3400", 310=>x"4800", 311=>x"1e00", 312=>x"7000", 313=>x"a700", 314=>x"4500", 315=>x"4e00",
---- 316=>x"2500", 317=>x"5300", 318=>x"a700", 319=>x"4c00", 320=>x"3f00", 321=>x"3900", 322=>x"5900", 323=>x"a600", 324=>x"5800",
---- 325=>x"4300", 326=>x"3600", 327=>x"2700", 328=>x"a900", 329=>x"5d00", 330=>x"4100", 331=>x"3200", 332=>x"2f00", 333=>x"a000",
---- 334=>x"6400", 335=>x"4600", 336=>x"3800", 337=>x"2700", 338=>x"9a00", 339=>x"6f00", 340=>x"4300", 341=>x"3f00", 342=>x"1a00",
---- 343=>x"8500", 344=>x"8400", 345=>x"4100", 346=>x"4900", 347=>x"2600", 348=>x"7800", 349=>x"9500", 350=>x"4800", 351=>x"4600",
---- 352=>x"4700", 353=>x"7200", 354=>x"9e00", 355=>x"4a00", 356=>x"4600", 357=>x"2b00", 358=>x"6f00", 359=>x"9f00", 360=>x"4b00",
---- 361=>x"4b00", 362=>x"3200", 363=>x"6700", 364=>x"a300", 365=>x"4a00", 366=>x"5200", 367=>x"3900", 368=>x"6400", 369=>x"ad00",
---- 370=>x"5b00", 371=>x"5b00", 372=>x"3f00", 373=>x"6100", 374=>x"ac00", 375=>x"5600", 376=>x"6900", 377=>x"4000", 378=>x"6e00",
---- 379=>x"a700", 380=>x"5800", 381=>x"5500", 382=>x"4000", 383=>x"7900", 384=>x"9b00", 385=>x"4e00", 386=>x"5100", 387=>x"3e00",
---- 388=>x"9700", 389=>x"8400", 390=>x"4900", 391=>x"6200", 392=>x"3600", 393=>x"9800", 394=>x"8800", 395=>x"4200", 396=>x"5000",
---- 397=>x"3b00", 398=>x"9300", 399=>x"8d00", 400=>x"3d00", 401=>x"4c00", 402=>x"2e00", 403=>x"9100", 404=>x"8e00", 405=>x"3200",
---- 406=>x"4500", 407=>x"4300", 408=>x"9d00", 409=>x"8e00", 410=>x"1f00", 411=>x"2f00", 412=>x"3700", 413=>x"9900", 414=>x"9100",
---- 415=>x"2c00", 416=>x"1f00", 417=>x"4400", 418=>x"9c00", 419=>x"8a00", 420=>x"8600", 421=>x"a00", 422=>x"5500", 423=>x"9600",
---- 424=>x"9600", 425=>x"c700", 426=>x"3200", 427=>x"5f00", 428=>x"9500", 429=>x"9600", 430=>x"ed00", 431=>x"1f00", 432=>x"6a00",
---- 433=>x"9300", 434=>x"8e00", 435=>x"e700", 436=>x"6000", 437=>x"7000", 438=>x"9300", 439=>x"9400", 440=>x"db00", 441=>x"a700",
---- 442=>x"6f00", 443=>x"9300", 444=>x"9500", 445=>x"d500", 446=>x"d500", 447=>x"8900", 448=>x"6d00", 449=>x"7400", 450=>x"d900",
---- 451=>x"e300", 452=>x"8200", 453=>x"4300", 454=>x"4900", 455=>x"d400", 456=>x"e100", 457=>x"9b00", 458=>x"4b00", 459=>x"5400",
---- 460=>x"d400", 461=>x"de00", 462=>x"cd00", 463=>x"4a00", 464=>x"6800", 465=>x"d600", 466=>x"ae00", 467=>x"e900", 468=>x"5900",
---- 469=>x"6300", 470=>x"d200", 471=>x"d800", 472=>x"e400", 473=>x"8700", 474=>x"5500", 475=>x"d100", 476=>x"c900", 477=>x"c100",
---- 478=>x"b800", 479=>x"4a00", 480=>x"cd00", 481=>x"d400", 482=>x"d900", 483=>x"d600", 484=>x"4d00", 485=>x"c900", 486=>x"d100",
---- 487=>x"d200", 488=>x"e000", 489=>x"6100", 490=>x"c800", 491=>x"cc00", 492=>x"d100", 493=>x"dd00", 494=>x"9100", 495=>x"c400",
---- 496=>x"ca00", 497=>x"cf00", 498=>x"d900", 499=>x"9d00"),
---- 15  => (0=>x"9c00", 1=>x"9b00", 2=>x"9d00", 3=>x"9b00", 4=>x"d300", 5=>x"9900", 6=>x"9a00", 7=>x"9a00", 8=>x"9500", 9=>x"c100",
---- 10=>x"9100", 11=>x"9800", 12=>x"9900", 13=>x"9600", 14=>x"9b00", 15=>x"9000", 16=>x"9900", 17=>x"9700", 18=>x"9700",
---- 19=>x"8f00", 20=>x"9b00", 21=>x"9700", 22=>x"9800", 23=>x"9700", 24=>x"9500", 25=>x"9700", 26=>x"9a00", 27=>x"8800",
---- 28=>x"9800", 29=>x"9600", 30=>x"9500", 31=>x"9b00", 32=>x"9500", 33=>x"9a00", 34=>x"9700", 35=>x"9d00", 36=>x"9c00",
---- 37=>x"9c00", 38=>x"9b00", 39=>x"9600", 40=>x"9900", 41=>x"9d00", 42=>x"8f00", 43=>x"8b00", 44=>x"9300", 45=>x"9b00",
---- 46=>x"9700", 47=>x"9600", 48=>x"9300", 49=>x"9100", 50=>x"9600", 51=>x"9400", 52=>x"8f00", 53=>x"9000", 54=>x"8600",
---- 55=>x"9000", 56=>x"9200", 57=>x"9000", 58=>x"8d00", 59=>x"8c00", 60=>x"8d00", 61=>x"9000", 62=>x"8f00", 63=>x"8f00",
---- 64=>x"8e00", 65=>x"8c00", 66=>x"8f00", 67=>x"9200", 68=>x"8d00", 69=>x"8d00", 70=>x"8f00", 71=>x"9200", 72=>x"9200",
---- 73=>x"8d00", 74=>x"8d00", 75=>x"9100", 76=>x"9100", 77=>x"9200", 78=>x"8e00", 79=>x"8f00", 80=>x"9500", 81=>x"8e00",
---- 82=>x"9200", 83=>x"8d00", 84=>x"8f00", 85=>x"9500", 86=>x"9200", 87=>x"9000", 88=>x"8f00", 89=>x"9000", 90=>x"8800",
---- 91=>x"9300", 92=>x"9100", 93=>x"8d00", 94=>x"8f00", 95=>x"7900", 96=>x"9000", 97=>x"9500", 98=>x"8f00", 99=>x"8d00",
---- 100=>x"7600", 101=>x"8500", 102=>x"8b00", 103=>x"8800", 104=>x"8b00", 105=>x"3700", 106=>x"5e00", 107=>x"8500", 108=>x"9a00",
---- 109=>x"8700", 110=>x"e00", 111=>x"7700", 112=>x"dd00", 113=>x"d200", 114=>x"cc00", 115=>x"9200", 116=>x"cf00", 117=>x"b800",
---- 118=>x"d700", 119=>x"e400", 120=>x"c400", 121=>x"c700", 122=>x"cf00", 123=>x"d100", 124=>x"d600", 125=>x"b000", 126=>x"ab00",
---- 127=>x"d500", 128=>x"ca00", 129=>x"ab00", 130=>x"bc00", 131=>x"cb00", 132=>x"c800", 133=>x"cd00", 134=>x"b700", 135=>x"c900",
---- 136=>x"ca00", 137=>x"cc00", 138=>x"ce00", 139=>x"da00", 140=>x"c900", 141=>x"cd00", 142=>x"c900", 143=>x"ca00", 144=>x"d500",
---- 145=>x"ce00", 146=>x"d000", 147=>x"b400", 148=>x"ca00", 149=>x"d600", 150=>x"d300", 151=>x"b500", 152=>x"8e00", 153=>x"af00",
---- 154=>x"c500", 155=>x"cb00", 156=>x"9900", 157=>x"ac00", 158=>x"8600", 159=>x"cc00", 160=>x"a100", 161=>x"a800", 162=>x"9b00",
---- 163=>x"9900", 164=>x"db00", 165=>x"a100", 166=>x"7f00", 167=>x"5f00", 168=>x"a500", 169=>x"b600", 170=>x"5600", 171=>x"4b00",
---- 172=>x"7f00", 173=>x"c500", 174=>x"4400", 175=>x"5200", 176=>x"8a00", 177=>x"d800", 178=>x"9b00", 179=>x"1800", 180=>x"a000",
---- 181=>x"c500", 182=>x"6b00", 183=>x"3f00", 184=>x"2b00", 185=>x"bc00", 186=>x"6700", 187=>x"1c00", 188=>x"2e00", 189=>x"3400",
---- 190=>x"8700", 191=>x"1800", 192=>x"2e00", 193=>x"3400", 194=>x"4f00", 195=>x"1700", 196=>x"2c00", 197=>x"3300", 198=>x"3800",
---- 199=>x"3200", 200=>x"2b00", 201=>x"3600", 202=>x"2f00", 203=>x"3500", 204=>x"5300", 205=>x"3000", 206=>x"3500", 207=>x"5b00",
---- 208=>x"3400", 209=>x"2700", 210=>x"5800", 211=>x"3500", 212=>x"3b00", 213=>x"3400", 214=>x"2a00", 215=>x"3100", 216=>x"3800",
---- 217=>x"3d00", 218=>x"2900", 219=>x"2b00", 220=>x"4900", 221=>x"4900", 222=>x"4d00", 223=>x"5b00", 224=>x"3000", 225=>x"3900",
---- 226=>x"3c00", 227=>x"3600", 228=>x"2900", 229=>x"3600", 230=>x"3d00", 231=>x"3f00", 232=>x"2e00", 233=>x"3400", 234=>x"2e00",
---- 235=>x"4100", 236=>x"3b00", 237=>x"3000", 238=>x"3600", 239=>x"2600", 240=>x"4100", 241=>x"3300", 242=>x"2d00", 243=>x"3300",
---- 244=>x"4200", 245=>x"3f00", 246=>x"2d00", 247=>x"5300", 248=>x"3100", 249=>x"3b00", 250=>x"3600", 251=>x"2d00", 252=>x"4600",
---- 253=>x"3100", 254=>x"5700", 255=>x"3300", 256=>x"2f00", 257=>x"3200", 258=>x"2800", 259=>x"7600", 260=>x"4d00", 261=>x"3200",
---- 262=>x"2a00", 263=>x"5700", 264=>x"8e00", 265=>x"2b00", 266=>x"3200", 267=>x"2c00", 268=>x"4c00", 269=>x"9100", 270=>x"2d00",
---- 271=>x"3400", 272=>x"2e00", 273=>x"7a00", 274=>x"8700", 275=>x"2b00", 276=>x"5600", 277=>x"2700", 278=>x"8900", 279=>x"8500",
---- 280=>x"2d00", 281=>x"2b00", 282=>x"6400", 283=>x"8a00", 284=>x"8d00", 285=>x"3000", 286=>x"2500", 287=>x"6900", 288=>x"8b00",
---- 289=>x"9800", 290=>x"3c00", 291=>x"2500", 292=>x"8100", 293=>x"8c00", 294=>x"a400", 295=>x"3500", 296=>x"5200", 297=>x"8c00",
---- 298=>x"8f00", 299=>x"a000", 300=>x"2a00", 301=>x"5300", 302=>x"8e00", 303=>x"9900", 304=>x"9b00", 305=>x"2100", 306=>x"7700",
---- 307=>x"8e00", 308=>x"9e00", 309=>x"9c00", 310=>x"2000", 311=>x"8e00", 312=>x"9100", 313=>x"9f00", 314=>x"9b00", 315=>x"3f00",
---- 316=>x"9800", 317=>x"9400", 318=>x"9f00", 319=>x"9900", 320=>x"5b00", 321=>x"9700", 322=>x"9800", 323=>x"9c00", 324=>x"9b00",
---- 325=>x"7b00", 326=>x"9300", 327=>x"9d00", 328=>x"9900", 329=>x"7b00", 330=>x"8d00", 331=>x"9200", 332=>x"9c00", 333=>x"9a00",
---- 334=>x"9a00", 335=>x"9000", 336=>x"9200", 337=>x"9c00", 338=>x"9900", 339=>x"9600", 340=>x"9400", 341=>x"9400", 342=>x"9d00",
---- 343=>x"9700", 344=>x"9700", 345=>x"9400", 346=>x"9800", 347=>x"9b00", 348=>x"9700", 349=>x"9800", 350=>x"9700", 351=>x"9800",
---- 352=>x"9d00", 353=>x"9a00", 354=>x"9900", 355=>x"9500", 356=>x"9a00", 357=>x"8f00", 358=>x"9700", 359=>x"9a00", 360=>x"9300",
---- 361=>x"9c00", 362=>x"9e00", 363=>x"9100", 364=>x"9a00", 365=>x"9100", 366=>x"9f00", 367=>x"9b00", 368=>x"9800", 369=>x"9600",
---- 370=>x"9300", 371=>x"9900", 372=>x"9a00", 373=>x"9500", 374=>x"9800", 375=>x"7800", 376=>x"7800", 377=>x"8400", 378=>x"8c00",
---- 379=>x"8900", 380=>x"6c00", 381=>x"6b00", 382=>x"7000", 383=>x"7300", 384=>x"7600", 385=>x"8000", 386=>x"8400", 387=>x"7900",
---- 388=>x"7200", 389=>x"6b00", 390=>x"8e00", 391=>x"8d00", 392=>x"8700", 393=>x"8200", 394=>x"8100", 395=>x"9600", 396=>x"9100",
---- 397=>x"8e00", 398=>x"8c00", 399=>x"8900", 400=>x"8d00", 401=>x"9100", 402=>x"8600", 403=>x"8f00", 404=>x"8c00", 405=>x"9500",
---- 406=>x"9100", 407=>x"8b00", 408=>x"8f00", 409=>x"8d00", 410=>x"9100", 411=>x"9000", 412=>x"9000", 413=>x"8c00", 414=>x"8d00",
---- 415=>x"9600", 416=>x"9000", 417=>x"8f00", 418=>x"8e00", 419=>x"8a00", 420=>x"8900", 421=>x"9300", 422=>x"9000", 423=>x"8b00",
---- 424=>x"8700", 425=>x"9100", 426=>x"8800", 427=>x"8d00", 428=>x"8b00", 429=>x"8900", 430=>x"8800", 431=>x"8e00", 432=>x"8a00",
---- 433=>x"8b00", 434=>x"8b00", 435=>x"8f00", 436=>x"8e00", 437=>x"8900", 438=>x"8a00", 439=>x"8b00", 440=>x"9100", 441=>x"9100",
---- 442=>x"8f00", 443=>x"8d00", 444=>x"8c00", 445=>x"7f00", 446=>x"8b00", 447=>x"9200", 448=>x"9200", 449=>x"9000", 450=>x"5300",
---- 451=>x"6300", 452=>x"7300", 453=>x"7d00", 454=>x"8600", 455=>x"6500", 456=>x"4600", 457=>x"4400", 458=>x"4400", 459=>x"4c00",
---- 460=>x"6200", 461=>x"5a00", 462=>x"4900", 463=>x"5400", 464=>x"2a00", 465=>x"7e00", 466=>x"6600", 467=>x"5e00", 468=>x"4e00",
---- 469=>x"3e00", 470=>x"6b00", 471=>x"6900", 472=>x"6000", 473=>x"5d00", 474=>x"4e00", 475=>x"6300", 476=>x"6700", 477=>x"6300",
---- 478=>x"6f00", 479=>x"5900", 480=>x"5a00", 481=>x"6400", 482=>x"6d00", 483=>x"6800", 484=>x"6700", 485=>x"5300", 486=>x"6300",
---- 487=>x"7100", 488=>x"7000", 489=>x"7600", 490=>x"4700", 491=>x"6100", 492=>x"6700", 493=>x"7200", 494=>x"7800", 495=>x"4f00",
---- 496=>x"5a00", 497=>x"5e00", 498=>x"6c00", 499=>x"7800"),
---- 16  => (0=>x"b300", 1=>x"e100", 2=>x"a000", 3=>x"6300", 4=>x"7000", 5=>x"dc00", 6=>x"e100", 7=>x"9400", 8=>x"6800", 9=>x"7200",
---- 10=>x"d100", 11=>x"db00", 12=>x"e000", 13=>x"9a00", 14=>x"6000", 15=>x"b600", 16=>x"da00", 17=>x"de00", 18=>x"d200",
---- 19=>x"6a00", 20=>x"8b00", 21=>x"cd00", 22=>x"dc00", 23=>x"e400", 24=>x"a800", 25=>x"8e00", 26=>x"ae00", 27=>x"ca00",
---- 28=>x"ce00", 29=>x"e000", 30=>x"9300", 31=>x"8b00", 32=>x"ac00", 33=>x"b600", 34=>x"be00", 35=>x"9300", 36=>x"8900",
---- 37=>x"a200", 38=>x"dd00", 39=>x"e300", 40=>x"8f00", 41=>x"8b00", 42=>x"8800", 43=>x"c400", 44=>x"e100", 45=>x"8f00",
---- 46=>x"8e00", 47=>x"8b00", 48=>x"9900", 49=>x"d800", 50=>x"8600", 51=>x"8c00", 52=>x"8c00", 53=>x"8600", 54=>x"bb00",
---- 55=>x"8b00", 56=>x"8b00", 57=>x"8d00", 58=>x"8a00", 59=>x"8700", 60=>x"8c00", 61=>x"8c00", 62=>x"9000", 63=>x"9000",
---- 64=>x"8600", 65=>x"8c00", 66=>x"8f00", 67=>x"8e00", 68=>x"8600", 69=>x"9100", 70=>x"8f00", 71=>x"9100", 72=>x"8a00",
---- 73=>x"9300", 74=>x"8f00", 75=>x"9000", 76=>x"9000", 77=>x"8a00", 78=>x"9500", 79=>x"9b00", 80=>x"9100", 81=>x"9100",
---- 82=>x"9200", 83=>x"9500", 84=>x"a300", 85=>x"8d00", 86=>x"8a00", 87=>x"9200", 88=>x"a100", 89=>x"6b00", 90=>x"9100",
---- 91=>x"9200", 92=>x"9500", 93=>x"9300", 94=>x"2100", 95=>x"8a00", 96=>x"8b00", 97=>x"9f00", 98=>x"4300", 99=>x"2100",
---- 100=>x"8700", 101=>x"9c00", 102=>x"7000", 103=>x"1f00", 104=>x"2800", 105=>x"9200", 106=>x"8f00", 107=>x"2700", 108=>x"2600",
---- 109=>x"5300", 110=>x"db00", 111=>x"6500", 112=>x"2100", 113=>x"2f00", 114=>x"2f00", 115=>x"f300", 116=>x"9200", 117=>x"1d00",
---- 118=>x"2b00", 119=>x"3700", 120=>x"df00", 121=>x"ce00", 122=>x"1400", 123=>x"5300", 124=>x"3100", 125=>x"e300", 126=>x"d700",
---- 127=>x"1400", 128=>x"2e00", 129=>x"3700", 130=>x"dd00", 131=>x"be00", 132=>x"1700", 133=>x"3000", 134=>x"3400", 135=>x"e900",
---- 136=>x"8d00", 137=>x"4800", 138=>x"3100", 139=>x"3100", 140=>x"ee00", 141=>x"6900", 142=>x"2400", 143=>x"3200", 144=>x"3600",
---- 145=>x"e800", 146=>x"3600", 147=>x"2700", 148=>x"2f00", 149=>x"3400", 150=>x"bd00", 151=>x"1a00", 152=>x"2f00", 153=>x"3000",
---- 154=>x"2a00", 155=>x"6b00", 156=>x"1d00", 157=>x"3500", 158=>x"5300", 159=>x"2800", 160=>x"2400", 161=>x"2c00", 162=>x"3000",
---- 163=>x"3100", 164=>x"3300", 165=>x"3900", 166=>x"2d00", 167=>x"3200", 168=>x"3000", 169=>x"3c00", 170=>x"3700", 171=>x"2e00",
---- 172=>x"2c00", 173=>x"3200", 174=>x"3100", 175=>x"3f00", 176=>x"3100", 177=>x"2d00", 178=>x"3500", 179=>x"2200", 180=>x"3100",
---- 181=>x"2d00", 182=>x"3400", 183=>x"3500", 184=>x"2e00", 185=>x"3100", 186=>x"2900", 187=>x"3900", 188=>x"3300", 189=>x"5b00",
---- 190=>x"3300", 191=>x"2f00", 192=>x"3300", 193=>x"2700", 194=>x"8a00", 195=>x"2d00", 196=>x"3c00", 197=>x"2d00", 198=>x"4900",
---- 199=>x"9200", 200=>x"2700", 201=>x"4800", 202=>x"3100", 203=>x"6e00", 204=>x"8200", 205=>x"3000", 206=>x"2c00", 207=>x"4200",
---- 208=>x"8500", 209=>x"7800", 210=>x"3b00", 211=>x"3e00", 212=>x"7d00", 213=>x"8700", 214=>x"8100", 215=>x"2f00", 216=>x"3100",
---- 217=>x"8700", 218=>x"8300", 219=>x"8a00", 220=>x"2b00", 221=>x"4800", 222=>x"9300", 223=>x"8700", 224=>x"a600", 225=>x"2500",
---- 226=>x"7a00", 227=>x"8c00", 228=>x"8d00", 229=>x"a800", 230=>x"3d00", 231=>x"9000", 232=>x"8100", 233=>x"a300", 234=>x"a200",
---- 235=>x"6100", 236=>x"8d00", 237=>x"8a00", 238=>x"a300", 239=>x"a300", 240=>x"8400", 241=>x"8200", 242=>x"9800", 243=>x"a400",
---- 244=>x"8f00", 245=>x"8d00", 246=>x"8100", 247=>x"a100", 248=>x"a000", 249=>x"9f00", 250=>x"8d00", 251=>x"8b00", 252=>x"a200",
---- 253=>x"9e00", 254=>x"9900", 255=>x"8c00", 256=>x"9b00", 257=>x"9f00", 258=>x"9d00", 259=>x"8100", 260=>x"8a00", 261=>x"9e00",
---- 262=>x"9d00", 263=>x"9e00", 264=>x"8900", 265=>x"9100", 266=>x"9f00", 267=>x"9b00", 268=>x"9900", 269=>x"8e00", 270=>x"9a00",
---- 271=>x"9d00", 272=>x"9a00", 273=>x"9800", 274=>x"9700", 275=>x"9e00", 276=>x"9b00", 277=>x"9800", 278=>x"9600", 279=>x"8c00",
---- 280=>x"a000", 281=>x"8e00", 282=>x"9800", 283=>x"9800", 284=>x"9700", 285=>x"9d00", 286=>x"9a00", 287=>x"9800", 288=>x"9800",
---- 289=>x"9600", 290=>x"9b00", 291=>x"9900", 292=>x"9900", 293=>x"8c00", 294=>x"9000", 295=>x"9a00", 296=>x"9a00", 297=>x"9800",
---- 298=>x"9500", 299=>x"9300", 300=>x"9900", 301=>x"9900", 302=>x"9900", 303=>x"9700", 304=>x"9400", 305=>x"9800", 306=>x"9700",
---- 307=>x"9800", 308=>x"9700", 309=>x"9500", 310=>x"9900", 311=>x"9700", 312=>x"8100", 313=>x"9600", 314=>x"9500", 315=>x"9500",
---- 316=>x"9500", 317=>x"9800", 318=>x"9400", 319=>x"9300", 320=>x"9700", 321=>x"9600", 322=>x"8b00", 323=>x"9600", 324=>x"9200",
---- 325=>x"9700", 326=>x"9400", 327=>x"9500", 328=>x"9100", 329=>x"9300", 330=>x"9500", 331=>x"9400", 332=>x"9400", 333=>x"9000",
---- 334=>x"8c00", 335=>x"9000", 336=>x"8e00", 337=>x"9400", 338=>x"9200", 339=>x"9200", 340=>x"9500", 341=>x"9400", 342=>x"9300",
---- 343=>x"9400", 344=>x"8800", 345=>x"9500", 346=>x"8f00", 347=>x"8900", 348=>x"9300", 349=>x"9300", 350=>x"9700", 351=>x"9700",
---- 352=>x"9600", 353=>x"9200", 354=>x"8c00", 355=>x"9a00", 356=>x"9a00", 357=>x"9500", 358=>x"9300", 359=>x"8e00", 360=>x"9800",
---- 361=>x"9900", 362=>x"9400", 363=>x"9400", 364=>x"9000", 365=>x"9500", 366=>x"9500", 367=>x"9800", 368=>x"8b00", 369=>x"8e00",
---- 370=>x"9400", 371=>x"9200", 372=>x"9400", 373=>x"9000", 374=>x"8b00", 375=>x"9400", 376=>x"9600", 377=>x"9200", 378=>x"8e00",
---- 379=>x"8700", 380=>x"7c00", 381=>x"8500", 382=>x"8400", 383=>x"8b00", 384=>x"8a00", 385=>x"6600", 386=>x"6500", 387=>x"6c00",
---- 388=>x"6f00", 389=>x"8200", 390=>x"7c00", 391=>x"6a00", 392=>x"6100", 393=>x"5c00", 394=>x"5d00", 395=>x"8300", 396=>x"7d00",
---- 397=>x"7400", 398=>x"6b00", 399=>x"6900", 400=>x"8900", 401=>x"8400", 402=>x"8100", 403=>x"7b00", 404=>x"7500", 405=>x"8c00",
---- 406=>x"8600", 407=>x"8400", 408=>x"7e00", 409=>x"7d00", 410=>x"8400", 411=>x"8900", 412=>x"8400", 413=>x"7f00", 414=>x"7800",
---- 415=>x"8700", 416=>x"8600", 417=>x"8100", 418=>x"7900", 419=>x"8300", 420=>x"8500", 421=>x"8200", 422=>x"7f00", 423=>x"7500",
---- 424=>x"a400", 425=>x"8400", 426=>x"8100", 427=>x"7b00", 428=>x"6f00", 429=>x"d800", 430=>x"8700", 431=>x"7f00", 432=>x"7900",
---- 433=>x"8600", 434=>x"d900", 435=>x"8700", 436=>x"7f00", 437=>x"7d00", 438=>x"8a00", 439=>x"d900", 440=>x"8700", 441=>x"8000",
---- 442=>x"8500", 443=>x"8400", 444=>x"af00", 445=>x"8c00", 446=>x"8100", 447=>x"9100", 448=>x"9000", 449=>x"8100", 450=>x"8d00",
---- 451=>x"9300", 452=>x"9f00", 453=>x"8800", 454=>x"7f00", 455=>x"5800", 456=>x"7e00", 457=>x"9300", 458=>x"9e00", 459=>x"9300",
---- 460=>x"2300", 461=>x"3100", 462=>x"9d00", 463=>x"cc00", 464=>x"9000", 465=>x"2700", 466=>x"1f00", 467=>x"c000", 468=>x"c500",
---- 469=>x"ae00", 470=>x"4100", 471=>x"3c00", 472=>x"a800", 473=>x"d500", 474=>x"c400", 475=>x"5f00", 476=>x"5400", 477=>x"a800",
---- 478=>x"d600", 479=>x"8c00", 480=>x"7300", 481=>x"6b00", 482=>x"7600", 483=>x"7600", 484=>x"4c00", 485=>x"7500", 486=>x"7200",
---- 487=>x"7100", 488=>x"5f00", 489=>x"6500", 490=>x"7a00", 491=>x"7300", 492=>x"6e00", 493=>x"6d00", 494=>x"7900", 495=>x"8200",
---- 496=>x"7900", 497=>x"7b00", 498=>x"8600", 499=>x"8100"),
---- 17  => (0=>x"7800", 1=>x"7900", 2=>x"7a00", 3=>x"7a00", 4=>x"7800", 5=>x"7800", 6=>x"7a00", 7=>x"7a00", 8=>x"7a00", 9=>x"7800",
---- 10=>x"6f00", 11=>x"7b00", 12=>x"7700", 13=>x"7900", 14=>x"7700", 15=>x"7200", 16=>x"7300", 17=>x"7600", 18=>x"7c00",
---- 19=>x"7a00", 20=>x"6000", 21=>x"7000", 22=>x"7600", 23=>x"7600", 24=>x"7900", 25=>x"7a00", 26=>x"6900", 27=>x"7600",
---- 28=>x"7a00", 29=>x"7c00", 30=>x"c900", 31=>x"6300", 32=>x"7000", 33=>x"7600", 34=>x"7900", 35=>x"e700", 36=>x"9300",
---- 37=>x"5f00", 38=>x"7100", 39=>x"7700", 40=>x"b700", 41=>x"d900", 42=>x"6400", 43=>x"6900", 44=>x"6f00", 45=>x"e900",
---- 46=>x"bc00", 47=>x"aa00", 48=>x"6300", 49=>x"7b00", 50=>x"b700", 51=>x"cb00", 52=>x"d400", 53=>x"8400", 54=>x"6800",
---- 55=>x"d600", 56=>x"e300", 57=>x"eb00", 58=>x"cc00", 59=>x"2100", 60=>x"a500", 61=>x"e100", 62=>x"f600", 63=>x"8f00",
---- 64=>x"1900", 65=>x"8d00", 66=>x"da00", 67=>x"aa00", 68=>x"1d00", 69=>x"2600", 70=>x"9c00", 71=>x"8200", 72=>x"2000",
---- 73=>x"2600", 74=>x"5200", 75=>x"9a00", 76=>x"2e00", 77=>x"2600", 78=>x"2b00", 79=>x"2d00", 80=>x"4400", 81=>x"1e00",
---- 82=>x"3d00", 83=>x"2f00", 84=>x"3600", 85=>x"2900", 86=>x"2900", 87=>x"3f00", 88=>x"3600", 89=>x"3700", 90=>x"2900",
---- 91=>x"4d00", 92=>x"5300", 93=>x"3100", 94=>x"2d00", 95=>x"2900", 96=>x"3600", 97=>x"3500", 98=>x"3700", 99=>x"2d00",
---- 100=>x"3100", 101=>x"3700", 102=>x"3400", 103=>x"4800", 104=>x"4900", 105=>x"3100", 106=>x"3400", 107=>x"3100", 108=>x"2b00",
---- 109=>x"5400", 110=>x"5200", 111=>x"3200", 112=>x"5600", 113=>x"3200", 114=>x"2b00", 115=>x"3800", 116=>x"3300", 117=>x"3300",
---- 118=>x"3b00", 119=>x"3300", 120=>x"3500", 121=>x"2f00", 122=>x"2e00", 123=>x"3c00", 124=>x"3700", 125=>x"2c00", 126=>x"2900",
---- 127=>x"5300", 128=>x"3000", 129=>x"2a00", 130=>x"3400", 131=>x"2c00", 132=>x"3000", 133=>x"3300", 134=>x"1600", 135=>x"2f00",
---- 136=>x"2900", 137=>x"2f00", 138=>x"4a00", 139=>x"6900", 140=>x"2b00", 141=>x"2f00", 142=>x"3300", 143=>x"3b00", 144=>x"7c00",
---- 145=>x"2500", 146=>x"3600", 147=>x"2900", 148=>x"5c00", 149=>x"9400", 150=>x"7700", 151=>x"2800", 152=>x"3700", 153=>x"8a00",
---- 154=>x"9600", 155=>x"2800", 156=>x"3400", 157=>x"6e00", 158=>x"9b00", 159=>x"9100", 160=>x"2e00", 161=>x"4700", 162=>x"9700",
---- 163=>x"9400", 164=>x"8900", 165=>x"3000", 166=>x"6d00", 167=>x"9d00", 168=>x"9000", 169=>x"9e00", 170=>x"3d00", 171=>x"9600",
---- 172=>x"9300", 173=>x"9900", 174=>x"a200", 175=>x"6600", 176=>x"9a00", 177=>x"8800", 178=>x"a300", 179=>x"a000", 180=>x"8700",
---- 181=>x"8a00", 182=>x"9d00", 183=>x"a400", 184=>x"a300", 185=>x"9c00", 186=>x"9100", 187=>x"a500", 188=>x"a500", 189=>x"9000",
---- 190=>x"9300", 191=>x"9800", 192=>x"a600", 193=>x"a600", 194=>x"a600", 195=>x"8900", 196=>x"a500", 197=>x"a700", 198=>x"9300",
---- 199=>x"a400", 200=>x"8e00", 201=>x"aa00", 202=>x"a500", 203=>x"a300", 204=>x"a200", 205=>x"9d00", 206=>x"a800", 207=>x"a600",
---- 208=>x"a300", 209=>x"a200", 210=>x"a000", 211=>x"a600", 212=>x"a500", 213=>x"a500", 214=>x"a100", 215=>x"9200", 216=>x"9900",
---- 217=>x"a100", 218=>x"a400", 219=>x"a300", 220=>x"9900", 221=>x"9700", 222=>x"8900", 223=>x"9500", 224=>x"9800", 225=>x"a200",
---- 226=>x"9c00", 227=>x"9800", 228=>x"9600", 229=>x"9500", 230=>x"a200", 231=>x"9f00", 232=>x"a400", 233=>x"9d00", 234=>x"9e00",
---- 235=>x"a000", 236=>x"a000", 237=>x"a500", 238=>x"9b00", 239=>x"a500", 240=>x"9f00", 241=>x"9a00", 242=>x"9c00", 243=>x"a000",
---- 244=>x"a100", 245=>x"9e00", 246=>x"8b00", 247=>x"9900", 248=>x"9c00", 249=>x"9a00", 250=>x"9800", 251=>x"9d00", 252=>x"9b00",
---- 253=>x"9b00", 254=>x"9e00", 255=>x"9900", 256=>x"9900", 257=>x"9b00", 258=>x"9b00", 259=>x"8f00", 260=>x"9500", 261=>x"9700",
---- 262=>x"9900", 263=>x"9900", 264=>x"8d00", 265=>x"9a00", 266=>x"9e00", 267=>x"9700", 268=>x"9a00", 269=>x"9800", 270=>x"9600",
---- 271=>x"9a00", 272=>x"9600", 273=>x"9700", 274=>x"9900", 275=>x"9700", 276=>x"9600", 277=>x"9600", 278=>x"9700", 279=>x"8a00",
---- 280=>x"9900", 281=>x"8b00", 282=>x"9600", 283=>x"9300", 284=>x"9100", 285=>x"9700", 286=>x"9400", 287=>x"9200", 288=>x"8800",
---- 289=>x"8900", 290=>x"8f00", 291=>x"9400", 292=>x"9200", 293=>x"9200", 294=>x"8600", 295=>x"9300", 296=>x"8900", 297=>x"8a00",
---- 298=>x"8800", 299=>x"8a00", 300=>x"9300", 301=>x"9100", 302=>x"8e00", 303=>x"8b00", 304=>x"8400", 305=>x"9500", 306=>x"9300",
---- 307=>x"8e00", 308=>x"8600", 309=>x"8000", 310=>x"8a00", 311=>x"8b00", 312=>x"9000", 313=>x"8500", 314=>x"8500", 315=>x"8a00",
---- 316=>x"9200", 317=>x"8600", 318=>x"8000", 319=>x"a100", 320=>x"9000", 321=>x"8f00", 322=>x"8d00", 323=>x"7f00", 324=>x"b100",
---- 325=>x"9200", 326=>x"8e00", 327=>x"8500", 328=>x"8300", 329=>x"b900", 330=>x"8e00", 331=>x"8e00", 332=>x"8400", 333=>x"8900",
---- 334=>x"c100", 335=>x"9000", 336=>x"8c00", 337=>x"8400", 338=>x"8b00", 339=>x"c100", 340=>x"9100", 341=>x"8e00", 342=>x"7d00",
---- 343=>x"8200", 344=>x"c300", 345=>x"8900", 346=>x"8e00", 347=>x"7e00", 348=>x"9a00", 349=>x"d100", 350=>x"9000", 351=>x"8c00",
---- 352=>x"7c00", 353=>x"8f00", 354=>x"d900", 355=>x"8e00", 356=>x"8800", 357=>x"7500", 358=>x"9900", 359=>x"dc00", 360=>x"8d00",
---- 361=>x"8300", 362=>x"7300", 363=>x"9700", 364=>x"e200", 365=>x"8b00", 366=>x"8600", 367=>x"7300", 368=>x"9100", 369=>x"b200",
---- 370=>x"8a00", 371=>x"8200", 372=>x"6f00", 373=>x"c000", 374=>x"e600", 375=>x"8600", 376=>x"7f00", 377=>x"7600", 378=>x"ab00",
---- 379=>x"e000", 380=>x"8600", 381=>x"7600", 382=>x"8900", 383=>x"df00", 384=>x"d700", 385=>x"7300", 386=>x"7500", 387=>x"8200",
---- 388=>x"ca00", 389=>x"ce00", 390=>x"7000", 391=>x"5800", 392=>x"6800", 393=>x"cf00", 394=>x"cc00", 395=>x"8700", 396=>x"5d00",
---- 397=>x"7c00", 398=>x"d800", 399=>x"d200", 400=>x"8300", 401=>x"6800", 402=>x"ae00", 403=>x"d700", 404=>x"d500", 405=>x"8900",
---- 406=>x"7b00", 407=>x"a500", 408=>x"da00", 409=>x"d500", 410=>x"8a00", 411=>x"9d00", 412=>x"d200", 413=>x"d700", 414=>x"d500",
---- 415=>x"b500", 416=>x"cc00", 417=>x"ad00", 418=>x"dc00", 419=>x"d700", 420=>x"ca00", 421=>x"cd00", 422=>x"db00", 423=>x"d800",
---- 424=>x"d300", 425=>x"dc00", 426=>x"d300", 427=>x"d900", 428=>x"da00", 429=>x"c100", 430=>x"d300", 431=>x"c200", 432=>x"8d00",
---- 433=>x"dd00", 434=>x"9900", 435=>x"d100", 436=>x"cd00", 437=>x"b800", 438=>x"ca00", 439=>x"7a00", 440=>x"bd00", 441=>x"d400",
---- 442=>x"dd00", 443=>x"b600", 444=>x"6f00", 445=>x"9e00", 446=>x"df00", 447=>x"da00", 448=>x"a100", 449=>x"6d00", 450=>x"9600",
---- 451=>x"cc00", 452=>x"c700", 453=>x"8800", 454=>x"6100", 455=>x"ce00", 456=>x"b700", 457=>x"a700", 458=>x"6300", 459=>x"4000",
---- 460=>x"cc00", 461=>x"cd00", 462=>x"8f00", 463=>x"5000", 464=>x"3c00", 465=>x"db00", 466=>x"ad00", 467=>x"3500", 468=>x"5400",
---- 469=>x"4600", 470=>x"9c00", 471=>x"4400", 472=>x"2f00", 473=>x"3e00", 474=>x"5c00", 475=>x"4a00", 476=>x"3800", 477=>x"4600",
---- 478=>x"5f00", 479=>x"5400", 480=>x"4f00", 481=>x"6300", 482=>x"4f00", 483=>x"4d00", 484=>x"6d00", 485=>x"7800", 486=>x"5600",
---- 487=>x"4f00", 488=>x"6200", 489=>x"5600", 490=>x"7900", 491=>x"5e00", 492=>x"6500", 493=>x"5c00", 494=>x"4c00", 495=>x"6200",
---- 496=>x"6c00", 497=>x"5000", 498=>x"4f00", 499=>x"5a00"),
---- 18  => (0=>x"7900", 1=>x"7b00", 2=>x"7d00", 3=>x"7900", 4=>x"7e00", 5=>x"7c00", 6=>x"7d00", 7=>x"7a00", 8=>x"7a00", 9=>x"7c00",
---- 10=>x"7900", 11=>x"7800", 12=>x"7b00", 13=>x"7b00", 14=>x"7c00", 15=>x"7900", 16=>x"7b00", 17=>x"7c00", 18=>x"7e00",
---- 19=>x"8100", 20=>x"7700", 21=>x"7a00", 22=>x"8100", 23=>x"8200", 24=>x"8e00", 25=>x"7b00", 26=>x"7a00", 27=>x"7c00",
---- 28=>x"8c00", 29=>x"6f00", 30=>x"7900", 31=>x"7d00", 32=>x"8a00", 33=>x"6d00", 34=>x"4400", 35=>x"7c00", 36=>x"8700",
---- 37=>x"6b00", 38=>x"2200", 39=>x"3800", 40=>x"8200", 41=>x"6e00", 42=>x"2700", 43=>x"2600", 44=>x"4000", 45=>x"6600",
---- 46=>x"2300", 47=>x"3f00", 48=>x"4000", 49=>x"3c00", 50=>x"4d00", 51=>x"2400", 52=>x"3b00", 53=>x"2e00", 54=>x"3400",
---- 55=>x"2400", 56=>x"2c00", 57=>x"3200", 58=>x"3500", 59=>x"3500", 60=>x"2b00", 61=>x"3000", 62=>x"3300", 63=>x"3600",
---- 64=>x"2e00", 65=>x"2b00", 66=>x"2b00", 67=>x"5200", 68=>x"2f00", 69=>x"2d00", 70=>x"2c00", 71=>x"7a00", 72=>x"2b00",
---- 73=>x"5100", 74=>x"3600", 75=>x"3500", 76=>x"2b00", 77=>x"2a00", 78=>x"3400", 79=>x"2f00", 80=>x"3400", 81=>x"2a00",
---- 82=>x"3300", 83=>x"2f00", 84=>x"5200", 85=>x"2e00", 86=>x"3200", 87=>x"3500", 88=>x"2a00", 89=>x"3600", 90=>x"2c00",
---- 91=>x"3a00", 92=>x"2e00", 93=>x"3400", 94=>x"3800", 95=>x"3600", 96=>x"2900", 97=>x"3400", 98=>x"3500", 99=>x"3800",
---- 100=>x"4f00", 101=>x"5500", 102=>x"3000", 103=>x"4000", 104=>x"6600", 105=>x"2a00", 106=>x"3300", 107=>x"2100", 108=>x"4a00",
---- 109=>x"9600", 110=>x"3700", 111=>x"4800", 112=>x"4a00", 113=>x"8c00", 114=>x"9400", 115=>x"3500", 116=>x"2900", 117=>x"7700",
---- 118=>x"9c00", 119=>x"8b00", 120=>x"2c00", 121=>x"5300", 122=>x"9f00", 123=>x"8700", 124=>x"9600", 125=>x"2a00", 126=>x"9700",
---- 127=>x"9600", 128=>x"9400", 129=>x"a300", 130=>x"6700", 131=>x"a100", 132=>x"8f00", 133=>x"a000", 134=>x"a100", 135=>x"8a00",
---- 136=>x"9400", 137=>x"9800", 138=>x"a200", 139=>x"9f00", 140=>x"9a00", 141=>x"9100", 142=>x"a000", 143=>x"9f00", 144=>x"9e00",
---- 145=>x"9000", 146=>x"9c00", 147=>x"a100", 148=>x"a000", 149=>x"9f00", 150=>x"9600", 151=>x"a100", 152=>x"a200", 153=>x"9f00",
---- 154=>x"a000", 155=>x"9e00", 156=>x"a100", 157=>x"a100", 158=>x"9f00", 159=>x"9f00", 160=>x"a100", 161=>x"a000", 162=>x"8f00",
---- 163=>x"9200", 164=>x"9000", 165=>x"a000", 166=>x"9d00", 167=>x"9d00", 168=>x"9c00", 169=>x"9e00", 170=>x"9f00", 171=>x"9e00",
---- 172=>x"9b00", 173=>x"9d00", 174=>x"9c00", 175=>x"9f00", 176=>x"a000", 177=>x"9e00", 178=>x"9c00", 179=>x"8d00", 180=>x"a000",
---- 181=>x"9f00", 182=>x"9e00", 183=>x"9200", 184=>x"9d00", 185=>x"a300", 186=>x"a000", 187=>x"a000", 188=>x"a000", 189=>x"9c00",
---- 190=>x"a200", 191=>x"a400", 192=>x"9000", 193=>x"9400", 194=>x"9d00", 195=>x"a400", 196=>x"9200", 197=>x"a400", 198=>x"9c00",
---- 199=>x"9d00", 200=>x"a400", 201=>x"9b00", 202=>x"9900", 203=>x"a000", 204=>x"9f00", 205=>x"a400", 206=>x"a200", 207=>x"a300",
---- 208=>x"a200", 209=>x"9100", 210=>x"a200", 211=>x"a200", 212=>x"a200", 213=>x"a100", 214=>x"a100", 215=>x"a100", 216=>x"a100",
---- 217=>x"a400", 218=>x"a100", 219=>x"9e00", 220=>x"9d00", 221=>x"9700", 222=>x"9b00", 223=>x"a300", 224=>x"a200", 225=>x"9200",
---- 226=>x"9200", 227=>x"8900", 228=>x"9d00", 229=>x"8600", 230=>x"9b00", 231=>x"9000", 232=>x"9300", 233=>x"8f00", 234=>x"8e00",
---- 235=>x"9d00", 236=>x"9a00", 237=>x"9500", 238=>x"9000", 239=>x"9000", 240=>x"9c00", 241=>x"9b00", 242=>x"9b00", 243=>x"9900",
---- 244=>x"9800", 245=>x"9300", 246=>x"9a00", 247=>x"9a00", 248=>x"9b00", 249=>x"9e00", 250=>x"9b00", 251=>x"9700", 252=>x"9a00",
---- 253=>x"9a00", 254=>x"8e00", 255=>x"9a00", 256=>x"9a00", 257=>x"8e00", 258=>x"9000", 259=>x"9600", 260=>x"9900", 261=>x"9600",
---- 262=>x"9500", 263=>x"9300", 264=>x"9100", 265=>x"9600", 266=>x"9400", 267=>x"9300", 268=>x"8e00", 269=>x"8c00", 270=>x"9300",
---- 271=>x"9000", 272=>x"8a00", 273=>x"8700", 274=>x"8200", 275=>x"9100", 276=>x"8e00", 277=>x"8800", 278=>x"8000", 279=>x"9e00",
---- 280=>x"8d00", 281=>x"8a00", 282=>x"7e00", 283=>x"a400", 284=>x"c300", 285=>x"8900", 286=>x"8000", 287=>x"9b00", 288=>x"ad00",
---- 289=>x"c700", 290=>x"8400", 291=>x"8600", 292=>x"bc00", 293=>x"c800", 294=>x"c000", 295=>x"7d00", 296=>x"ad00", 297=>x"c800",
---- 298=>x"c100", 299=>x"c000", 300=>x"8500", 301=>x"c600", 302=>x"a500", 303=>x"c200", 304=>x"c300", 305=>x"b200", 306=>x"c800",
---- 307=>x"c400", 308=>x"c100", 309=>x"cc00", 310=>x"b500", 311=>x"be00", 312=>x"c100", 313=>x"c500", 314=>x"ce00", 315=>x"c800",
---- 316=>x"ae00", 317=>x"c600", 318=>x"ce00", 319=>x"d100", 320=>x"c700", 321=>x"bb00", 322=>x"cc00", 323=>x"d300", 324=>x"ac00",
---- 325=>x"c600", 326=>x"b600", 327=>x"d400", 328=>x"cf00", 329=>x"d200", 330=>x"c600", 331=>x"bd00", 332=>x"c100", 333=>x"d000",
---- 334=>x"d100", 335=>x"ca00", 336=>x"d300", 337=>x"d200", 338=>x"d000", 339=>x"d400", 340=>x"d500", 341=>x"d300", 342=>x"d100",
---- 343=>x"d400", 344=>x"cf00", 345=>x"aa00", 346=>x"d600", 347=>x"d100", 348=>x"b100", 349=>x"b000", 350=>x"bd00", 351=>x"d800",
---- 352=>x"d300", 353=>x"da00", 354=>x"d400", 355=>x"de00", 356=>x"af00", 357=>x"d800", 358=>x"da00", 359=>x"d300", 360=>x"da00",
---- 361=>x"d900", 362=>x"d700", 363=>x"d800", 364=>x"d300", 365=>x"de00", 366=>x"d300", 367=>x"d300", 368=>x"b300", 369=>x"da00",
---- 370=>x"d700", 371=>x"d200", 372=>x"d600", 373=>x"da00", 374=>x"d400", 375=>x"d600", 376=>x"d600", 377=>x"d300", 378=>x"d300",
---- 379=>x"d500", 380=>x"b000", 381=>x"ac00", 382=>x"d400", 383=>x"d100", 384=>x"a800", 385=>x"cf00", 386=>x"d400", 387=>x"d300",
---- 388=>x"c800", 389=>x"a600", 390=>x"d100", 391=>x"d000", 392=>x"cd00", 393=>x"ae00", 394=>x"6200", 395=>x"d500", 396=>x"d300",
---- 397=>x"b000", 398=>x"2d00", 399=>x"3500", 400=>x"d500", 401=>x"c800", 402=>x"7700", 403=>x"2800", 404=>x"5d00", 405=>x"d600",
---- 406=>x"ae00", 407=>x"4a00", 408=>x"5600", 409=>x"5c00", 410=>x"d800", 411=>x"7d00", 412=>x"5000", 413=>x"5a00", 414=>x"6200",
---- 415=>x"a400", 416=>x"5c00", 417=>x"6400", 418=>x"5c00", 419=>x"6900", 420=>x"9500", 421=>x"5300", 422=>x"5900", 423=>x"6b00",
---- 424=>x"7700", 425=>x"6f00", 426=>x"5f00", 427=>x"5800", 428=>x"6a00", 429=>x"7100", 430=>x"7000", 431=>x"6300", 432=>x"6a00",
---- 433=>x"6c00", 434=>x"6c00", 435=>x"7700", 436=>x"6500", 437=>x"6200", 438=>x"6900", 439=>x"5900", 440=>x"6d00", 441=>x"5f00",
---- 442=>x"5f00", 443=>x"6a00", 444=>x"5600", 445=>x"6300", 446=>x"6000", 447=>x"6100", 448=>x"4900", 449=>x"6100", 450=>x"4d00",
---- 451=>x"6d00", 452=>x"4900", 453=>x"5500", 454=>x"6700", 455=>x"5100", 456=>x"5900", 457=>x"5200", 458=>x"6a00", 459=>x"5c00",
---- 460=>x"5000", 461=>x"4c00", 462=>x"6d00", 463=>x"6300", 464=>x"5500", 465=>x"4300", 466=>x"6200", 467=>x"6900", 468=>x"4d00",
---- 469=>x"4e00", 470=>x"5700", 471=>x"6b00", 472=>x"5300", 473=>x"4800", 474=>x"5200", 475=>x"7000", 476=>x"5a00", 477=>x"4300",
---- 478=>x"4800", 479=>x"6400", 480=>x"5e00", 481=>x"4400", 482=>x"3b00", 483=>x"5d00", 484=>x"7300", 485=>x"4800", 486=>x"4700",
---- 487=>x"4900", 488=>x"7200", 489=>x"7b00", 490=>x"4800", 491=>x"4a00", 492=>x"6a00", 493=>x"8000", 494=>x"7100", 495=>x"5000",
---- 496=>x"6200", 497=>x"8100", 498=>x"7f00", 499=>x"5c00"),
---- 19  => (0=>x"7e00", 1=>x"7a00", 2=>x"7200", 3=>x"8800", 4=>x"af00", 5=>x"7d00", 6=>x"7e00", 7=>x"7e00", 8=>x"7a00", 9=>x"4a00",
---- 10=>x"7c00", 11=>x"8800", 12=>x"7600", 13=>x"3100", 14=>x"2900", 15=>x"8c00", 16=>x"6d00", 17=>x"2800", 18=>x"2a00",
---- 19=>x"2d00", 20=>x"6f00", 21=>x"2a00", 22=>x"5100", 23=>x"4900", 24=>x"2f00", 25=>x"2e00", 26=>x"2d00", 27=>x"2700",
---- 28=>x"3300", 29=>x"3500", 30=>x"5000", 31=>x"3900", 32=>x"3200", 33=>x"2e00", 34=>x"3500", 35=>x"2f00", 36=>x"3800",
---- 37=>x"3100", 38=>x"5500", 39=>x"2c00", 40=>x"3400", 41=>x"3600", 42=>x"3200", 43=>x"2800", 44=>x"2d00", 45=>x"5700",
---- 46=>x"4400", 47=>x"4e00", 48=>x"3e00", 49=>x"2d00", 50=>x"3000", 51=>x"3200", 52=>x"3700", 53=>x"3b00", 54=>x"2a00",
---- 55=>x"3000", 56=>x"3800", 57=>x"4300", 58=>x"2c00", 59=>x"2f00", 60=>x"2a00", 61=>x"3100", 62=>x"2a00", 63=>x"2e00",
---- 64=>x"3500", 65=>x"3200", 66=>x"4e00", 67=>x"2a00", 68=>x"3e00", 69=>x"1c00", 70=>x"2c00", 71=>x"5300", 72=>x"3f00",
---- 73=>x"2800", 74=>x"3d00", 75=>x"2d00", 76=>x"3d00", 77=>x"3b00", 78=>x"2800", 79=>x"9b00", 80=>x"3400", 81=>x"4800",
---- 82=>x"3700", 83=>x"8700", 84=>x"9600", 85=>x"4500", 86=>x"4800", 87=>x"7d00", 88=>x"9c00", 89=>x"8b00", 90=>x"4c00",
---- 91=>x"7700", 92=>x"9200", 93=>x"9000", 94=>x"9900", 95=>x"6f00", 96=>x"9500", 97=>x"9400", 98=>x"9600", 99=>x"a500",
---- 100=>x"9700", 101=>x"8a00", 102=>x"9000", 103=>x"a700", 104=>x"a500", 105=>x"8f00", 106=>x"8a00", 107=>x"a100", 108=>x"a300",
---- 109=>x"9400", 110=>x"8800", 111=>x"a100", 112=>x"a200", 113=>x"9f00", 114=>x"9f00", 115=>x"9f00", 116=>x"a400", 117=>x"9f00",
---- 118=>x"9e00", 119=>x"9d00", 120=>x"9300", 121=>x"9f00", 122=>x"a000", 123=>x"9c00", 124=>x"9f00", 125=>x"9f00", 126=>x"9f00",
---- 127=>x"9000", 128=>x"9d00", 129=>x"9000", 130=>x"9c00", 131=>x"9b00", 132=>x"9d00", 133=>x"9b00", 134=>x"9a00", 135=>x"9d00",
---- 136=>x"9e00", 137=>x"9c00", 138=>x"9b00", 139=>x"9900", 140=>x"9d00", 141=>x"9000", 142=>x"9000", 143=>x"8e00", 144=>x"9b00",
---- 145=>x"9d00", 146=>x"9f00", 147=>x"9e00", 148=>x"9c00", 149=>x"9d00", 150=>x"9d00", 151=>x"9900", 152=>x"9e00", 153=>x"9f00",
---- 154=>x"9c00", 155=>x"9f00", 156=>x"9400", 157=>x"9d00", 158=>x"9d00", 159=>x"9c00", 160=>x"9e00", 161=>x"9700", 162=>x"9f00",
---- 163=>x"9c00", 164=>x"9c00", 165=>x"9c00", 166=>x"9600", 167=>x"8f00", 168=>x"9d00", 169=>x"9a00", 170=>x"9a00", 171=>x"9a00",
---- 172=>x"9c00", 173=>x"8d00", 174=>x"9a00", 175=>x"9b00", 176=>x"9b00", 177=>x"9900", 178=>x"9a00", 179=>x"9a00", 180=>x"9b00",
---- 181=>x"9900", 182=>x"9900", 183=>x"9a00", 184=>x"9100", 185=>x"9b00", 186=>x"9a00", 187=>x"9a00", 188=>x"9b00", 189=>x"9400",
---- 190=>x"9b00", 191=>x"9a00", 192=>x"9a00", 193=>x"9900", 194=>x"9800", 195=>x"9d00", 196=>x"9e00", 197=>x"9b00", 198=>x"9800",
---- 199=>x"9700", 200=>x"a100", 201=>x"8f00", 202=>x"9c00", 203=>x"9a00", 204=>x"9800", 205=>x"9300", 206=>x"9f00", 207=>x"9c00",
---- 208=>x"9900", 209=>x"9700", 210=>x"9f00", 211=>x"9e00", 212=>x"9f00", 213=>x"9b00", 214=>x"9700", 215=>x"9d00", 216=>x"9f00",
---- 217=>x"8f00", 218=>x"9c00", 219=>x"9700", 220=>x"9e00", 221=>x"9b00", 222=>x"9e00", 223=>x"9600", 224=>x"9100", 225=>x"9e00",
---- 226=>x"9a00", 227=>x"9900", 228=>x"9a00", 229=>x"9600", 230=>x"9000", 231=>x"8800", 232=>x"9900", 233=>x"9500", 234=>x"9100",
---- 235=>x"8700", 236=>x"8e00", 237=>x"8d00", 238=>x"9000", 239=>x"9400", 240=>x"9500", 241=>x"8f00", 242=>x"8d00", 243=>x"8500",
---- 244=>x"8600", 245=>x"9d00", 246=>x"8b00", 247=>x"9500", 248=>x"8a00", 249=>x"8400", 250=>x"9a00", 251=>x"9300", 252=>x"9300",
---- 253=>x"8f00", 254=>x"8a00", 255=>x"9200", 256=>x"8f00", 257=>x"8a00", 258=>x"8800", 259=>x"8500", 260=>x"8a00", 261=>x"8800",
---- 262=>x"7e00", 263=>x"7e00", 264=>x"8000", 265=>x"8300", 266=>x"7f00", 267=>x"9000", 268=>x"a600", 269=>x"b100", 270=>x"8a00",
---- 271=>x"a900", 272=>x"ba00", 273=>x"be00", 274=>x"bd00", 275=>x"be00", 276=>x"c300", 277=>x"c000", 278=>x"bd00", 279=>x"bf00",
---- 280=>x"c800", 281=>x"c100", 282=>x"bd00", 283=>x"be00", 284=>x"a400", 285=>x"c400", 286=>x"c100", 287=>x"bd00", 288=>x"c100",
---- 289=>x"c500", 290=>x"c300", 291=>x"c100", 292=>x"c300", 293=>x"c900", 294=>x"cc00", 295=>x"c400", 296=>x"c800", 297=>x"cf00",
---- 298=>x"cd00", 299=>x"ca00", 300=>x"ac00", 301=>x"c900", 302=>x"d200", 303=>x"cd00", 304=>x"cb00", 305=>x"b500", 306=>x"d100",
---- 307=>x"cc00", 308=>x"d100", 309=>x"d000", 310=>x"d100", 311=>x"cd00", 312=>x"cf00", 313=>x"c600", 314=>x"be00", 315=>x"cf00",
---- 316=>x"d400", 317=>x"d700", 318=>x"9600", 319=>x"d800", 320=>x"c700", 321=>x"ad00", 322=>x"d700", 323=>x"ba00", 324=>x"bf00",
---- 325=>x"b900", 326=>x"d600", 327=>x"d100", 328=>x"d400", 329=>x"d800", 330=>x"d300", 331=>x"d100", 332=>x"d400", 333=>x"d400",
---- 334=>x"af00", 335=>x"b700", 336=>x"cc00", 337=>x"d900", 338=>x"d300", 339=>x"d700", 340=>x"ba00", 341=>x"a900", 342=>x"bf00",
---- 343=>x"d700", 344=>x"d500", 345=>x"dc00", 346=>x"d900", 347=>x"d700", 348=>x"d300", 349=>x"d400", 350=>x"bb00", 351=>x"d700",
---- 352=>x"d200", 353=>x"ce00", 354=>x"cc00", 355=>x"b600", 356=>x"c300", 357=>x"b000", 358=>x"d200", 359=>x"c800", 360=>x"d500",
---- 361=>x"cf00", 362=>x"c400", 363=>x"d500", 364=>x"bb00", 365=>x"d300", 366=>x"d100", 367=>x"d000", 368=>x"d300", 369=>x"d400",
---- 370=>x"d200", 371=>x"d100", 372=>x"d400", 373=>x"a500", 374=>x"9500", 375=>x"aa00", 376=>x"b300", 377=>x"6e00", 378=>x"2800",
---- 379=>x"1c00", 380=>x"a900", 381=>x"4000", 382=>x"1b00", 383=>x"2d00", 384=>x"4600", 385=>x"6300", 386=>x"2100", 387=>x"3900",
---- 388=>x"5000", 389=>x"5500", 390=>x"3800", 391=>x"4800", 392=>x"4a00", 393=>x"6800", 394=>x"5500", 395=>x"5600", 396=>x"4e00",
---- 397=>x"5c00", 398=>x"5d00", 399=>x"5100", 400=>x"5a00", 401=>x"5a00", 402=>x"6f00", 403=>x"5c00", 404=>x"5a00", 405=>x"5c00",
---- 406=>x"7100", 407=>x"6d00", 408=>x"5a00", 409=>x"6500", 410=>x"6c00", 411=>x"6c00", 412=>x"5600", 413=>x"6300", 414=>x"6800",
---- 415=>x"7200", 416=>x"5a00", 417=>x"5b00", 418=>x"6800", 419=>x"6400", 420=>x"6c00", 421=>x"5700", 422=>x"6600", 423=>x"6400",
---- 424=>x"6f00", 425=>x"5d00", 426=>x"5f00", 427=>x"6a00", 428=>x"6400", 429=>x"5c00", 430=>x"5800", 431=>x"7000", 432=>x"6600",
---- 433=>x"6b00", 434=>x"5100", 435=>x"5800", 436=>x"6b00", 437=>x"6000", 438=>x"5800", 439=>x"5c00", 440=>x"6a00", 441=>x"6b00",
---- 442=>x"5900", 443=>x"6f00", 444=>x"5e00", 445=>x"6800", 446=>x"5700", 447=>x"5a00", 448=>x"6000", 449=>x"5300", 450=>x"5e00",
---- 451=>x"5900", 452=>x"6900", 453=>x"5b00", 454=>x"3e00", 455=>x"5b00", 456=>x"6200", 457=>x"6400", 458=>x"5a00", 459=>x"3300",
---- 460=>x"5600", 461=>x"6700", 462=>x"5f00", 463=>x"5f00", 464=>x"3000", 465=>x"5b00", 466=>x"7200", 467=>x"5800", 468=>x"4700",
---- 469=>x"3a00", 470=>x"6e00", 471=>x"6400", 472=>x"6a00", 473=>x"4000", 474=>x"4100", 475=>x"7900", 476=>x"6600", 477=>x"4800",
---- 478=>x"4000", 479=>x"4000", 480=>x"7200", 481=>x"6100", 482=>x"4500", 483=>x"3b00", 484=>x"5700", 485=>x"6900", 486=>x"5200",
---- 487=>x"4400", 488=>x"3400", 489=>x"2d00", 490=>x"5800", 491=>x"3a00", 492=>x"3100", 493=>x"5500", 494=>x"4300", 495=>x"3a00",
---- 496=>x"2c00", 497=>x"3200", 498=>x"4800", 499=>x"6500")
---- );
--
--constant c_PIXEL  : t_MATRIX := (
--0   => (0=>x"a200", 1=>x"a100", 2=>x"9f00", 3=>x"9d00", 4=>x"9b00", 5=>x"9e00", 6=>x"9f00", 7=>x"9c00",
--8=>x"a200", 9=>x"a200", 10=>x"a000", 11=>x"a000", 12=>x"a300", 13=>x"a100", 14=>x"9f00",
--15=>x"9f00", 16=>x"a300", 17=>x"a100", 18=>x"a000", 19=>x"a100", 20=>x"a200", 21=>x"9e00",
--22=>x"9e00", 23=>x"9d00", 24=>x"a200", 25=>x"9f00", 26=>x"9e00", 27=>x"9e00", 28=>x"9f00",
--29=>x"a000", 30=>x"9b00", 31=>x"9900", 32=>x"9c00", 33=>x"9d00", 34=>x"9e00", 35=>x"9d00",
--36=>x"9f00", 37=>x"9e00", 38=>x"9d00", 39=>x"9a00", 40=>x"9b00", 41=>x"9d00", 42=>x"9d00",
--43=>x"9700", 44=>x"9d00", 45=>x"9d00", 46=>x"9d00", 47=>x"9c00", 48=>x"9d00", 49=>x"9d00",
--50=>x"9d00", 51=>x"9a00", 52=>x"9d00", 53=>x"9d00", 54=>x"9b00", 55=>x"9c00", 56=>x"9e00",
--57=>x"9e00", 58=>x"9d00", 59=>x"9c00", 60=>x"6300", 61=>x"9b00", 62=>x"9c00", 63=>x"9b00",
--64=>x"9d00", 65=>x"6100", 66=>x"9c00", 67=>x"9a00", 68=>x"9c00", 69=>x"9d00", 70=>x"9c00",
--71=>x"9c00", 72=>x"9c00", 73=>x"9c00", 74=>x"9f00", 75=>x"9a00", 76=>x"9c00", 77=>x"9c00",
--78=>x"9c00", 79=>x"9e00", 80=>x"9b00", 81=>x"9c00", 82=>x"9d00", 83=>x"9c00", 84=>x"9b00",
--85=>x"9d00", 86=>x"9e00", 87=>x"9e00", 88=>x"9e00", 89=>x"9d00", 90=>x"9900", 91=>x"9c00",
--92=>x"9d00", 93=>x"9b00", 94=>x"9e00", 95=>x"9d00", 96=>x"9c00", 97=>x"9a00", 98=>x"9900",
--99=>x"9d00", 100=>x"9f00", 101=>x"9f00", 102=>x"9d00", 103=>x"9e00", 104=>x"9a00", 105=>x"9a00",
--106=>x"9900", 107=>x"9c00", 108=>x"9e00", 109=>x"9f00", 110=>x"9f00", 111=>x"9d00", 112=>x"9e00",
--113=>x"9e00", 114=>x"9d00", 115=>x"9d00", 116=>x"9d00", 117=>x"9f00", 118=>x"9f00", 119=>x"9d00",
--120=>x"9d00", 121=>x"6000", 122=>x"6000", 123=>x"9e00", 124=>x"9f00", 125=>x"6100", 126=>x"a100",
--127=>x"9f00", 128=>x"9d00", 129=>x"9f00", 130=>x"9f00", 131=>x"9c00", 132=>x"9d00", 133=>x"9e00",
--134=>x"a000", 135=>x"a000", 136=>x"9f00", 137=>x"9f00", 138=>x"9d00", 139=>x"9c00", 140=>x"9d00",
--141=>x"9e00", 142=>x"9f00", 143=>x"a100", 144=>x"a000", 145=>x"9d00", 146=>x"9e00", 147=>x"6000",
--148=>x"a100", 149=>x"a400", 150=>x"a300", 151=>x"a100", 152=>x"a100", 153=>x"a000", 154=>x"a100",
--155=>x"6100", 156=>x"a100", 157=>x"a300", 158=>x"a000", 159=>x"a100", 160=>x"a500", 161=>x"a200",
--162=>x"a200", 163=>x"a000", 164=>x"9f00", 165=>x"a200", 166=>x"a200", 167=>x"a100", 168=>x"a000",
--169=>x"a000", 170=>x"a200", 171=>x"a100", 172=>x"9f00", 173=>x"a100", 174=>x"a100", 175=>x"a400",
--176=>x"a100", 177=>x"9f00", 178=>x"a100", 179=>x"a200", 180=>x"a000", 181=>x"a000", 182=>x"a200",
--183=>x"a700", 184=>x"a300", 185=>x"a000", 186=>x"a200", 187=>x"a000", 188=>x"9e00", 189=>x"a100",
--190=>x"a300", 191=>x"5700", 192=>x"a300", 193=>x"a200", 194=>x"a200", 195=>x"a100", 196=>x"9f00",
--197=>x"a200", 198=>x"a600", 199=>x"a900", 200=>x"a200", 201=>x"a300", 202=>x"a000", 203=>x"a000",
--204=>x"9f00", 205=>x"a300", 206=>x"aa00", 207=>x"ac00", 208=>x"a100", 209=>x"9f00", 210=>x"9d00",
--211=>x"a100", 212=>x"a100", 213=>x"a600", 214=>x"aa00", 215=>x"aa00", 216=>x"a100", 217=>x"a200",
--218=>x"a000", 219=>x"a300", 220=>x"a600", 221=>x"a800", 222=>x"a900", 223=>x"a700", 224=>x"9e00",
--225=>x"a000", 226=>x"a000", 227=>x"a400", 228=>x"a800", 229=>x"ab00", 230=>x"a900", 231=>x"a500",
--232=>x"5f00", 233=>x"5f00", 234=>x"a200", 235=>x"a600", 236=>x"aa00", 237=>x"ad00", 238=>x"a700",
--239=>x"a100", 240=>x"a100", 241=>x"a200", 242=>x"a700", 243=>x"aa00", 244=>x"ac00", 245=>x"a800",
--246=>x"a400", 247=>x"9d00", 248=>x"a200", 249=>x"a300", 250=>x"a800", 251=>x"ab00", 252=>x"ab00",
--253=>x"a700", 254=>x"a000", 255=>x"9800", 256=>x"a500", 257=>x"a700", 258=>x"ac00", 259=>x"ae00",
--260=>x"a900", 261=>x"a300", 262=>x"9d00", 263=>x"9600", 264=>x"a700", 265=>x"ab00", 266=>x"b000",
--267=>x"ad00", 268=>x"a700", 269=>x"9f00", 270=>x"9900", 271=>x"9300", 272=>x"a900", 273=>x"ad00",
--274=>x"ae00", 275=>x"aa00", 276=>x"a300", 277=>x"9c00", 278=>x"9600", 279=>x"8b00", 280=>x"ad00",
--281=>x"ac00", 282=>x"ab00", 283=>x"a600", 284=>x"a000", 285=>x"9a00", 286=>x"9200", 287=>x"8300",
--288=>x"ad00", 289=>x"ab00", 290=>x"a900", 291=>x"a400", 292=>x"9e00", 293=>x"9400", 294=>x"8b00",
--295=>x"7e00", 296=>x"ad00", 297=>x"ad00", 298=>x"a700", 299=>x"9f00", 300=>x"9a00", 301=>x"8f00",
--302=>x"8000", 303=>x"7000", 304=>x"aa00", 305=>x"a700", 306=>x"a300", 307=>x"9e00", 308=>x"9500",
--309=>x"8a00", 310=>x"7700", 311=>x"6000", 312=>x"a700", 313=>x"a400", 314=>x"9f00", 315=>x"9900",
--316=>x"8f00", 317=>x"8100", 318=>x"6d00", 319=>x"5200", 320=>x"a200", 321=>x"a200", 322=>x"6600",
--323=>x"9300", 324=>x"8600", 325=>x"7600", 326=>x"6100", 327=>x"5100", 328=>x"a200", 329=>x"9f00",
--330=>x"9700", 331=>x"8c00", 332=>x"7b00", 333=>x"6a00", 334=>x"5500", 335=>x"5000", 336=>x"9b00",
--337=>x"9900", 338=>x"9200", 339=>x"8400", 340=>x"8e00", 341=>x"5e00", 342=>x"4f00", 343=>x"5200",
--344=>x"9700", 345=>x"9400", 346=>x"8900", 347=>x"7700", 348=>x"6200", 349=>x"5100", 350=>x"5300",
--351=>x"5600", 352=>x"9400", 353=>x"8d00", 354=>x"7e00", 355=>x"6a00", 356=>x"5700", 357=>x"5100",
--358=>x"5600", 359=>x"5900", 360=>x"8b00", 361=>x"7900", 362=>x"7300", 363=>x"5d00", 364=>x"5300",
--365=>x"5400", 366=>x"5800", 367=>x"5800", 368=>x"8300", 369=>x"7c00", 370=>x"6700", 371=>x"5500",
--372=>x"5400", 373=>x"5700", 374=>x"5d00", 375=>x"5900", 376=>x"7b00", 377=>x"6f00", 378=>x"5800",
--379=>x"5300", 380=>x"5500", 381=>x"5b00", 382=>x"6000", 383=>x"5c00", 384=>x"6d00", 385=>x"6100",
--386=>x"5100", 387=>x"5500", 388=>x"5700", 389=>x"a500", 390=>x"5b00", 391=>x"5b00", 392=>x"6100",
--393=>x"5700", 394=>x"5400", 395=>x"5600", 396=>x"5700", 397=>x"5b00", 398=>x"6000", 399=>x"5d00",
--400=>x"5800", 401=>x"5400", 402=>x"5500", 403=>x"5b00", 404=>x"5800", 405=>x"5900", 406=>x"5c00",
--407=>x"5800", 408=>x"5b00", 409=>x"5800", 410=>x"5600", 411=>x"5c00", 412=>x"5d00", 413=>x"5b00",
--414=>x"5b00", 415=>x"5d00", 416=>x"5500", 417=>x"5700", 418=>x"5900", 419=>x"5d00", 420=>x"5d00",
--421=>x"5b00", 422=>x"5d00", 423=>x"5d00", 424=>x"5600", 425=>x"5400", 426=>x"5500", 427=>x"5d00",
--428=>x"5d00", 429=>x"5c00", 430=>x"5d00", 431=>x"5f00", 432=>x"5b00", 433=>x"5900", 434=>x"5a00",
--435=>x"5e00", 436=>x"5c00", 437=>x"5c00", 438=>x"5b00", 439=>x"5a00", 440=>x"5b00", 441=>x"5b00",
--442=>x"5a00", 443=>x"5d00", 444=>x"5e00", 445=>x"5a00", 446=>x"5b00", 447=>x"5d00", 448=>x"5c00",
--449=>x"5f00", 450=>x"5a00", 451=>x"5b00", 452=>x"5c00", 453=>x"5c00", 454=>x"5d00", 455=>x"5d00",
--456=>x"5c00", 457=>x"5f00", 458=>x"5b00", 459=>x"5900", 460=>x"5b00", 461=>x"5900", 462=>x"5700",
--463=>x"5900", 464=>x"5700", 465=>x"5900", 466=>x"5a00", 467=>x"5a00", 468=>x"5a00", 469=>x"5900",
--470=>x"5600", 471=>x"5900", 472=>x"5d00", 473=>x"5a00", 474=>x"a700", 475=>x"5a00", 476=>x"5800",
--477=>x"5700", 478=>x"5800", 479=>x"5a00", 480=>x"5900", 481=>x"5900", 482=>x"5900", 483=>x"5900",
--484=>x"5a00", 485=>x"5c00", 486=>x"5b00", 487=>x"5b00", 488=>x"5700", 489=>x"5700", 490=>x"5900",
--491=>x"5900", 492=>x"5c00", 493=>x"5a00", 494=>x"5c00", 495=>x"5e00", 496=>x"5c00", 497=>x"5b00",
--498=>x"5a00", 499=>x"5d00"),
--1  => (0=>x"9b00", 1=>x"a000", 2=>x"9d00", 3=>x"9b00", 4=>x"9c00", 5=>x"9a00", 6=>x"9a00", 7=>x"9b00",
--8=>x"9b00", 9=>x"a200", 10=>x"9c00", 11=>x"9a00", 12=>x"9c00", 13=>x"9900", 14=>x"9a00",
--15=>x"9900", 16=>x"9a00", 17=>x"9f00", 18=>x"9b00", 19=>x"9a00", 20=>x"9c00", 21=>x"9a00",
--22=>x"9a00", 23=>x"9a00", 24=>x"9b00", 25=>x"9b00", 26=>x"9a00", 27=>x"9700", 28=>x"9a00",
--29=>x"9a00", 30=>x"9800", 31=>x"9a00", 32=>x"9b00", 33=>x"9c00", 34=>x"9b00", 35=>x"9a00",
--36=>x"9b00", 37=>x"9a00", 38=>x"9800", 39=>x"9a00", 40=>x"9b00", 41=>x"9b00", 42=>x"9d00",
--43=>x"9c00", 44=>x"9800", 45=>x"9900", 46=>x"9c00", 47=>x"9a00", 48=>x"9e00", 49=>x"9d00",
--50=>x"9c00", 51=>x"9c00", 52=>x"9a00", 53=>x"9900", 54=>x"6400", 55=>x"6400", 56=>x"9d00",
--57=>x"9c00", 58=>x"9b00", 59=>x"9a00", 60=>x"9a00", 61=>x"9a00", 62=>x"9b00", 63=>x"9c00",
--64=>x"9a00", 65=>x"9c00", 66=>x"9c00", 67=>x"9b00", 68=>x"9900", 69=>x"9800", 70=>x"9a00",
--71=>x"a100", 72=>x"9d00", 73=>x"9f00", 74=>x"9c00", 75=>x"9b00", 76=>x"9b00", 77=>x"9900",
--78=>x"9d00", 79=>x"a100", 80=>x"9f00", 81=>x"9f00", 82=>x"9b00", 83=>x"9c00", 84=>x"9b00",
--85=>x"9b00", 86=>x"9e00", 87=>x"a000", 88=>x"9f00", 89=>x"9e00", 90=>x"9c00", 91=>x"9c00",
--92=>x"9800", 93=>x"9b00", 94=>x"9c00", 95=>x"a200", 96=>x"9f00", 97=>x"9c00", 98=>x"9c00",
--99=>x"9e00", 100=>x"9d00", 101=>x"9e00", 102=>x"a100", 103=>x"a400", 104=>x"9e00", 105=>x"9f00",
--106=>x"9e00", 107=>x"9c00", 108=>x"9d00", 109=>x"a100", 110=>x"a300", 111=>x"a600", 112=>x"9f00",
--113=>x"9f00", 114=>x"9f00", 115=>x"9e00", 116=>x"9e00", 117=>x"a200", 118=>x"a700", 119=>x"a800",
--120=>x"9e00", 121=>x"a000", 122=>x"a000", 123=>x"a100", 124=>x"a300", 125=>x"a700", 126=>x"a700",
--127=>x"a800", 128=>x"9f00", 129=>x"a200", 130=>x"a000", 131=>x"a300", 132=>x"a700", 133=>x"a800",
--134=>x"a800", 135=>x"aa00", 136=>x"a100", 137=>x"a100", 138=>x"a300", 139=>x"a500", 140=>x"a800",
--141=>x"a700", 142=>x"a800", 143=>x"a800", 144=>x"a300", 145=>x"a400", 146=>x"a500", 147=>x"a700",
--148=>x"a800", 149=>x"a800", 150=>x"a800", 151=>x"a900", 152=>x"a300", 153=>x"5900", 154=>x"a800",
--155=>x"a900", 156=>x"a700", 157=>x"a800", 158=>x"a700", 159=>x"a400", 160=>x"a400", 161=>x"a700",
--162=>x"a900", 163=>x"a700", 164=>x"a500", 165=>x"a400", 166=>x"5e00", 167=>x"a200", 168=>x"a800",
--169=>x"a900", 170=>x"a900", 171=>x"a200", 172=>x"a200", 173=>x"a200", 174=>x"9e00", 175=>x"a100",
--176=>x"ab00", 177=>x"ab00", 178=>x"a700", 179=>x"a000", 180=>x"9c00", 181=>x"9e00", 182=>x"9a00",
--183=>x"9d00", 184=>x"a900", 185=>x"a500", 186=>x"a000", 187=>x"9c00", 188=>x"9a00", 189=>x"9a00",
--190=>x"9900", 191=>x"9700", 192=>x"ab00", 193=>x"a400", 194=>x"9e00", 195=>x"6500", 196=>x"9700",
--197=>x"9500", 198=>x"9400", 199=>x"9500", 200=>x"a900", 201=>x"a200", 202=>x"9c00", 203=>x"9600",
--204=>x"9200", 205=>x"6e00", 206=>x"8e00", 207=>x"9100", 208=>x"a800", 209=>x"a000", 210=>x"9900",
--211=>x"6d00", 212=>x"8c00", 213=>x"8c00", 214=>x"8d00", 215=>x"8a00", 216=>x"a300", 217=>x"9f00",
--218=>x"9500", 219=>x"8f00", 220=>x"8700", 221=>x"8200", 222=>x"8700", 223=>x"8a00", 224=>x"9e00",
--225=>x"9900", 226=>x"9000", 227=>x"8700", 228=>x"8100", 229=>x"7e00", 230=>x"8000", 231=>x"8a00",
--232=>x"9b00", 233=>x"9300", 234=>x"8b00", 235=>x"7e00", 236=>x"7900", 237=>x"7800", 238=>x"8000",
--239=>x"8f00", 240=>x"9800", 241=>x"8f00", 242=>x"7f00", 243=>x"7300", 244=>x"6d00", 245=>x"6f00",
--246=>x"8000", 247=>x"9000", 248=>x"6a00", 249=>x"8700", 250=>x"7700", 251=>x"6800", 252=>x"6100",
--253=>x"7000", 254=>x"8100", 255=>x"8d00", 256=>x"8f00", 257=>x"7d00", 258=>x"6b00", 259=>x"5c00",
--260=>x"5a00", 261=>x"7000", 262=>x"8000", 263=>x"8e00", 264=>x"8800", 265=>x"7400", 266=>x"6100",
--267=>x"4f00", 268=>x"5900", 269=>x"7000", 270=>x"8100", 271=>x"8e00", 272=>x"7f00", 273=>x"6900",
--274=>x"5300", 275=>x"4a00", 276=>x"5700", 277=>x"6f00", 278=>x"8200", 279=>x"8e00", 280=>x"7100",
--281=>x"5600", 282=>x"4a00", 283=>x"4c00", 284=>x"5a00", 285=>x"7200", 286=>x"8000", 287=>x"8a00",
--288=>x"6600", 289=>x"5000", 290=>x"b600", 291=>x"5000", 292=>x"6000", 293=>x"6e00", 294=>x"8000",
--295=>x"8c00", 296=>x"5700", 297=>x"4d00", 298=>x"4d00", 299=>x"ae00", 300=>x"6000", 301=>x"7200",
--302=>x"8000", 303=>x"8c00", 304=>x"5300", 305=>x"5300", 306=>x"4c00", 307=>x"5100", 308=>x"5f00",
--309=>x"7400", 310=>x"8100", 311=>x"8b00", 312=>x"5400", 313=>x"5700", 314=>x"5100", 315=>x"4f00",
--316=>x"5e00", 317=>x"7100", 318=>x"8200", 319=>x"8c00", 320=>x"5200", 321=>x"5300", 322=>x"5600",
--323=>x"5200", 324=>x"6000", 325=>x"7400", 326=>x"8200", 327=>x"8e00", 328=>x"5300", 329=>x"5400",
--330=>x"5200", 331=>x"5500", 332=>x"5f00", 333=>x"7300", 334=>x"8400", 335=>x"8e00", 336=>x"5600",
--337=>x"5500", 338=>x"5300", 339=>x"5700", 340=>x"6000", 341=>x"7200", 342=>x"7f00", 343=>x"8d00",
--344=>x"5900", 345=>x"5b00", 346=>x"5400", 347=>x"5700", 348=>x"5f00", 349=>x"7000", 350=>x"8000",
--351=>x"8d00", 352=>x"5b00", 353=>x"5900", 354=>x"5300", 355=>x"5600", 356=>x"6300", 357=>x"8d00",
--358=>x"8200", 359=>x"7200", 360=>x"5800", 361=>x"5700", 362=>x"5600", 363=>x"5700", 364=>x"9f00",
--365=>x"7000", 366=>x"7f00", 367=>x"8e00", 368=>x"5900", 369=>x"5700", 370=>x"5800", 371=>x"5600",
--372=>x"5d00", 373=>x"7000", 374=>x"7e00", 375=>x"8c00", 376=>x"5900", 377=>x"5900", 378=>x"5600",
--379=>x"5500", 380=>x"5d00", 381=>x"6e00", 382=>x"8000", 383=>x"8c00", 384=>x"5b00", 385=>x"5800",
--386=>x"5400", 387=>x"5600", 388=>x"5d00", 389=>x"6f00", 390=>x"8200", 391=>x"8c00", 392=>x"5b00",
--393=>x"5b00", 394=>x"5500", 395=>x"5600", 396=>x"6000", 397=>x"6e00", 398=>x"7e00", 399=>x"8700",
--400=>x"5c00", 401=>x"5b00", 402=>x"5600", 403=>x"5500", 404=>x"5e00", 405=>x"6c00", 406=>x"7b00",
--407=>x"8900", 408=>x"5c00", 409=>x"5a00", 410=>x"5700", 411=>x"5800", 412=>x"5f00", 413=>x"6d00",
--414=>x"7d00", 415=>x"8c00", 416=>x"5a00", 417=>x"5b00", 418=>x"5700", 419=>x"5a00", 420=>x"6100",
--421=>x"6e00", 422=>x"8000", 423=>x"8b00", 424=>x"5d00", 425=>x"5a00", 426=>x"5900", 427=>x"5b00",
--428=>x"6300", 429=>x"7100", 430=>x"8000", 431=>x"8a00", 432=>x"5b00", 433=>x"5b00", 434=>x"5900",
--435=>x"5700", 436=>x"5f00", 437=>x"7100", 438=>x"7f00", 439=>x"8a00", 440=>x"5c00", 441=>x"5700",
--442=>x"5600", 443=>x"5700", 444=>x"5c00", 445=>x"6f00", 446=>x"7d00", 447=>x"8c00", 448=>x"5b00",
--449=>x"5a00", 450=>x"5700", 451=>x"5500", 452=>x"5c00", 453=>x"6a00", 454=>x"7d00", 455=>x"8d00",
--456=>x"5600", 457=>x"5500", 458=>x"5400", 459=>x"5300", 460=>x"5c00", 461=>x"6b00", 462=>x"8000",
--463=>x"8c00", 464=>x"a300", 465=>x"5900", 466=>x"5400", 467=>x"5400", 468=>x"a600", 469=>x"6a00",
--470=>x"7a00", 471=>x"8800", 472=>x"5b00", 473=>x"5800", 474=>x"5300", 475=>x"5400", 476=>x"5600",
--477=>x"6900", 478=>x"7b00", 479=>x"8800", 480=>x"5c00", 481=>x"5b00", 482=>x"5800", 483=>x"5400",
--484=>x"5b00", 485=>x"6c00", 486=>x"7d00", 487=>x"8700", 488=>x"6000", 489=>x"5c00", 490=>x"5900",
--491=>x"5900", 492=>x"5b00", 493=>x"6d00", 494=>x"7c00", 495=>x"8600", 496=>x"6100", 497=>x"5b00",
--498=>x"5a00", 499=>x"5600"),
--2  => (0=>x"9b00", 1=>x"9c00", 2=>x"a000", 3=>x"a400", 4=>x"a600", 5=>x"a700", 6=>x"ae00", 7=>x"ad00",
--8=>x"9b00", 9=>x"9c00", 10=>x"5d00", 11=>x"a400", 12=>x"a600", 13=>x"a700", 14=>x"ad00",
--15=>x"ad00", 16=>x"9c00", 17=>x"9b00", 18=>x"9f00", 19=>x"a300", 20=>x"a400", 21=>x"a700",
--22=>x"ac00", 23=>x"ad00", 24=>x"9d00", 25=>x"9900", 26=>x"9c00", 27=>x"a200", 28=>x"a600",
--29=>x"a900", 30=>x"ab00", 31=>x"ac00", 32=>x"9b00", 33=>x"9a00", 34=>x"a100", 35=>x"a400",
--36=>x"a800", 37=>x"ab00", 38=>x"ac00", 39=>x"ac00", 40=>x"9900", 41=>x"9d00", 42=>x"a100",
--43=>x"a600", 44=>x"a800", 45=>x"a800", 46=>x"ab00", 47=>x"ab00", 48=>x"9b00", 49=>x"a000",
--50=>x"a300", 51=>x"a600", 52=>x"a900", 53=>x"a900", 54=>x"a900", 55=>x"a800", 56=>x"9f00",
--57=>x"a300", 58=>x"a700", 59=>x"a800", 60=>x"a900", 61=>x"a800", 62=>x"a900", 63=>x"a800",
--64=>x"a200", 65=>x"a500", 66=>x"a800", 67=>x"a600", 68=>x"a700", 69=>x"a900", 70=>x"a500",
--71=>x"a700", 72=>x"a200", 73=>x"a700", 74=>x"a700", 75=>x"a600", 76=>x"a700", 77=>x"a400",
--78=>x"a600", 79=>x"a400", 80=>x"a400", 81=>x"a600", 82=>x"a400", 83=>x"a500", 84=>x"a700",
--85=>x"a400", 86=>x"a500", 87=>x"a200", 88=>x"a600", 89=>x"a600", 90=>x"a500", 91=>x"a200",
--92=>x"a600", 93=>x"a500", 94=>x"a400", 95=>x"a300", 96=>x"a700", 97=>x"a600", 98=>x"a800",
--99=>x"a500", 100=>x"5b00", 101=>x"a400", 102=>x"a300", 103=>x"9f00", 104=>x"a600", 105=>x"a700",
--106=>x"a600", 107=>x"5900", 108=>x"a100", 109=>x"a100", 110=>x"a100", 111=>x"9e00", 112=>x"a800",
--113=>x"a800", 114=>x"a600", 115=>x"a400", 116=>x"a000", 117=>x"9e00", 118=>x"9e00", 119=>x"9e00",
--120=>x"a900", 121=>x"a700", 122=>x"a600", 123=>x"a300", 124=>x"a000", 125=>x"9f00", 126=>x"9d00",
--127=>x"9d00", 128=>x"aa00", 129=>x"a700", 130=>x"a700", 131=>x"a200", 132=>x"9f00", 133=>x"9f00",
--134=>x"9e00", 135=>x"9e00", 136=>x"a700", 137=>x"a700", 138=>x"a900", 139=>x"a100", 140=>x"a000",
--141=>x"a100", 142=>x"9d00", 143=>x"9e00", 144=>x"a600", 145=>x"a600", 146=>x"a500", 147=>x"a000",
--148=>x"9c00", 149=>x"9e00", 150=>x"9e00", 151=>x"9f00", 152=>x"a500", 153=>x"a300", 154=>x"a200",
--155=>x"a100", 156=>x"9e00", 157=>x"9e00", 158=>x"a000", 159=>x"a100", 160=>x"a400", 161=>x"a300",
--162=>x"a000", 163=>x"a000", 164=>x"9f00", 165=>x"9f00", 166=>x"a100", 167=>x"a100", 168=>x"a000",
--169=>x"9c00", 170=>x"a000", 171=>x"a300", 172=>x"a000", 173=>x"9e00", 174=>x"a000", 175=>x"a000",
--176=>x"9c00", 177=>x"9c00", 178=>x"9d00", 179=>x"a200", 180=>x"a100", 181=>x"9f00", 182=>x"9f00",
--183=>x"9f00", 184=>x"9a00", 185=>x"9b00", 186=>x"a000", 187=>x"a400", 188=>x"a500", 189=>x"a300",
--190=>x"a000", 191=>x"a100", 192=>x"9500", 193=>x"9a00", 194=>x"a100", 195=>x"a200", 196=>x"a200",
--197=>x"a100", 198=>x"9f00", 199=>x"a100", 200=>x"9200", 201=>x"6500", 202=>x"a100", 203=>x"a600",
--204=>x"a300", 205=>x"a100", 206=>x"a100", 207=>x"a100", 208=>x"9000", 209=>x"9a00", 210=>x"a300",
--211=>x"a400", 212=>x"a400", 213=>x"a200", 214=>x"a200", 215=>x"a200", 216=>x"9100", 217=>x"9b00",
--218=>x"a200", 219=>x"a300", 220=>x"a400", 221=>x"a200", 222=>x"a200", 223=>x"5c00", 224=>x"9400",
--225=>x"9b00", 226=>x"a300", 227=>x"a600", 228=>x"a400", 229=>x"a300", 230=>x"a200", 231=>x"a600",
--232=>x"9700", 233=>x"9d00", 234=>x"a300", 235=>x"a400", 236=>x"a500", 237=>x"a600", 238=>x"a400",
--239=>x"a400", 240=>x"9700", 241=>x"9d00", 242=>x"a400", 243=>x"a800", 244=>x"a400", 245=>x"a700",
--246=>x"a400", 247=>x"a300", 248=>x"9800", 249=>x"9d00", 250=>x"a500", 251=>x"a800", 252=>x"a500",
--253=>x"a500", 254=>x"a600", 255=>x"a500", 256=>x"9900", 257=>x"9f00", 258=>x"a500", 259=>x"a700",
--260=>x"a600", 261=>x"a500", 262=>x"a400", 263=>x"a500", 264=>x"9900", 265=>x"a100", 266=>x"a600",
--267=>x"a600", 268=>x"a500", 269=>x"a600", 270=>x"a900", 271=>x"a300", 272=>x"9600", 273=>x"a200",
--274=>x"a400", 275=>x"a800", 276=>x"a700", 277=>x"a400", 278=>x"a500", 279=>x"a300", 280=>x"9400",
--281=>x"a000", 282=>x"a700", 283=>x"a600", 284=>x"a800", 285=>x"a400", 286=>x"a400", 287=>x"a600",
--288=>x"9600", 289=>x"9f00", 290=>x"a400", 291=>x"a800", 292=>x"ab00", 293=>x"a600", 294=>x"a600",
--295=>x"a500", 296=>x"9800", 297=>x"5f00", 298=>x"a600", 299=>x"a900", 300=>x"a700", 301=>x"a600",
--302=>x"5900", 303=>x"a400", 304=>x"9800", 305=>x"a000", 306=>x"a600", 307=>x"a700", 308=>x"a600",
--309=>x"a800", 310=>x"a700", 311=>x"a400", 312=>x"9700", 313=>x"9e00", 314=>x"a400", 315=>x"a800",
--316=>x"a800", 317=>x"a900", 318=>x"a800", 319=>x"a600", 320=>x"9700", 321=>x"9d00", 322=>x"a500",
--323=>x"a600", 324=>x"a800", 325=>x"a800", 326=>x"a700", 327=>x"a700", 328=>x"9700", 329=>x"9d00",
--330=>x"a400", 331=>x"a700", 332=>x"a700", 333=>x"a700", 334=>x"a900", 335=>x"a700", 336=>x"9700",
--337=>x"9c00", 338=>x"a300", 339=>x"a800", 340=>x"a800", 341=>x"a800", 342=>x"5700", 343=>x"a600",
--344=>x"9600", 345=>x"9f00", 346=>x"a500", 347=>x"a800", 348=>x"a700", 349=>x"a800", 350=>x"a700",
--351=>x"a600", 352=>x"9600", 353=>x"9f00", 354=>x"a400", 355=>x"a600", 356=>x"a800", 357=>x"a600",
--358=>x"a600", 359=>x"a500", 360=>x"9400", 361=>x"9b00", 362=>x"a200", 363=>x"a600", 364=>x"a700",
--365=>x"a800", 366=>x"a400", 367=>x"a600", 368=>x"9600", 369=>x"9c00", 370=>x"a200", 371=>x"a500",
--372=>x"a500", 373=>x"a800", 374=>x"a600", 375=>x"a400", 376=>x"9500", 377=>x"9c00", 378=>x"a000",
--379=>x"a400", 380=>x"a700", 381=>x"a700", 382=>x"a600", 383=>x"a600", 384=>x"9300", 385=>x"9b00",
--386=>x"a000", 387=>x"a500", 388=>x"a500", 389=>x"a700", 390=>x"a800", 391=>x"a700", 392=>x"9400",
--393=>x"9a00", 394=>x"a100", 395=>x"a400", 396=>x"a500", 397=>x"a700", 398=>x"a500", 399=>x"a600",
--400=>x"9300", 401=>x"9b00", 402=>x"a000", 403=>x"a300", 404=>x"a600", 405=>x"a600", 406=>x"a500",
--407=>x"a500", 408=>x"9300", 409=>x"9c00", 410=>x"a100", 411=>x"a700", 412=>x"a500", 413=>x"a500",
--414=>x"a800", 415=>x"a700", 416=>x"9300", 417=>x"9b00", 418=>x"9f00", 419=>x"a200", 420=>x"a600",
--421=>x"a600", 422=>x"a700", 423=>x"a600", 424=>x"9200", 425=>x"9b00", 426=>x"9f00", 427=>x"a400",
--428=>x"a400", 429=>x"a200", 430=>x"a400", 431=>x"a600", 432=>x"9400", 433=>x"9d00", 434=>x"9e00",
--435=>x"a200", 436=>x"a500", 437=>x"a300", 438=>x"a300", 439=>x"a300", 440=>x"9400", 441=>x"9c00",
--442=>x"a000", 443=>x"a200", 444=>x"a500", 445=>x"a500", 446=>x"a600", 447=>x"a300", 448=>x"9100",
--449=>x"9900", 450=>x"9f00", 451=>x"a400", 452=>x"a500", 453=>x"a500", 454=>x"a500", 455=>x"a400",
--456=>x"9500", 457=>x"9a00", 458=>x"9f00", 459=>x"a200", 460=>x"a500", 461=>x"a300", 462=>x"a300",
--463=>x"a200", 464=>x"9300", 465=>x"9c00", 466=>x"a000", 467=>x"a300", 468=>x"a600", 469=>x"a300",
--470=>x"a400", 471=>x"a400", 472=>x"9200", 473=>x"9b00", 474=>x"a000", 475=>x"a400", 476=>x"a300",
--477=>x"a500", 478=>x"a400", 479=>x"a200", 480=>x"9000", 481=>x"9b00", 482=>x"a000", 483=>x"a300",
--484=>x"a500", 485=>x"a400", 486=>x"a400", 487=>x"a300", 488=>x"9000", 489=>x"9900", 490=>x"a000",
--491=>x"a200", 492=>x"a500", 493=>x"a700", 494=>x"a700", 495=>x"a600", 496=>x"9300", 497=>x"9900",
--498=>x"9f00", 499=>x"a500"),
--3  => (0=>x"ab00", 1=>x"ab00", 2=>x"a900", 3=>x"a200", 4=>x"9700", 5=>x"9600", 6=>x"8200", 7=>x"7300",
--8=>x"5400", 9=>x"ab00", 10=>x"a900", 11=>x"a300", 12=>x"9700", 13=>x"9700", 14=>x"8300",
--15=>x"7200", 16=>x"ab00", 17=>x"ac00", 18=>x"a900", 19=>x"a200", 20=>x"9800", 21=>x"9500",
--22=>x"8000", 23=>x"7000", 24=>x"ad00", 25=>x"ab00", 26=>x"a600", 27=>x"a000", 28=>x"9700",
--29=>x"8b00", 30=>x"7c00", 31=>x"7100", 32=>x"ac00", 33=>x"a900", 34=>x"a600", 35=>x"9e00",
--36=>x"9500", 37=>x"8b00", 38=>x"7d00", 39=>x"7300", 40=>x"aa00", 41=>x"a900", 42=>x"a700",
--43=>x"9d00", 44=>x"9100", 45=>x"8800", 46=>x"8000", 47=>x"7000", 48=>x"a800", 49=>x"a700",
--50=>x"a600", 51=>x"9d00", 52=>x"8e00", 53=>x"8900", 54=>x"7d00", 55=>x"6c00", 56=>x"a700",
--57=>x"a500", 58=>x"9f00", 59=>x"9b00", 60=>x"9300", 61=>x"8800", 62=>x"7d00", 63=>x"7200",
--64=>x"a600", 65=>x"a300", 66=>x"9f00", 67=>x"9b00", 68=>x"9000", 69=>x"8800", 70=>x"7c00",
--71=>x"6d00", 72=>x"a500", 73=>x"a300", 74=>x"9e00", 75=>x"9800", 76=>x"9000", 77=>x"8a00",
--78=>x"7f00", 79=>x"6f00", 80=>x"a200", 81=>x"a300", 82=>x"9d00", 83=>x"9a00", 84=>x"9100",
--85=>x"8b00", 86=>x"8400", 87=>x"7900", 88=>x"9f00", 89=>x"a100", 90=>x"9f00", 91=>x"9a00",
--92=>x"9300", 93=>x"8900", 94=>x"8200", 95=>x"7100", 96=>x"9f00", 97=>x"a200", 98=>x"9f00",
--99=>x"9900", 100=>x"9500", 101=>x"8b00", 102=>x"8000", 103=>x"7200", 104=>x"a000", 105=>x"a100",
--106=>x"a000", 107=>x"9900", 108=>x"9400", 109=>x"8b00", 110=>x"7b00", 111=>x"6c00", 112=>x"a000",
--113=>x"a200", 114=>x"a100", 115=>x"9c00", 116=>x"9400", 117=>x"8a00", 118=>x"7b00", 119=>x"6d00",
--120=>x"a000", 121=>x"a400", 122=>x"a300", 123=>x"a000", 124=>x"9400", 125=>x"8900", 126=>x"7e00",
--127=>x"6e00", 128=>x"a000", 129=>x"a100", 130=>x"a100", 131=>x"9d00", 132=>x"9600", 133=>x"8c00",
--134=>x"8000", 135=>x"6f00", 136=>x"a000", 137=>x"a300", 138=>x"a200", 139=>x"9b00", 140=>x"9300",
--141=>x"8800", 142=>x"7c00", 143=>x"6c00", 144=>x"9f00", 145=>x"a100", 146=>x"a100", 147=>x"9c00",
--148=>x"9200", 149=>x"8700", 150=>x"7f00", 151=>x"6d00", 152=>x"5d00", 153=>x"a100", 154=>x"a000",
--155=>x"9a00", 156=>x"9100", 157=>x"8900", 158=>x"7f00", 159=>x"6d00", 160=>x"a100", 161=>x"a100",
--162=>x"9f00", 163=>x"9b00", 164=>x"9400", 165=>x"8700", 166=>x"7b00", 167=>x"6900", 168=>x"5f00",
--169=>x"a100", 170=>x"a000", 171=>x"9a00", 172=>x"9100", 173=>x"8900", 174=>x"7b00", 175=>x"6900",
--176=>x"a000", 177=>x"a200", 178=>x"a000", 179=>x"9900", 180=>x"9400", 181=>x"8900", 182=>x"7c00",
--183=>x"6a00", 184=>x"a200", 185=>x"a400", 186=>x"a100", 187=>x"9a00", 188=>x"9500", 189=>x"8b00",
--190=>x"7d00", 191=>x"6b00", 192=>x"a400", 193=>x"5d00", 194=>x"a000", 195=>x"9c00", 196=>x"9500",
--197=>x"8a00", 198=>x"8200", 199=>x"7000", 200=>x"a400", 201=>x"a400", 202=>x"a100", 203=>x"9c00",
--204=>x"9500", 205=>x"8900", 206=>x"8100", 207=>x"6c00", 208=>x"a500", 209=>x"a400", 210=>x"a200",
--211=>x"9b00", 212=>x"9300", 213=>x"8a00", 214=>x"7f00", 215=>x"6c00", 216=>x"a600", 217=>x"a400",
--218=>x"a200", 219=>x"9d00", 220=>x"9100", 221=>x"8d00", 222=>x"7e00", 223=>x"6c00", 224=>x"a600",
--225=>x"a500", 226=>x"a400", 227=>x"9f00", 228=>x"9500", 229=>x"8b00", 230=>x"8000", 231=>x"6c00",
--232=>x"a500", 233=>x"a400", 234=>x"a000", 235=>x"9c00", 236=>x"6900", 237=>x"8b00", 238=>x"7e00",
--239=>x"6800", 240=>x"a400", 241=>x"a500", 242=>x"a100", 243=>x"9f00", 244=>x"9600", 245=>x"8d00",
--246=>x"8000", 247=>x"6b00", 248=>x"a600", 249=>x"a500", 250=>x"a300", 251=>x"9d00", 252=>x"9600",
--253=>x"8b00", 254=>x"8000", 255=>x"6e00", 256=>x"a600", 257=>x"a600", 258=>x"a400", 259=>x"9d00",
--260=>x"9600", 261=>x"8b00", 262=>x"7d00", 263=>x"6a00", 264=>x"a300", 265=>x"a300", 266=>x"a200",
--267=>x"9b00", 268=>x"9400", 269=>x"8b00", 270=>x"7e00", 271=>x"6d00", 272=>x"a300", 273=>x"a300",
--274=>x"a100", 275=>x"9a00", 276=>x"9100", 277=>x"8800", 278=>x"7f00", 279=>x"6b00", 280=>x"a600",
--281=>x"a500", 282=>x"a000", 283=>x"9b00", 284=>x"8f00", 285=>x"8800", 286=>x"7d00", 287=>x"6b00",
--288=>x"a200", 289=>x"a200", 290=>x"a000", 291=>x"9a00", 292=>x"9100", 293=>x"8900", 294=>x"7c00",
--295=>x"6a00", 296=>x"a500", 297=>x"a300", 298=>x"a000", 299=>x"9900", 300=>x"9200", 301=>x"8700",
--302=>x"8200", 303=>x"6c00", 304=>x"a400", 305=>x"a300", 306=>x"a000", 307=>x"9900", 308=>x"9300",
--309=>x"8900", 310=>x"7a00", 311=>x"6700", 312=>x"a300", 313=>x"a100", 314=>x"a000", 315=>x"9c00",
--316=>x"9400", 317=>x"8a00", 318=>x"7b00", 319=>x"6b00", 320=>x"a400", 321=>x"a300", 322=>x"5f00",
--323=>x"9a00", 324=>x"9300", 325=>x"8900", 326=>x"7900", 327=>x"6800", 328=>x"a600", 329=>x"a300",
--330=>x"9f00", 331=>x"9a00", 332=>x"9100", 333=>x"8600", 334=>x"7900", 335=>x"6700", 336=>x"a600",
--337=>x"a200", 338=>x"9d00", 339=>x"9800", 340=>x"8f00", 341=>x"8600", 342=>x"7500", 343=>x"6b00",
--344=>x"a600", 345=>x"a500", 346=>x"9e00", 347=>x"9800", 348=>x"9000", 349=>x"8600", 350=>x"7900",
--351=>x"6a00", 352=>x"a800", 353=>x"a500", 354=>x"9e00", 355=>x"9800", 356=>x"9000", 357=>x"8300",
--358=>x"7c00", 359=>x"6b00", 360=>x"a700", 361=>x"a400", 362=>x"9f00", 363=>x"9800", 364=>x"9000",
--365=>x"8400", 366=>x"7700", 367=>x"6a00", 368=>x"a400", 369=>x"a300", 370=>x"a000", 371=>x"9a00",
--372=>x"9000", 373=>x"8500", 374=>x"7900", 375=>x"6800", 376=>x"a600", 377=>x"a200", 378=>x"9f00",
--379=>x"9b00", 380=>x"9100", 381=>x"8400", 382=>x"7600", 383=>x"6700", 384=>x"a300", 385=>x"a400",
--386=>x"9e00", 387=>x"9a00", 388=>x"9200", 389=>x"8800", 390=>x"7800", 391=>x"6c00", 392=>x"a200",
--393=>x"a200", 394=>x"a000", 395=>x"9900", 396=>x"8e00", 397=>x"8500", 398=>x"7a00", 399=>x"6800",
--400=>x"a600", 401=>x"a300", 402=>x"a100", 403=>x"9800", 404=>x"9000", 405=>x"8600", 406=>x"7800",
--407=>x"6a00", 408=>x"a600", 409=>x"a300", 410=>x"a000", 411=>x"9a00", 412=>x"9100", 413=>x"8500",
--414=>x"7a00", 415=>x"6b00", 416=>x"a400", 417=>x"a300", 418=>x"9f00", 419=>x"6500", 420=>x"9200",
--421=>x"8600", 422=>x"7a00", 423=>x"6800", 424=>x"a000", 425=>x"a200", 426=>x"9f00", 427=>x"9a00",
--428=>x"9200", 429=>x"8900", 430=>x"7900", 431=>x"6900", 432=>x"a300", 433=>x"a300", 434=>x"a100",
--435=>x"9c00", 436=>x"6f00", 437=>x"8800", 438=>x"7900", 439=>x"6a00", 440=>x"a200", 441=>x"a400",
--442=>x"a400", 443=>x"9b00", 444=>x"9300", 445=>x"8800", 446=>x"7b00", 447=>x"6a00", 448=>x"a300",
--449=>x"a500", 450=>x"a400", 451=>x"9d00", 452=>x"9200", 453=>x"8700", 454=>x"7800", 455=>x"6c00",
--456=>x"a300", 457=>x"a300", 458=>x"a400", 459=>x"9b00", 460=>x"9200", 461=>x"8900", 462=>x"7d00",
--463=>x"7000", 464=>x"a300", 465=>x"a200", 466=>x"a100", 467=>x"9900", 468=>x"9300", 469=>x"8600",
--470=>x"7b00", 471=>x"6c00", 472=>x"a200", 473=>x"a400", 474=>x"a100", 475=>x"9a00", 476=>x"9100",
--477=>x"8800", 478=>x"7800", 479=>x"6800", 480=>x"a400", 481=>x"a500", 482=>x"a200", 483=>x"9a00",
--484=>x"9100", 485=>x"8600", 486=>x"7a00", 487=>x"6a00", 488=>x"a300", 489=>x"a200", 490=>x"a000",
--491=>x"9c00", 492=>x"9300", 493=>x"8600", 494=>x"7b00", 495=>x"6500", 496=>x"a400", 497=>x"a400",
--498=>x"a100", 499=>x"9a00"),
--4  => (0=>x"6300", 1=>x"5d00", 2=>x"5b00", 3=>x"6400", 4=>x"6400", 5=>x"6700", 6=>x"6900", 7=>x"6900",
--8=>x"6300", 9=>x"5e00", 10=>x"5b00", 11=>x"6500", 12=>x"6400", 13=>x"6700", 14=>x"6900",
--15=>x"6900", 16=>x"6400", 17=>x"5e00", 18=>x"5c00", 19=>x"6300", 20=>x"9c00", 21=>x"6600",
--22=>x"6900", 23=>x"6900", 24=>x"6300", 25=>x"5b00", 26=>x"5a00", 27=>x"5e00", 28=>x"6100",
--29=>x"6000", 30=>x"6900", 31=>x"6c00", 32=>x"6300", 33=>x"5a00", 34=>x"5800", 35=>x"5a00",
--36=>x"5f00", 37=>x"6400", 38=>x"6600", 39=>x"6800", 40=>x"6000", 41=>x"5b00", 42=>x"5900",
--43=>x"5b00", 44=>x"6200", 45=>x"6100", 46=>x"6300", 47=>x"6700", 48=>x"6300", 49=>x"5900",
--50=>x"5900", 51=>x"5b00", 52=>x"5d00", 53=>x"6000", 54=>x"6300", 55=>x"6900", 56=>x"6400",
--57=>x"5a00", 58=>x"5c00", 59=>x"5b00", 60=>x"5d00", 61=>x"6500", 62=>x"6500", 63=>x"6600",
--64=>x"6100", 65=>x"5900", 66=>x"5700", 67=>x"5b00", 68=>x"5c00", 69=>x"6500", 70=>x"9700",
--71=>x"6200", 72=>x"6100", 73=>x"5b00", 74=>x"5700", 75=>x"5d00", 76=>x"5f00", 77=>x"6400",
--78=>x"6600", 79=>x"6200", 80=>x"6600", 81=>x"a300", 82=>x"5700", 83=>x"5d00", 84=>x"5e00",
--85=>x"6100", 86=>x"6700", 87=>x"6700", 88=>x"6100", 89=>x"5a00", 90=>x"5b00", 91=>x"5f00",
--92=>x"6100", 93=>x"6200", 94=>x"6400", 95=>x"6600", 96=>x"6300", 97=>x"5800", 98=>x"5600",
--99=>x"5d00", 100=>x"6000", 101=>x"6000", 102=>x"6300", 103=>x"6800", 104=>x"5c00", 105=>x"5800",
--106=>x"5200", 107=>x"5600", 108=>x"5d00", 109=>x"6000", 110=>x"6500", 111=>x"6700", 112=>x"5f00",
--113=>x"5700", 114=>x"5500", 115=>x"5700", 116=>x"5f00", 117=>x"6200", 118=>x"6400", 119=>x"6700",
--120=>x"6100", 121=>x"5a00", 122=>x"5600", 123=>x"5a00", 124=>x"6100", 125=>x"6200", 126=>x"6200",
--127=>x"6800", 128=>x"6100", 129=>x"5a00", 130=>x"5700", 131=>x"5e00", 132=>x"5f00", 133=>x"6000",
--134=>x"6400", 135=>x"6400", 136=>x"5f00", 137=>x"5800", 138=>x"5a00", 139=>x"5d00", 140=>x"5f00",
--141=>x"6400", 142=>x"6200", 143=>x"6700", 144=>x"6000", 145=>x"5600", 146=>x"5600", 147=>x"5a00",
--148=>x"6100", 149=>x"6100", 150=>x"6500", 151=>x"6600", 152=>x"5b00", 153=>x"5300", 154=>x"5300",
--155=>x"5700", 156=>x"5f00", 157=>x"5f00", 158=>x"6400", 159=>x"6500", 160=>x"5d00", 161=>x"5400",
--162=>x"5100", 163=>x"5b00", 164=>x"5e00", 165=>x"6000", 166=>x"6800", 167=>x"6800", 168=>x"5d00",
--169=>x"5400", 170=>x"5300", 171=>x"5900", 172=>x"5c00", 173=>x"6200", 174=>x"6700", 175=>x"6700",
--176=>x"5d00", 177=>x"5300", 178=>x"5300", 179=>x"5b00", 180=>x"5e00", 181=>x"6200", 182=>x"6400",
--183=>x"6500", 184=>x"5e00", 185=>x"5400", 186=>x"5100", 187=>x"5b00", 188=>x"5d00", 189=>x"5f00",
--190=>x"6200", 191=>x"6600", 192=>x"6100", 193=>x"5800", 194=>x"5300", 195=>x"5900", 196=>x"5e00",
--197=>x"6000", 198=>x"6200", 199=>x"6500", 200=>x"5c00", 201=>x"5600", 202=>x"5500", 203=>x"5900",
--204=>x"5c00", 205=>x"6000", 206=>x"6100", 207=>x"6300", 208=>x"5e00", 209=>x"5200", 210=>x"ae00",
--211=>x"5700", 212=>x"5e00", 213=>x"5c00", 214=>x"6200", 215=>x"6500", 216=>x"5c00", 217=>x"5100",
--218=>x"5500", 219=>x"5800", 220=>x"5d00", 221=>x"5e00", 222=>x"6300", 223=>x"6200", 224=>x"5900",
--225=>x"4f00", 226=>x"5000", 227=>x"5600", 228=>x"5600", 229=>x"5b00", 230=>x"6000", 231=>x"6000",
--232=>x"5900", 233=>x"4c00", 234=>x"4e00", 235=>x"5300", 236=>x"5a00", 237=>x"5f00", 238=>x"9c00",
--239=>x"6000", 240=>x"a600", 241=>x"5100", 242=>x"4e00", 243=>x"5300", 244=>x"5f00", 245=>x"5b00",
--246=>x"5e00", 247=>x"6100", 248=>x"5900", 249=>x"5200", 250=>x"4d00", 251=>x"5000", 252=>x"5700",
--253=>x"5600", 254=>x"5a00", 255=>x"5c00", 256=>x"5a00", 257=>x"4c00", 258=>x"4c00", 259=>x"5100",
--260=>x"5300", 261=>x"5600", 262=>x"5b00", 263=>x"5e00", 264=>x"5700", 265=>x"4b00", 266=>x"4900",
--267=>x"5100", 268=>x"5200", 269=>x"5700", 270=>x"5b00", 271=>x"5d00", 272=>x"5900", 273=>x"4e00",
--274=>x"4700", 275=>x"5000", 276=>x"5200", 277=>x"5a00", 278=>x"5e00", 279=>x"5d00", 280=>x"5500",
--281=>x"4b00", 282=>x"4700", 283=>x"5000", 284=>x"5700", 285=>x"5800", 286=>x"5900", 287=>x"5d00",
--288=>x"5300", 289=>x"4b00", 290=>x"4800", 291=>x"5000", 292=>x"5600", 293=>x"5800", 294=>x"5b00",
--295=>x"5f00", 296=>x"5300", 297=>x"4b00", 298=>x"4800", 299=>x"5000", 300=>x"5600", 301=>x"5a00",
--302=>x"5e00", 303=>x"6000", 304=>x"5400", 305=>x"4900", 306=>x"4b00", 307=>x"5100", 308=>x"5400",
--309=>x"5800", 310=>x"5c00", 311=>x"6000", 312=>x"5700", 313=>x"4a00", 314=>x"4e00", 315=>x"5100",
--316=>x"5800", 317=>x"5600", 318=>x"5c00", 319=>x"6200", 320=>x"5600", 321=>x"4d00", 322=>x"4700",
--323=>x"5000", 324=>x"5500", 325=>x"5900", 326=>x"5f00", 327=>x"6100", 328=>x"5400", 329=>x"4d00",
--330=>x"4a00", 331=>x"5000", 332=>x"5800", 333=>x"5a00", 334=>x"5e00", 335=>x"5f00", 336=>x"5900",
--337=>x"4c00", 338=>x"4a00", 339=>x"5000", 340=>x"5600", 341=>x"5a00", 342=>x"6100", 343=>x"5f00",
--344=>x"5b00", 345=>x"5000", 346=>x"4f00", 347=>x"5300", 348=>x"5800", 349=>x"5a00", 350=>x"5c00",
--351=>x"5c00", 352=>x"5900", 353=>x"4f00", 354=>x"4a00", 355=>x"5000", 356=>x"5500", 357=>x"5b00",
--358=>x"5c00", 359=>x"5e00", 360=>x"5800", 361=>x"4b00", 362=>x"4900", 363=>x"5200", 364=>x"5800",
--365=>x"5b00", 366=>x"5d00", 367=>x"6200", 368=>x"5a00", 369=>x"4c00", 370=>x"4b00", 371=>x"5300",
--372=>x"5800", 373=>x"5a00", 374=>x"6000", 375=>x"6100", 376=>x"a500", 377=>x"4d00", 378=>x"4e00",
--379=>x"5200", 380=>x"5800", 381=>x"5f00", 382=>x"6200", 383=>x"6100", 384=>x"5c00", 385=>x"4900",
--386=>x"4e00", 387=>x"5300", 388=>x"5900", 389=>x"5b00", 390=>x"6200", 391=>x"5d00", 392=>x"5a00",
--393=>x"4d00", 394=>x"4c00", 395=>x"4d00", 396=>x"5600", 397=>x"5c00", 398=>x"6000", 399=>x"6100",
--400=>x"5900", 401=>x"4c00", 402=>x"4b00", 403=>x"4d00", 404=>x"5600", 405=>x"5900", 406=>x"5e00",
--407=>x"6100", 408=>x"5e00", 409=>x"4e00", 410=>x"b700", 411=>x"4f00", 412=>x"5600", 413=>x"5800",
--414=>x"5e00", 415=>x"5f00", 416=>x"5e00", 417=>x"4e00", 418=>x"4900", 419=>x"5000", 420=>x"5500",
--421=>x"5a00", 422=>x"5e00", 423=>x"5e00", 424=>x"5900", 425=>x"5000", 426=>x"4c00", 427=>x"4e00",
--428=>x"5500", 429=>x"5b00", 430=>x"5e00", 431=>x"5f00", 432=>x"5e00", 433=>x"4f00", 434=>x"4b00",
--435=>x"5100", 436=>x"5500", 437=>x"5a00", 438=>x"5c00", 439=>x"5b00", 440=>x"a400", 441=>x"4e00",
--442=>x"4a00", 443=>x"5200", 444=>x"5500", 445=>x"5400", 446=>x"5a00", 447=>x"5d00", 448=>x"5900",
--449=>x"4c00", 450=>x"4a00", 451=>x"5100", 452=>x"5600", 453=>x"5600", 454=>x"5c00", 455=>x"6000",
--456=>x"5c00", 457=>x"5000", 458=>x"4b00", 459=>x"5000", 460=>x"5400", 461=>x"5a00", 462=>x"5d00",
--463=>x"5f00", 464=>x"5c00", 465=>x"4900", 466=>x"4700", 467=>x"4f00", 468=>x"5000", 469=>x"5600",
--470=>x"5800", 471=>x"5800", 472=>x"5600", 473=>x"4600", 474=>x"4700", 475=>x"4f00", 476=>x"5300",
--477=>x"5500", 478=>x"5800", 479=>x"5800", 480=>x"5300", 481=>x"4800", 482=>x"4600", 483=>x"4b00",
--484=>x"4f00", 485=>x"5300", 486=>x"5900", 487=>x"5c00", 488=>x"5600", 489=>x"4700", 490=>x"4500",
--491=>x"4a00", 492=>x"4d00", 493=>x"5200", 494=>x"5b00", 495=>x"5f00", 496=>x"5500", 497=>x"4d00",
--498=>x"4900", 499=>x"4c00"),
--5  => (0=>x"6d00", 1=>x"6a00", 2=>x"6900", 3=>x"6d00", 4=>x"6c00", 5=>x"6a00", 6=>x"6d00", 7=>x"6c00",
--8=>x"6e00", 9=>x"6a00", 10=>x"6900", 11=>x"6e00", 12=>x"6c00", 13=>x"6b00", 14=>x"6d00",
--15=>x"6b00", 16=>x"6d00", 17=>x"6a00", 18=>x"6800", 19=>x"6c00", 20=>x"6b00", 21=>x"6a00",
--22=>x"6d00", 23=>x"6b00", 24=>x"6700", 25=>x"6800", 26=>x"6700", 27=>x"6800", 28=>x"6700",
--29=>x"6800", 30=>x"6900", 31=>x"6800", 32=>x"9500", 33=>x"6900", 34=>x"6500", 35=>x"6a00",
--36=>x"6900", 37=>x"6800", 38=>x"6800", 39=>x"6700", 40=>x"9b00", 41=>x"6600", 42=>x"6700",
--43=>x"6700", 44=>x"6800", 45=>x"6b00", 46=>x"6700", 47=>x"6600", 48=>x"6600", 49=>x"6900",
--50=>x"6a00", 51=>x"6b00", 52=>x"6c00", 53=>x"6900", 54=>x"6600", 55=>x"6700", 56=>x"6900",
--57=>x"6e00", 58=>x"6b00", 59=>x"6b00", 60=>x"6b00", 61=>x"6b00", 62=>x"6600", 63=>x"6800",
--64=>x"6a00", 65=>x"6a00", 66=>x"6900", 67=>x"6a00", 68=>x"6700", 69=>x"9700", 70=>x"6700",
--71=>x"6a00", 72=>x"6600", 73=>x"6700", 74=>x"6a00", 75=>x"6b00", 76=>x"6900", 77=>x"6a00",
--78=>x"6900", 79=>x"6a00", 80=>x"6b00", 81=>x"6c00", 82=>x"6b00", 83=>x"6c00", 84=>x"6800",
--85=>x"6800", 86=>x"6600", 87=>x"6500", 88=>x"7000", 89=>x"6700", 90=>x"6700", 91=>x"6700",
--92=>x"6700", 93=>x"9500", 94=>x"6500", 95=>x"6600", 96=>x"6a00", 97=>x"6800", 98=>x"6900",
--99=>x"6600", 100=>x"6400", 101=>x"6a00", 102=>x"6700", 103=>x"6800", 104=>x"6900", 105=>x"6900",
--106=>x"6900", 107=>x"6900", 108=>x"6900", 109=>x"6a00", 110=>x"6600", 111=>x"6600", 112=>x"6700",
--113=>x"6800", 114=>x"6800", 115=>x"6b00", 116=>x"6a00", 117=>x"6900", 118=>x"6800", 119=>x"6700",
--120=>x"6b00", 121=>x"6b00", 122=>x"6c00", 123=>x"6700", 124=>x"6900", 125=>x"6a00", 126=>x"6600",
--127=>x"6700", 128=>x"6900", 129=>x"6b00", 130=>x"6c00", 131=>x"6c00", 132=>x"6b00", 133=>x"6a00",
--134=>x"6400", 135=>x"6600", 136=>x"6800", 137=>x"6900", 138=>x"6800", 139=>x"6a00", 140=>x"6900",
--141=>x"6700", 142=>x"6700", 143=>x"6700", 144=>x"6800", 145=>x"6700", 146=>x"6600", 147=>x"6500",
--148=>x"6700", 149=>x"6700", 150=>x"6700", 151=>x"6400", 152=>x"6600", 153=>x"6900", 154=>x"6500",
--155=>x"6500", 156=>x"6600", 157=>x"6800", 158=>x"6600", 159=>x"6600", 160=>x"6700", 161=>x"6700",
--162=>x"6400", 163=>x"6700", 164=>x"6600", 165=>x"6500", 166=>x"6500", 167=>x"6700", 168=>x"6700",
--169=>x"9a00", 170=>x"6600", 171=>x"6700", 172=>x"6600", 173=>x"6a00", 174=>x"6400", 175=>x"9800",
--176=>x"6700", 177=>x"6600", 178=>x"6900", 179=>x"6700", 180=>x"6700", 181=>x"6800", 182=>x"6a00",
--183=>x"6600", 184=>x"6800", 185=>x"6900", 186=>x"6900", 187=>x"6b00", 188=>x"6700", 189=>x"6600",
--190=>x"6900", 191=>x"6700", 192=>x"6700", 193=>x"6900", 194=>x"6900", 195=>x"6c00", 196=>x"6700",
--197=>x"6600", 198=>x"6800", 199=>x"6600", 200=>x"6700", 201=>x"6700", 202=>x"6600", 203=>x"6700",
--204=>x"6600", 205=>x"6400", 206=>x"6700", 207=>x"6900", 208=>x"6800", 209=>x"6900", 210=>x"6700",
--211=>x"6800", 212=>x"6600", 213=>x"6a00", 214=>x"6700", 215=>x"6600", 216=>x"6500", 217=>x"6900",
--218=>x"6500", 219=>x"6500", 220=>x"6800", 221=>x"6900", 222=>x"6600", 223=>x"6700", 224=>x"6300",
--225=>x"6400", 226=>x"6800", 227=>x"6300", 228=>x"6600", 229=>x"6600", 230=>x"6700", 231=>x"6500",
--232=>x"5f00", 233=>x"6100", 234=>x"6300", 235=>x"6600", 236=>x"6500", 237=>x"6300", 238=>x"9b00",
--239=>x"6200", 240=>x"6500", 241=>x"6500", 242=>x"6400", 243=>x"9d00", 244=>x"6300", 245=>x"6500",
--246=>x"6100", 247=>x"6400", 248=>x"6100", 249=>x"6400", 250=>x"6100", 251=>x"5f00", 252=>x"6300",
--253=>x"6200", 254=>x"6200", 255=>x"6500", 256=>x"5f00", 257=>x"5e00", 258=>x"5d00", 259=>x"6200",
--260=>x"6400", 261=>x"6300", 262=>x"6300", 263=>x"6300", 264=>x"5e00", 265=>x"5f00", 266=>x"5f00",
--267=>x"6200", 268=>x"6100", 269=>x"6300", 270=>x"6400", 271=>x"6500", 272=>x"5f00", 273=>x"6100",
--274=>x"6200", 275=>x"6100", 276=>x"6200", 277=>x"6500", 278=>x"6300", 279=>x"6300", 280=>x"6400",
--281=>x"6700", 282=>x"6600", 283=>x"6900", 284=>x"6300", 285=>x"6500", 286=>x"6500", 287=>x"6300",
--288=>x"6400", 289=>x"6500", 290=>x"6000", 291=>x"6700", 292=>x"6600", 293=>x"6400", 294=>x"6100",
--295=>x"9d00", 296=>x"6100", 297=>x"6200", 298=>x"6100", 299=>x"6600", 300=>x"6400", 301=>x"6600",
--302=>x"9c00", 303=>x"6300", 304=>x"6500", 305=>x"6200", 306=>x"6200", 307=>x"6400", 308=>x"6200",
--309=>x"6400", 310=>x"6300", 311=>x"6500", 312=>x"6900", 313=>x"6200", 314=>x"6300", 315=>x"6400",
--316=>x"9b00", 317=>x"6100", 318=>x"6500", 319=>x"6200", 320=>x"6100", 321=>x"6000", 322=>x"6000",
--323=>x"6100", 324=>x"6600", 325=>x"6400", 326=>x"6200", 327=>x"6400", 328=>x"5f00", 329=>x"6500",
--330=>x"6900", 331=>x"6000", 332=>x"6400", 333=>x"6500", 334=>x"6300", 335=>x"6300", 336=>x"6100",
--337=>x"6300", 338=>x"6300", 339=>x"6300", 340=>x"6300", 341=>x"6000", 342=>x"6800", 343=>x"6700",
--344=>x"6000", 345=>x"6300", 346=>x"6300", 347=>x"6300", 348=>x"6200", 349=>x"6400", 350=>x"6a00",
--351=>x"6700", 352=>x"5f00", 353=>x"5e00", 354=>x"6200", 355=>x"6600", 356=>x"6600", 357=>x"6600",
--358=>x"6900", 359=>x"6500", 360=>x"5f00", 361=>x"5e00", 362=>x"6500", 363=>x"6700", 364=>x"6500",
--365=>x"6500", 366=>x"6900", 367=>x"6600", 368=>x"6100", 369=>x"5f00", 370=>x"6200", 371=>x"6300",
--372=>x"6200", 373=>x"6300", 374=>x"6500", 375=>x"9c00", 376=>x"6700", 377=>x"6200", 378=>x"6100",
--379=>x"6100", 380=>x"6300", 381=>x"6200", 382=>x"6600", 383=>x"9e00", 384=>x"6400", 385=>x"6600",
--386=>x"6100", 387=>x"6300", 388=>x"6400", 389=>x"6400", 390=>x"6300", 391=>x"6600", 392=>x"6300",
--393=>x"6300", 394=>x"6300", 395=>x"6500", 396=>x"6200", 397=>x"6100", 398=>x"6200", 399=>x"6200",
--400=>x"6000", 401=>x"6600", 402=>x"6300", 403=>x"6400", 404=>x"6200", 405=>x"6500", 406=>x"6100",
--407=>x"6400", 408=>x"6200", 409=>x"6200", 410=>x"6200", 411=>x"6100", 412=>x"6200", 413=>x"6600",
--414=>x"6300", 415=>x"6400", 416=>x"6100", 417=>x"6000", 418=>x"6000", 419=>x"6600", 420=>x"6700",
--421=>x"6500", 422=>x"6300", 423=>x"6300", 424=>x"5f00", 425=>x"6000", 426=>x"6100", 427=>x"6100",
--428=>x"6900", 429=>x"6600", 430=>x"6300", 431=>x"6200", 432=>x"6000", 433=>x"6200", 434=>x"6400",
--435=>x"6200", 436=>x"6500", 437=>x"6400", 438=>x"6600", 439=>x"6400", 440=>x"5f00", 441=>x"6300",
--442=>x"6300", 443=>x"6200", 444=>x"6500", 445=>x"6400", 446=>x"6500", 447=>x"6600", 448=>x"5e00",
--449=>x"6100", 450=>x"5d00", 451=>x"6200", 452=>x"6400", 453=>x"6600", 454=>x"6a00", 455=>x"6500",
--456=>x"5c00", 457=>x"5d00", 458=>x"6100", 459=>x"6300", 460=>x"6500", 461=>x"6200", 462=>x"6600",
--463=>x"6300", 464=>x"5c00", 465=>x"5f00", 466=>x"5f00", 467=>x"5f00", 468=>x"6100", 469=>x"6000",
--470=>x"5f00", 471=>x"6000", 472=>x"5e00", 473=>x"5d00", 474=>x"5f00", 475=>x"6000", 476=>x"5f00",
--477=>x"6100", 478=>x"6000", 479=>x"5e00", 480=>x"5d00", 481=>x"6100", 482=>x"6200", 483=>x"6200",
--484=>x"6100", 485=>x"6200", 486=>x"6200", 487=>x"5f00", 488=>x"5b00", 489=>x"5e00", 490=>x"6200",
--491=>x"6200", 492=>x"6200", 493=>x"6500", 494=>x"6300", 495=>x"6300", 496=>x"5e00", 497=>x"6200",
--498=>x"6400", 499=>x"6300"),
--6  => (0=>x"6d00", 1=>x"6d00", 2=>x"6800", 3=>x"6a00", 4=>x"9200", 5=>x"7000", 6=>x"7100", 7=>x"7800",
--8=>x"6f00", 9=>x"6d00", 10=>x"6900", 11=>x"6a00", 12=>x"6e00", 13=>x"7200", 14=>x"7100",
--15=>x"7800", 16=>x"6c00", 17=>x"6c00", 18=>x"6900", 19=>x"6800", 20=>x"6d00", 21=>x"7200",
--22=>x"7200", 23=>x"7700", 24=>x"6a00", 25=>x"6a00", 26=>x"6800", 27=>x"6b00", 28=>x"6b00",
--29=>x"6e00", 30=>x"7400", 31=>x"7500", 32=>x"6700", 33=>x"6a00", 34=>x"6800", 35=>x"6b00",
--36=>x"6e00", 37=>x"6e00", 38=>x"7000", 39=>x"7400", 40=>x"6800", 41=>x"6600", 42=>x"6700",
--43=>x"6c00", 44=>x"6e00", 45=>x"6d00", 46=>x"7200", 47=>x"7400", 48=>x"6700", 49=>x"6700",
--50=>x"6500", 51=>x"6700", 52=>x"7000", 53=>x"8f00", 54=>x"7100", 55=>x"7400", 56=>x"6900",
--57=>x"6500", 58=>x"6600", 59=>x"6800", 60=>x"6e00", 61=>x"6e00", 62=>x"7000", 63=>x"7400",
--64=>x"6700", 65=>x"6800", 66=>x"6500", 67=>x"6700", 68=>x"6b00", 69=>x"6f00", 70=>x"7000",
--71=>x"7400", 72=>x"6500", 73=>x"6700", 74=>x"6600", 75=>x"6900", 76=>x"9200", 77=>x"7100",
--78=>x"7300", 79=>x"7500", 80=>x"6900", 81=>x"6800", 82=>x"6600", 83=>x"6500", 84=>x"6e00",
--85=>x"7100", 86=>x"7300", 87=>x"7100", 88=>x"6600", 89=>x"6700", 90=>x"6700", 91=>x"6900",
--92=>x"6d00", 93=>x"6f00", 94=>x"6f00", 95=>x"7300", 96=>x"6600", 97=>x"6600", 98=>x"6800",
--99=>x"6b00", 100=>x"6b00", 101=>x"6e00", 102=>x"6f00", 103=>x"6f00", 104=>x"6800", 105=>x"6600",
--106=>x"6700", 107=>x"6c00", 108=>x"6e00", 109=>x"6d00", 110=>x"6f00", 111=>x"7200", 112=>x"6700",
--113=>x"6500", 114=>x"6800", 115=>x"6b00", 116=>x"6b00", 117=>x"6c00", 118=>x"7100", 119=>x"7300",
--120=>x"6900", 121=>x"6600", 122=>x"6600", 123=>x"6b00", 124=>x"6c00", 125=>x"6b00", 126=>x"6e00",
--127=>x"7300", 128=>x"6700", 129=>x"6500", 130=>x"6800", 131=>x"6a00", 132=>x"6b00", 133=>x"6e00",
--134=>x"7100", 135=>x"7100", 136=>x"6400", 137=>x"6500", 138=>x"6600", 139=>x"6800", 140=>x"6b00",
--141=>x"6f00", 142=>x"6f00", 143=>x"7200", 144=>x"6600", 145=>x"6800", 146=>x"6800", 147=>x"6900",
--148=>x"6b00", 149=>x"6e00", 150=>x"7200", 151=>x"7000", 152=>x"6600", 153=>x"6900", 154=>x"6500",
--155=>x"6800", 156=>x"6b00", 157=>x"6e00", 158=>x"7000", 159=>x"7300", 160=>x"6600", 161=>x"6600",
--162=>x"6600", 163=>x"6700", 164=>x"6900", 165=>x"6f00", 166=>x"7200", 167=>x"7400", 168=>x"6500",
--169=>x"6500", 170=>x"6700", 171=>x"6700", 172=>x"6900", 173=>x"6d00", 174=>x"6f00", 175=>x"7100",
--176=>x"6700", 177=>x"6500", 178=>x"6700", 179=>x"6800", 180=>x"6d00", 181=>x"6c00", 182=>x"6f00",
--183=>x"7400", 184=>x"6600", 185=>x"6600", 186=>x"6800", 187=>x"6900", 188=>x"7000", 189=>x"6c00",
--190=>x"7200", 191=>x"7500", 192=>x"6500", 193=>x"6500", 194=>x"6700", 195=>x"6a00", 196=>x"6f00",
--197=>x"7000", 198=>x"7000", 199=>x"6f00", 200=>x"6700", 201=>x"6500", 202=>x"6700", 203=>x"6a00",
--204=>x"6e00", 205=>x"7200", 206=>x"7100", 207=>x"7100", 208=>x"6900", 209=>x"6900", 210=>x"6a00",
--211=>x"6d00", 212=>x"6c00", 213=>x"6f00", 214=>x"7100", 215=>x"7400", 216=>x"6a00", 217=>x"6700",
--218=>x"6800", 219=>x"6b00", 220=>x"6d00", 221=>x"7100", 222=>x"7700", 223=>x"7300", 224=>x"6800",
--225=>x"6800", 226=>x"6900", 227=>x"6800", 228=>x"6c00", 229=>x"6f00", 230=>x"7700", 231=>x"7300",
--232=>x"6200", 233=>x"6a00", 234=>x"6c00", 235=>x"9600", 236=>x"6a00", 237=>x"6e00", 238=>x"7100",
--239=>x"7100", 240=>x"6500", 241=>x"6800", 242=>x"6800", 243=>x"6a00", 244=>x"6b00", 245=>x"6e00",
--246=>x"7000", 247=>x"7100", 248=>x"9800", 249=>x"6400", 250=>x"6700", 251=>x"6900", 252=>x"6b00",
--253=>x"6e00", 254=>x"6e00", 255=>x"7200", 256=>x"6400", 257=>x"6600", 258=>x"6900", 259=>x"6800",
--260=>x"6900", 261=>x"6d00", 262=>x"6c00", 263=>x"6f00", 264=>x"6400", 265=>x"6600", 266=>x"6800",
--267=>x"6700", 268=>x"6700", 269=>x"6a00", 270=>x"6600", 271=>x"6d00", 272=>x"6500", 273=>x"6600",
--274=>x"6300", 275=>x"6400", 276=>x"6900", 277=>x"6a00", 278=>x"6c00", 279=>x"6f00", 280=>x"6500",
--281=>x"6500", 282=>x"6700", 283=>x"6800", 284=>x"6b00", 285=>x"6c00", 286=>x"6c00", 287=>x"6f00",
--288=>x"6400", 289=>x"6500", 290=>x"6100", 291=>x"6400", 292=>x"6800", 293=>x"6b00", 294=>x"6d00",
--295=>x"6d00", 296=>x"6300", 297=>x"6300", 298=>x"6300", 299=>x"6700", 300=>x"6900", 301=>x"6a00",
--302=>x"6d00", 303=>x"6d00", 304=>x"6400", 305=>x"6400", 306=>x"6600", 307=>x"6600", 308=>x"6800",
--309=>x"6800", 310=>x"6c00", 311=>x"6e00", 312=>x"6500", 313=>x"6500", 314=>x"6500", 315=>x"6800",
--316=>x"6700", 317=>x"6a00", 318=>x"6e00", 319=>x"7000", 320=>x"6700", 321=>x"6600", 322=>x"9b00",
--323=>x"6700", 324=>x"6a00", 325=>x"6c00", 326=>x"6d00", 327=>x"6e00", 328=>x"6400", 329=>x"6500",
--330=>x"6600", 331=>x"6800", 332=>x"6900", 333=>x"6b00", 334=>x"6e00", 335=>x"6e00", 336=>x"6300",
--337=>x"6500", 338=>x"6500", 339=>x"6700", 340=>x"6600", 341=>x"6900", 342=>x"7000", 343=>x"7000",
--344=>x"6600", 345=>x"6400", 346=>x"6400", 347=>x"6600", 348=>x"6700", 349=>x"6a00", 350=>x"6b00",
--351=>x"6e00", 352=>x"6600", 353=>x"6300", 354=>x"6500", 355=>x"6600", 356=>x"6900", 357=>x"6d00",
--358=>x"9200", 359=>x"6c00", 360=>x"6400", 361=>x"6400", 362=>x"6300", 363=>x"6500", 364=>x"6b00",
--365=>x"6e00", 366=>x"6c00", 367=>x"6c00", 368=>x"6200", 369=>x"6200", 370=>x"6600", 371=>x"6700",
--372=>x"6a00", 373=>x"6600", 374=>x"6b00", 375=>x"6e00", 376=>x"6600", 377=>x"6300", 378=>x"6300",
--379=>x"6a00", 380=>x"6900", 381=>x"6700", 382=>x"6b00", 383=>x"6e00", 384=>x"6500", 385=>x"6500",
--386=>x"6400", 387=>x"6800", 388=>x"6500", 389=>x"6700", 390=>x"6b00", 391=>x"6f00", 392=>x"6300",
--393=>x"6300", 394=>x"6700", 395=>x"6800", 396=>x"9800", 397=>x"6a00", 398=>x"6900", 399=>x"6d00",
--400=>x"6300", 401=>x"6600", 402=>x"6800", 403=>x"6600", 404=>x"6700", 405=>x"6a00", 406=>x"6e00",
--407=>x"6d00", 408=>x"6500", 409=>x"6800", 410=>x"6400", 411=>x"6600", 412=>x"6600", 413=>x"6a00",
--414=>x"6d00", 415=>x"6f00", 416=>x"6400", 417=>x"6600", 418=>x"6200", 419=>x"6500", 420=>x"6700",
--421=>x"6900", 422=>x"6d00", 423=>x"6e00", 424=>x"6200", 425=>x"6100", 426=>x"6600", 427=>x"6300",
--428=>x"6700", 429=>x"6a00", 430=>x"6b00", 431=>x"6e00", 432=>x"6200", 433=>x"6300", 434=>x"6500",
--435=>x"6500", 436=>x"6700", 437=>x"6800", 438=>x"6a00", 439=>x"6e00", 440=>x"9b00", 441=>x"6400",
--442=>x"6500", 443=>x"6400", 444=>x"6b00", 445=>x"6c00", 446=>x"6d00", 447=>x"6d00", 448=>x"6600",
--449=>x"6400", 450=>x"6700", 451=>x"6b00", 452=>x"6d00", 453=>x"6a00", 454=>x"6e00", 455=>x"6f00",
--456=>x"6000", 457=>x"6500", 458=>x"6800", 459=>x"6d00", 460=>x"6c00", 461=>x"6b00", 462=>x"6b00",
--463=>x"6c00", 464=>x"6300", 465=>x"6300", 466=>x"6300", 467=>x"6700", 468=>x"6400", 469=>x"6900",
--470=>x"6b00", 471=>x"6e00", 472=>x"6100", 473=>x"6100", 474=>x"6300", 475=>x"6a00", 476=>x"6700",
--477=>x"6800", 478=>x"6900", 479=>x"6a00", 480=>x"6300", 481=>x"6300", 482=>x"6400", 483=>x"6600",
--484=>x"6800", 485=>x"9700", 486=>x"6b00", 487=>x"6b00", 488=>x"6300", 489=>x"6400", 490=>x"6300",
--491=>x"6600", 492=>x"6800", 493=>x"6800", 494=>x"6900", 495=>x"6900", 496=>x"6300", 497=>x"6500",
--498=>x"6300", 499=>x"6500"),
--7  => (0=>x"7400", 1=>x"8500", 2=>x"7c00", 3=>x"7900", 4=>x"7d00", 5=>x"8000", 6=>x"7a00", 7=>x"8300",
--8=>x"7500", 9=>x"7a00", 10=>x"7a00", 11=>x"7900", 12=>x"7f00", 13=>x"8000", 14=>x"7b00",
--15=>x"8300", 16=>x"7500", 17=>x"7900", 18=>x"7b00", 19=>x"7a00", 20=>x"7e00", 21=>x"8000",
--22=>x"7b00", 23=>x"8100", 24=>x"8900", 25=>x"7900", 26=>x"7d00", 27=>x"7c00", 28=>x"7d00",
--29=>x"7b00", 30=>x"7c00", 31=>x"7c00", 32=>x"7700", 33=>x"7a00", 34=>x"7a00", 35=>x"7c00",
--36=>x"7d00", 37=>x"7d00", 38=>x"7b00", 39=>x"7c00", 40=>x"7400", 41=>x"7900", 42=>x"7b00",
--43=>x"7c00", 44=>x"7b00", 45=>x"7c00", 46=>x"7d00", 47=>x"8000", 48=>x"7700", 49=>x"7500",
--50=>x"7a00", 51=>x"7a00", 52=>x"7a00", 53=>x"7d00", 54=>x"7f00", 55=>x"7d00", 56=>x"7600",
--57=>x"7600", 58=>x"7a00", 59=>x"7800", 60=>x"7d00", 61=>x"7c00", 62=>x"7d00", 63=>x"8000",
--64=>x"7300", 65=>x"7800", 66=>x"7a00", 67=>x"7d00", 68=>x"7c00", 69=>x"7e00", 70=>x"7f00",
--71=>x"8000", 72=>x"7700", 73=>x"7700", 74=>x"7800", 75=>x"7a00", 76=>x"7b00", 77=>x"7d00",
--78=>x"7a00", 79=>x"7f00", 80=>x"7700", 81=>x"7800", 82=>x"7800", 83=>x"7700", 84=>x"7c00",
--85=>x"7c00", 86=>x"7a00", 87=>x"7d00", 88=>x"7400", 89=>x"7600", 90=>x"7700", 91=>x"7900",
--92=>x"7b00", 93=>x"7d00", 94=>x"7d00", 95=>x"7b00", 96=>x"7500", 97=>x"7900", 98=>x"7a00",
--99=>x"7800", 100=>x"7800", 101=>x"7800", 102=>x"7f00", 103=>x"7f00", 104=>x"7700", 105=>x"7900",
--106=>x"7700", 107=>x"7a00", 108=>x"7a00", 109=>x"7c00", 110=>x"7b00", 111=>x"7d00", 112=>x"7500",
--113=>x"7a00", 114=>x"7800", 115=>x"7800", 116=>x"7c00", 117=>x"7d00", 118=>x"7c00", 119=>x"7f00",
--120=>x"7400", 121=>x"7600", 122=>x"7a00", 123=>x"7a00", 124=>x"7a00", 125=>x"7c00", 126=>x"7d00",
--127=>x"7b00", 128=>x"7500", 129=>x"7700", 130=>x"7a00", 131=>x"7900", 132=>x"7c00", 133=>x"7800",
--134=>x"7a00", 135=>x"8200", 136=>x"7400", 137=>x"7500", 138=>x"7800", 139=>x"7a00", 140=>x"7c00",
--141=>x"7c00", 142=>x"7b00", 143=>x"7e00", 144=>x"7700", 145=>x"7400", 146=>x"7800", 147=>x"7800",
--148=>x"7600", 149=>x"7800", 150=>x"7d00", 151=>x"7b00", 152=>x"7300", 153=>x"7300", 154=>x"7900",
--155=>x"7900", 156=>x"7600", 157=>x"7700", 158=>x"7a00", 159=>x"7c00", 160=>x"7400", 161=>x"7700",
--162=>x"7700", 163=>x"7900", 164=>x"7900", 165=>x"7a00", 166=>x"7700", 167=>x"7800", 168=>x"7500",
--169=>x"7a00", 170=>x"7800", 171=>x"7700", 172=>x"7600", 173=>x"8500", 174=>x"8300", 175=>x"7a00",
--176=>x"7500", 177=>x"7800", 178=>x"7800", 179=>x"7800", 180=>x"7700", 181=>x"7a00", 182=>x"7d00",
--183=>x"7b00", 184=>x"7500", 185=>x"7800", 186=>x"7800", 187=>x"7900", 188=>x"7a00", 189=>x"7c00",
--190=>x"7a00", 191=>x"7b00", 192=>x"7200", 193=>x"7700", 194=>x"7900", 195=>x"7a00", 196=>x"8700",
--197=>x"7c00", 198=>x"7c00", 199=>x"7c00", 200=>x"7400", 201=>x"7900", 202=>x"7900", 203=>x"7900",
--204=>x"7800", 205=>x"8500", 206=>x"7e00", 207=>x"7c00", 208=>x"7600", 209=>x"7800", 210=>x"7900",
--211=>x"7b00", 212=>x"7800", 213=>x"7800", 214=>x"7a00", 215=>x"7c00", 216=>x"7500", 217=>x"7a00",
--218=>x"7900", 219=>x"7a00", 220=>x"7c00", 221=>x"7a00", 222=>x"7b00", 223=>x"7e00", 224=>x"7600",
--225=>x"7800", 226=>x"7800", 227=>x"7700", 228=>x"7a00", 229=>x"7a00", 230=>x"7e00", 231=>x"7b00",
--232=>x"7400", 233=>x"7500", 234=>x"7600", 235=>x"7900", 236=>x"7a00", 237=>x"7900", 238=>x"7b00",
--239=>x"7a00", 240=>x"7500", 241=>x"7500", 242=>x"7500", 243=>x"7500", 244=>x"7800", 245=>x"7b00",
--246=>x"7900", 247=>x"7900", 248=>x"7500", 249=>x"7500", 250=>x"7500", 251=>x"7500", 252=>x"7700",
--253=>x"7a00", 254=>x"7900", 255=>x"7700", 256=>x"7300", 257=>x"7500", 258=>x"7500", 259=>x"7200",
--260=>x"7800", 261=>x"7700", 262=>x"7900", 263=>x"7600", 264=>x"7000", 265=>x"7400", 266=>x"7500",
--267=>x"7200", 268=>x"7700", 269=>x"7400", 270=>x"7300", 271=>x"7500", 272=>x"7000", 273=>x"7100",
--274=>x"7000", 275=>x"8e00", 276=>x"7200", 277=>x"8900", 278=>x"7500", 279=>x"7600", 280=>x"7200",
--281=>x"7600", 282=>x"6f00", 283=>x"7100", 284=>x"7400", 285=>x"7500", 286=>x"7600", 287=>x"7700",
--288=>x"7100", 289=>x"7200", 290=>x"7200", 291=>x"7400", 292=>x"7300", 293=>x"7500", 294=>x"7300",
--295=>x"7600", 296=>x"7100", 297=>x"6f00", 298=>x"7300", 299=>x"8b00", 300=>x"7100", 301=>x"7200",
--302=>x"7400", 303=>x"7600", 304=>x"6d00", 305=>x"7100", 306=>x"7200", 307=>x"7600", 308=>x"8d00",
--309=>x"7300", 310=>x"7500", 311=>x"7a00", 312=>x"7200", 313=>x"7500", 314=>x"7400", 315=>x"7300",
--316=>x"7200", 317=>x"7100", 318=>x"7200", 319=>x"7400", 320=>x"7000", 321=>x"7200", 322=>x"7700",
--323=>x"7100", 324=>x"7400", 325=>x"7400", 326=>x"7800", 327=>x"7700", 328=>x"6e00", 329=>x"7000",
--330=>x"7200", 331=>x"7200", 332=>x"7100", 333=>x"7400", 334=>x"7500", 335=>x"7900", 336=>x"7100",
--337=>x"7500", 338=>x"7100", 339=>x"7300", 340=>x"7500", 341=>x"7500", 342=>x"7600", 343=>x"7600",
--344=>x"7000", 345=>x"7200", 346=>x"7200", 347=>x"7200", 348=>x"7400", 349=>x"7500", 350=>x"7500",
--351=>x"7600", 352=>x"6d00", 353=>x"7200", 354=>x"7300", 355=>x"7400", 356=>x"7500", 357=>x"7300",
--358=>x"7600", 359=>x"7800", 360=>x"6f00", 361=>x"7200", 362=>x"7400", 363=>x"7300", 364=>x"7400",
--365=>x"7500", 366=>x"7800", 367=>x"7b00", 368=>x"7000", 369=>x"7000", 370=>x"7400", 371=>x"7600",
--372=>x"7400", 373=>x"7600", 374=>x"7800", 375=>x"7800", 376=>x"7400", 377=>x"7200", 378=>x"7300",
--379=>x"7400", 380=>x"7400", 381=>x"7600", 382=>x"7700", 383=>x"7600", 384=>x"7000", 385=>x"7000",
--386=>x"7700", 387=>x"7800", 388=>x"7300", 389=>x"7400", 390=>x"7500", 391=>x"7500", 392=>x"7000",
--393=>x"7300", 394=>x"7900", 395=>x"7500", 396=>x"7400", 397=>x"7200", 398=>x"7600", 399=>x"7800",
--400=>x"6d00", 401=>x"7100", 402=>x"7400", 403=>x"7200", 404=>x"7200", 405=>x"7700", 406=>x"7700",
--407=>x"7500", 408=>x"7000", 409=>x"7400", 410=>x"7400", 411=>x"7600", 412=>x"7600", 413=>x"7600",
--414=>x"7600", 415=>x"7600", 416=>x"6e00", 417=>x"7100", 418=>x"7400", 419=>x"7500", 420=>x"7700",
--421=>x"7a00", 422=>x"7800", 423=>x"7300", 424=>x"7100", 425=>x"7000", 426=>x"7100", 427=>x"7500",
--428=>x"7600", 429=>x"7400", 430=>x"7500", 431=>x"7200", 432=>x"7300", 433=>x"7300", 434=>x"7600",
--435=>x"7300", 436=>x"7000", 437=>x"7300", 438=>x"7200", 439=>x"7100", 440=>x"7100", 441=>x"7200",
--442=>x"7000", 443=>x"7300", 444=>x"7500", 445=>x"7400", 446=>x"6e00", 447=>x"6b00", 448=>x"6d00",
--449=>x"7200", 450=>x"7300", 451=>x"7200", 452=>x"6f00", 453=>x"6e00", 454=>x"6d00", 455=>x"6700",
--456=>x"6e00", 457=>x"7000", 458=>x"7200", 459=>x"8d00", 460=>x"6f00", 461=>x"6f00", 462=>x"6b00",
--463=>x"6b00", 464=>x"6d00", 465=>x"7100", 466=>x"6f00", 467=>x"6f00", 468=>x"6c00", 469=>x"6b00",
--470=>x"6100", 471=>x"8300", 472=>x"6a00", 473=>x"6d00", 474=>x"6e00", 475=>x"6e00", 476=>x"6b00",
--477=>x"6500", 478=>x"6100", 479=>x"a700", 480=>x"6c00", 481=>x"6f00", 482=>x"7000", 483=>x"6c00",
--484=>x"6e00", 485=>x"6500", 486=>x"6f00", 487=>x"c700", 488=>x"6d00", 489=>x"7200", 490=>x"7000",
--491=>x"6e00", 492=>x"6c00", 493=>x"6200", 494=>x"8000", 495=>x"d100", 496=>x"6c00", 497=>x"7100",
--498=>x"7200", 499=>x"7500"),
--8  => (0=>x"7c00", 1=>x"8300", 2=>x"8000", 3=>x"8100", 4=>x"8500", 5=>x"8600", 6=>x"8300", 7=>x"8000",
--8=>x"8300", 9=>x"8300", 10=>x"8100", 11=>x"8100", 12=>x"8500", 13=>x"8600", 14=>x"8400",
--15=>x"8100", 16=>x"8200", 17=>x"8300", 18=>x"8200", 19=>x"8100", 20=>x"8400", 21=>x"8500",
--22=>x"8400", 23=>x"8200", 24=>x"7c00", 25=>x"8100", 26=>x"8400", 27=>x"8000", 28=>x"8100",
--29=>x"8200", 30=>x"8400", 31=>x"8100", 32=>x"7e00", 33=>x"8000", 34=>x"8000", 35=>x"8200",
--36=>x"8300", 37=>x"8200", 38=>x"8200", 39=>x"8200", 40=>x"7f00", 41=>x"8300", 42=>x"7f00",
--43=>x"8000", 44=>x"8100", 45=>x"8100", 46=>x"8000", 47=>x"8300", 48=>x"7e00", 49=>x"7e00",
--50=>x"7f00", 51=>x"8300", 52=>x"7e00", 53=>x"8200", 54=>x"8100", 55=>x"8400", 56=>x"7e00",
--57=>x"7d00", 58=>x"8000", 59=>x"8000", 60=>x"7d00", 61=>x"8300", 62=>x"8300", 63=>x"8300",
--64=>x"7f00", 65=>x"8100", 66=>x"7f00", 67=>x"8300", 68=>x"7f00", 69=>x"8200", 70=>x"8200",
--71=>x"8200", 72=>x"8000", 73=>x"8000", 74=>x"8000", 75=>x"8200", 76=>x"8100", 77=>x"8100",
--78=>x"8500", 79=>x"8400", 80=>x"7d00", 81=>x"7f00", 82=>x"8000", 83=>x"8100", 84=>x"8100",
--85=>x"8100", 86=>x"8300", 87=>x"8100", 88=>x"7c00", 89=>x"8000", 90=>x"8000", 91=>x"8200",
--92=>x"8200", 93=>x"8000", 94=>x"8300", 95=>x"8100", 96=>x"8000", 97=>x"8300", 98=>x"7f00",
--99=>x"7e00", 100=>x"8000", 101=>x"8300", 102=>x"8100", 103=>x"8200", 104=>x"7f00", 105=>x"8100",
--106=>x"8000", 107=>x"7d00", 108=>x"7f00", 109=>x"8100", 110=>x"8100", 111=>x"8200", 112=>x"8000",
--113=>x"7e00", 114=>x"7d00", 115=>x"7e00", 116=>x"8100", 117=>x"7e00", 118=>x"7e00", 119=>x"8100",
--120=>x"7e00", 121=>x"7e00", 122=>x"8000", 123=>x"7f00", 124=>x"7f00", 125=>x"8000", 126=>x"7f00",
--127=>x"7e00", 128=>x"7e00", 129=>x"7e00", 130=>x"8100", 131=>x"7d00", 132=>x"7e00", 133=>x"8100",
--134=>x"8000", 135=>x"7f00", 136=>x"7d00", 137=>x"7d00", 138=>x"7f00", 139=>x"8100", 140=>x"8000",
--141=>x"7f00", 142=>x"8000", 143=>x"8200", 144=>x"7a00", 145=>x"7c00", 146=>x"7f00", 147=>x"8000",
--148=>x"7f00", 149=>x"7d00", 150=>x"8200", 151=>x"8100", 152=>x"7c00", 153=>x"7d00", 154=>x"7e00",
--155=>x"7e00", 156=>x"7b00", 157=>x"7b00", 158=>x"8100", 159=>x"8100", 160=>x"7c00", 161=>x"7a00",
--162=>x"7900", 163=>x"7e00", 164=>x"7e00", 165=>x"7d00", 166=>x"7d00", 167=>x"7e00", 168=>x"7c00",
--169=>x"7d00", 170=>x"7800", 171=>x"7c00", 172=>x"7c00", 173=>x"8000", 174=>x"7e00", 175=>x"7a00",
--176=>x"7d00", 177=>x"7d00", 178=>x"7c00", 179=>x"7b00", 180=>x"8200", 181=>x"7e00", 182=>x"7d00",
--183=>x"7c00", 184=>x"7b00", 185=>x"7c00", 186=>x"7b00", 187=>x"7e00", 188=>x"7e00", 189=>x"7f00",
--190=>x"7d00", 191=>x"7b00", 192=>x"7b00", 193=>x"7d00", 194=>x"7c00", 195=>x"7f00", 196=>x"7f00",
--197=>x"7f00", 198=>x"8000", 199=>x"7f00", 200=>x"7f00", 201=>x"7c00", 202=>x"8400", 203=>x"7e00",
--204=>x"7d00", 205=>x"7e00", 206=>x"7d00", 207=>x"7f00", 208=>x"7f00", 209=>x"8000", 210=>x"7d00",
--211=>x"7d00", 212=>x"7b00", 213=>x"7d00", 214=>x"7d00", 215=>x"7d00", 216=>x"8200", 217=>x"7e00",
--218=>x"7f00", 219=>x"7c00", 220=>x"7c00", 221=>x"7c00", 222=>x"8000", 223=>x"8100", 224=>x"7f00",
--225=>x"7c00", 226=>x"7c00", 227=>x"7d00", 228=>x"7e00", 229=>x"7d00", 230=>x"8000", 231=>x"8000",
--232=>x"7c00", 233=>x"7900", 234=>x"7a00", 235=>x"7b00", 236=>x"7700", 237=>x"7e00", 238=>x"7e00",
--239=>x"7b00", 240=>x"7800", 241=>x"7a00", 242=>x"7d00", 243=>x"7a00", 244=>x"7b00", 245=>x"7900",
--246=>x"7e00", 247=>x"7e00", 248=>x"7a00", 249=>x"7a00", 250=>x"7d00", 251=>x"7b00", 252=>x"8300",
--253=>x"7c00", 254=>x"7c00", 255=>x"7d00", 256=>x"7b00", 257=>x"7900", 258=>x"7b00", 259=>x"7b00",
--260=>x"7800", 261=>x"7a00", 262=>x"7c00", 263=>x"7e00", 264=>x"7c00", 265=>x"7c00", 266=>x"7a00",
--267=>x"7c00", 268=>x"7b00", 269=>x"7b00", 270=>x"7c00", 271=>x"7c00", 272=>x"7900", 273=>x"7c00",
--274=>x"7800", 275=>x"7900", 276=>x"7a00", 277=>x"7d00", 278=>x"7a00", 279=>x"7b00", 280=>x"7600",
--281=>x"7700", 282=>x"7700", 283=>x"7700", 284=>x"7b00", 285=>x"7b00", 286=>x"7a00", 287=>x"7e00",
--288=>x"7700", 289=>x"7700", 290=>x"7500", 291=>x"7800", 292=>x"7900", 293=>x"7600", 294=>x"7b00",
--295=>x"7b00", 296=>x"7900", 297=>x"7900", 298=>x"7700", 299=>x"7700", 300=>x"7900", 301=>x"8500",
--302=>x"7a00", 303=>x"7c00", 304=>x"8800", 305=>x"7500", 306=>x"7700", 307=>x"7600", 308=>x"7800",
--309=>x"7b00", 310=>x"7800", 311=>x"7900", 312=>x"7800", 313=>x"7900", 314=>x"7800", 315=>x"7800",
--316=>x"7c00", 317=>x"7a00", 318=>x"7900", 319=>x"7900", 320=>x"7b00", 321=>x"7900", 322=>x"7d00",
--323=>x"7900", 324=>x"7b00", 325=>x"7d00", 326=>x"7600", 327=>x"7700", 328=>x"7900", 329=>x"7600",
--330=>x"7a00", 331=>x"7a00", 332=>x"7a00", 333=>x"7700", 334=>x"7900", 335=>x"7b00", 336=>x"7900",
--337=>x"7900", 338=>x"7900", 339=>x"7800", 340=>x"7c00", 341=>x"7900", 342=>x"7d00", 343=>x"7b00",
--344=>x"7800", 345=>x"7800", 346=>x"7800", 347=>x"7800", 348=>x"7b00", 349=>x"7a00", 350=>x"7e00",
--351=>x"7b00", 352=>x"7900", 353=>x"7700", 354=>x"7900", 355=>x"7900", 356=>x"7a00", 357=>x"7b00",
--358=>x"7b00", 359=>x"8100", 360=>x"7a00", 361=>x"7a00", 362=>x"7800", 363=>x"7c00", 364=>x"7800",
--365=>x"7700", 366=>x"8100", 367=>x"8100", 368=>x"7900", 369=>x"7c00", 370=>x"7800", 371=>x"7800",
--372=>x"8400", 373=>x"7b00", 374=>x"7f00", 375=>x"7200", 376=>x"7600", 377=>x"7800", 378=>x"7b00",
--379=>x"7c00", 380=>x"7b00", 381=>x"7f00", 382=>x"7900", 383=>x"7000", 384=>x"7700", 385=>x"7700",
--386=>x"7800", 387=>x"7a00", 388=>x"7f00", 389=>x"7e00", 390=>x"7400", 391=>x"7500", 392=>x"8500",
--393=>x"7900", 394=>x"7800", 395=>x"7a00", 396=>x"8900", 397=>x"7800", 398=>x"6f00", 399=>x"7100",
--400=>x"7b00", 401=>x"7700", 402=>x"7800", 403=>x"8500", 404=>x"8900", 405=>x"6f00", 406=>x"6b00",
--407=>x"6c00", 408=>x"7900", 409=>x"7600", 410=>x"7a00", 411=>x"8900", 412=>x"7b00", 413=>x"6d00",
--414=>x"6e00", 415=>x"6900", 416=>x"7300", 417=>x"7400", 418=>x"9400", 419=>x"8500", 420=>x"6d00",
--421=>x"6900", 422=>x"6700", 423=>x"6500", 424=>x"6f00", 425=>x"8700", 426=>x"b600", 427=>x"7b00",
--428=>x"6400", 429=>x"6500", 430=>x"6800", 431=>x"6700", 432=>x"6c00", 433=>x"9f00", 434=>x"b300",
--435=>x"7400", 436=>x"5f00", 437=>x"6700", 438=>x"6b00", 439=>x"6c00", 440=>x"7400", 441=>x"c000",
--442=>x"a900", 443=>x"6900", 444=>x"6200", 445=>x"6700", 446=>x"6d00", 447=>x"6900", 448=>x"9800",
--449=>x"cf00", 450=>x"9400", 451=>x"6400", 452=>x"6600", 453=>x"6900", 454=>x"6700", 455=>x"6900",
--456=>x"be00", 457=>x"c700", 458=>x"8a00", 459=>x"6100", 460=>x"6600", 461=>x"6b00", 462=>x"6700",
--463=>x"6700", 464=>x"d600", 465=>x"b600", 466=>x"7a00", 467=>x"6000", 468=>x"6700", 469=>x"6800",
--470=>x"6600", 471=>x"6a00", 472=>x"d900", 473=>x"a000", 474=>x"7b00", 475=>x"6600", 476=>x"6300",
--477=>x"6700", 478=>x"6700", 479=>x"6a00", 480=>x"c800", 481=>x"a700", 482=>x"8400", 483=>x"6700",
--484=>x"6100", 485=>x"6800", 486=>x"6800", 487=>x"6a00", 488=>x"c300", 489=>x"a200", 490=>x"7a00",
--491=>x"6600", 492=>x"9a00", 493=>x"6200", 494=>x"6400", 495=>x"6a00", 496=>x"be00", 497=>x"9600",
--498=>x"7300", 499=>x"6000"),
--9  => (0=>x"8300", 1=>x"7f00", 2=>x"8400", 3=>x"8200", 4=>x"8300", 5=>x"8100", 6=>x"8500", 7=>x"8700",
--8=>x"8200", 9=>x"7f00", 10=>x"8300", 11=>x"8200", 12=>x"8200", 13=>x"8000", 14=>x"8600",
--15=>x"8700", 16=>x"8300", 17=>x"7e00", 18=>x"8300", 19=>x"8200", 20=>x"8100", 21=>x"8100",
--22=>x"8600", 23=>x"8700", 24=>x"8100", 25=>x"8300", 26=>x"7b00", 27=>x"8200", 28=>x"8000",
--29=>x"8400", 30=>x"8300", 31=>x"8300", 32=>x"8300", 33=>x"8200", 34=>x"8300", 35=>x"8200",
--36=>x"8200", 37=>x"8200", 38=>x"8200", 39=>x"8300", 40=>x"8300", 41=>x"8300", 42=>x"8300",
--43=>x"8000", 44=>x"8200", 45=>x"8200", 46=>x"8000", 47=>x"8300", 48=>x"8400", 49=>x"8400",
--50=>x"8200", 51=>x"8100", 52=>x"8300", 53=>x"7d00", 54=>x"8100", 55=>x"8600", 56=>x"8200",
--57=>x"7c00", 58=>x"8200", 59=>x"8100", 60=>x"8200", 61=>x"8100", 62=>x"8300", 63=>x"8300",
--64=>x"8300", 65=>x"8300", 66=>x"8200", 67=>x"8300", 68=>x"8300", 69=>x"8300", 70=>x"8000",
--71=>x"8200", 72=>x"8100", 73=>x"8300", 74=>x"8500", 75=>x"8400", 76=>x"8500", 77=>x"8300",
--78=>x"8100", 79=>x"8200", 80=>x"8000", 81=>x"8500", 82=>x"8200", 83=>x"8300", 84=>x"8400",
--85=>x"8300", 86=>x"8200", 87=>x"8300", 88=>x"8100", 89=>x"8200", 90=>x"8200", 91=>x"8000",
--92=>x"8100", 93=>x"8000", 94=>x"8200", 95=>x"8200", 96=>x"8200", 97=>x"8100", 98=>x"8200",
--99=>x"8400", 100=>x"8000", 101=>x"8000", 102=>x"8100", 103=>x"8100", 104=>x"8000", 105=>x"8000",
--106=>x"7f00", 107=>x"8100", 108=>x"8000", 109=>x"8200", 110=>x"8400", 111=>x"8000", 112=>x"7f00",
--113=>x"7f00", 114=>x"8200", 115=>x"8000", 116=>x"8300", 117=>x"8200", 118=>x"8100", 119=>x"8300",
--120=>x"7f00", 121=>x"7d00", 122=>x"8000", 123=>x"8000", 124=>x"8000", 125=>x"8200", 126=>x"8100",
--127=>x"8000", 128=>x"7e00", 129=>x"7c00", 130=>x"7f00", 131=>x"8100", 132=>x"7f00", 133=>x"8300",
--134=>x"8100", 135=>x"8100", 136=>x"7f00", 137=>x"8100", 138=>x"7f00", 139=>x"7f00", 140=>x"7e00",
--141=>x"7f00", 142=>x"8100", 143=>x"8300", 144=>x"7f00", 145=>x"8000", 146=>x"7c00", 147=>x"7e00",
--148=>x"7b00", 149=>x"7d00", 150=>x"8100", 151=>x"8100", 152=>x"7d00", 153=>x"7d00", 154=>x"7a00",
--155=>x"7e00", 156=>x"7e00", 157=>x"7f00", 158=>x"7f00", 159=>x"8000", 160=>x"8000", 161=>x"7c00",
--162=>x"7b00", 163=>x"7c00", 164=>x"7d00", 165=>x"7d00", 166=>x"8100", 167=>x"7f00", 168=>x"7c00",
--169=>x"7d00", 170=>x"7e00", 171=>x"7e00", 172=>x"7f00", 173=>x"7f00", 174=>x"8100", 175=>x"7f00",
--176=>x"7c00", 177=>x"7d00", 178=>x"7d00", 179=>x"8000", 180=>x"8000", 181=>x"8200", 182=>x"8300",
--183=>x"8000", 184=>x"7e00", 185=>x"8000", 186=>x"7f00", 187=>x"8300", 188=>x"8000", 189=>x"7f00",
--190=>x"8300", 191=>x"8100", 192=>x"7d00", 193=>x"7e00", 194=>x"7f00", 195=>x"8100", 196=>x"7f00",
--197=>x"8200", 198=>x"8000", 199=>x"7e00", 200=>x"7e00", 201=>x"8100", 202=>x"8200", 203=>x"8000",
--204=>x"8100", 205=>x"8200", 206=>x"8200", 207=>x"7c00", 208=>x"7e00", 209=>x"8400", 210=>x"8100",
--211=>x"8000", 212=>x"8000", 213=>x"8100", 214=>x"8100", 215=>x"7d00", 216=>x"8300", 217=>x"8200",
--218=>x"7e00", 219=>x"7e00", 220=>x"7e00", 221=>x"8000", 222=>x"8300", 223=>x"8100", 224=>x"7f00",
--225=>x"7d00", 226=>x"8100", 227=>x"7e00", 228=>x"8000", 229=>x"8100", 230=>x"8000", 231=>x"8000",
--232=>x"7d00", 233=>x"7f00", 234=>x"7d00", 235=>x"7e00", 236=>x"7f00", 237=>x"8000", 238=>x"8000",
--239=>x"8000", 240=>x"7c00", 241=>x"8000", 242=>x"7e00", 243=>x"8000", 244=>x"7f00", 245=>x"7f00",
--246=>x"7b00", 247=>x"7b00", 248=>x"7f00", 249=>x"7e00", 250=>x"7e00", 251=>x"7d00", 252=>x"7d00",
--253=>x"7f00", 254=>x"7800", 255=>x"8500", 256=>x"7d00", 257=>x"7a00", 258=>x"7d00", 259=>x"7c00",
--260=>x"7b00", 261=>x"7b00", 262=>x"7b00", 263=>x"a900", 264=>x"7d00", 265=>x"8300", 266=>x"7d00",
--267=>x"7a00", 268=>x"7900", 269=>x"7600", 270=>x"9b00", 271=>x"a800", 272=>x"7c00", 273=>x"7c00",
--274=>x"7c00", 275=>x"7c00", 276=>x"7d00", 277=>x"7500", 278=>x"6400", 279=>x"8e00", 280=>x"7f00",
--281=>x"7a00", 282=>x"7e00", 283=>x"7f00", 284=>x"7d00", 285=>x"8600", 286=>x"7400", 287=>x"6a00",
--288=>x"7d00", 289=>x"7900", 290=>x"7a00", 291=>x"7700", 292=>x"8100", 293=>x"9100", 294=>x"7000",
--295=>x"6f00", 296=>x"7c00", 297=>x"7b00", 298=>x"7a00", 299=>x"7900", 300=>x"ac00", 301=>x"8900",
--302=>x"6a00", 303=>x"7300", 304=>x"7d00", 305=>x"7d00", 306=>x"7600", 307=>x"8a00", 308=>x"a500",
--309=>x"7400", 310=>x"7200", 311=>x"7300", 312=>x"7c00", 313=>x"7c00", 314=>x"7900", 315=>x"9500",
--316=>x"8400", 317=>x"7000", 318=>x"7300", 319=>x"6b00", 320=>x"7c00", 321=>x"7e00", 322=>x"8300",
--323=>x"8500", 324=>x"7700", 325=>x"7000", 326=>x"6c00", 327=>x"6d00", 328=>x"7c00", 329=>x"7d00",
--330=>x"8200", 331=>x"7b00", 332=>x"6d00", 333=>x"6d00", 334=>x"6c00", 335=>x"6e00", 336=>x"7c00",
--337=>x"8400", 338=>x"7c00", 339=>x"6d00", 340=>x"6d00", 341=>x"6a00", 342=>x"6f00", 343=>x"6d00",
--344=>x"7e00", 345=>x"8000", 346=>x"7000", 347=>x"6800", 348=>x"6a00", 349=>x"6c00", 350=>x"6f00",
--351=>x"7000", 352=>x"7c00", 353=>x"7200", 354=>x"6e00", 355=>x"6c00", 356=>x"6a00", 357=>x"6b00",
--358=>x"6f00", 359=>x"7300", 360=>x"7000", 361=>x"6c00", 362=>x"6a00", 363=>x"6b00", 364=>x"6d00",
--365=>x"6d00", 366=>x"6f00", 367=>x"7300", 368=>x"6a00", 369=>x"6e00", 370=>x"6b00", 371=>x"6e00",
--372=>x"7300", 373=>x"7100", 374=>x"7100", 375=>x"6f00", 376=>x"6d00", 377=>x"6900", 378=>x"6f00",
--379=>x"7500", 380=>x"6f00", 381=>x"6f00", 382=>x"7400", 383=>x"7000", 384=>x"6f00", 385=>x"7000",
--386=>x"6e00", 387=>x"7100", 388=>x"7200", 389=>x"7000", 390=>x"7000", 391=>x"7400", 392=>x"7200",
--393=>x"7500", 394=>x"6e00", 395=>x"9200", 396=>x"6e00", 397=>x"7000", 398=>x"7100", 399=>x"7400",
--400=>x"6d00", 401=>x"7400", 402=>x"7400", 403=>x"6d00", 404=>x"6d00", 405=>x"6e00", 406=>x"7100",
--407=>x"7100", 408=>x"6b00", 409=>x"7100", 410=>x"7400", 411=>x"7100", 412=>x"7200", 413=>x"7000",
--414=>x"7000", 415=>x"6f00", 416=>x"6700", 417=>x"6c00", 418=>x"7600", 419=>x"7400", 420=>x"7300",
--421=>x"7100", 422=>x"7100", 423=>x"7500", 424=>x"6900", 425=>x"6c00", 426=>x"7000", 427=>x"7100",
--428=>x"7300", 429=>x"7000", 430=>x"6e00", 431=>x"6f00", 432=>x"6800", 433=>x"7200", 434=>x"6f00",
--435=>x"7000", 436=>x"6f00", 437=>x"7100", 438=>x"7100", 439=>x"7200", 440=>x"6c00", 441=>x"6d00",
--442=>x"6d00", 443=>x"7100", 444=>x"6c00", 445=>x"7000", 446=>x"7300", 447=>x"7100", 448=>x"6c00",
--449=>x"6d00", 450=>x"6b00", 451=>x"6f00", 452=>x"6e00", 453=>x"8e00", 454=>x"7200", 455=>x"7200",
--456=>x"6900", 457=>x"7000", 458=>x"6f00", 459=>x"6d00", 460=>x"7300", 461=>x"7100", 462=>x"6c00",
--463=>x"6b00", 464=>x"6b00", 465=>x"6c00", 466=>x"7400", 467=>x"7700", 468=>x"6f00", 469=>x"6e00",
--470=>x"7400", 471=>x"6c00", 472=>x"6e00", 473=>x"6d00", 474=>x"7000", 475=>x"7400", 476=>x"7000",
--477=>x"7100", 478=>x"7500", 479=>x"7500", 480=>x"7000", 481=>x"6c00", 482=>x"6900", 483=>x"7400",
--484=>x"7300", 485=>x"7400", 486=>x"7300", 487=>x"7800", 488=>x"6e00", 489=>x"6700", 490=>x"6f00",
--491=>x"7b00", 492=>x"6e00", 493=>x"7000", 494=>x"7400", 495=>x"7300", 496=>x"6900", 497=>x"6d00",
--498=>x"7200", 499=>x"8600"),
--10 => (0=>x"8100", 1=>x"8600", 2=>x"8500", 3=>x"8600", 4=>x"8600", 5=>x"8500", 6=>x"8600", 7=>x"8600",
--8=>x"8200", 9=>x"8400", 10=>x"8500", 11=>x"8600", 12=>x"8500", 13=>x"8600", 14=>x"8600",
--15=>x"8400", 16=>x"8300", 17=>x"7900", 18=>x"8600", 19=>x"8700", 20=>x"8600", 21=>x"8400",
--22=>x"8600", 23=>x"8500", 24=>x"8300", 25=>x"8500", 26=>x"8700", 27=>x"8700", 28=>x"8500",
--29=>x"8400", 30=>x"8500", 31=>x"7800", 32=>x"8400", 33=>x"8300", 34=>x"8300", 35=>x"8500",
--36=>x"8500", 37=>x"8500", 38=>x"8600", 39=>x"8500", 40=>x"8200", 41=>x"8300", 42=>x"7b00",
--43=>x"8600", 44=>x"8400", 45=>x"8400", 46=>x"8500", 47=>x"8500", 48=>x"8000", 49=>x"8300",
--50=>x"8500", 51=>x"8400", 52=>x"8400", 53=>x"8300", 54=>x"8400", 55=>x"8400", 56=>x"8100",
--57=>x"8300", 58=>x"8000", 59=>x"8200", 60=>x"8100", 61=>x"8500", 62=>x"8600", 63=>x"8500",
--64=>x"8400", 65=>x"8600", 66=>x"8700", 67=>x"8400", 68=>x"8300", 69=>x"8700", 70=>x"8400",
--71=>x"8600", 72=>x"8300", 73=>x"8300", 74=>x"8600", 75=>x"8200", 76=>x"8300", 77=>x"8400",
--78=>x"8600", 79=>x"8500", 80=>x"8200", 81=>x"8000", 82=>x"8300", 83=>x"8300", 84=>x"8300",
--85=>x"8100", 86=>x"8400", 87=>x"8400", 88=>x"8100", 89=>x"8300", 90=>x"8400", 91=>x"8400",
--92=>x"8100", 93=>x"8300", 94=>x"8300", 95=>x"8400", 96=>x"8100", 97=>x"8100", 98=>x"8300",
--99=>x"8200", 100=>x"8000", 101=>x"8300", 102=>x"8600", 103=>x"8500", 104=>x"8100", 105=>x"8300",
--106=>x"8100", 107=>x"8000", 108=>x"7e00", 109=>x"8100", 110=>x"8000", 111=>x"8200", 112=>x"8200",
--113=>x"8200", 114=>x"8100", 115=>x"8400", 116=>x"8100", 117=>x"8100", 118=>x"8000", 119=>x"8400",
--120=>x"8000", 121=>x"8300", 122=>x"8200", 123=>x"8100", 124=>x"8200", 125=>x"8200", 126=>x"8000",
--127=>x"8300", 128=>x"8400", 129=>x"8200", 130=>x"8300", 131=>x"8300", 132=>x"8300", 133=>x"7d00",
--134=>x"8300", 135=>x"8200", 136=>x"8400", 137=>x"8200", 138=>x"8100", 139=>x"7f00", 140=>x"8100",
--141=>x"8300", 142=>x"8400", 143=>x"7f00", 144=>x"8000", 145=>x"7d00", 146=>x"8100", 147=>x"7f00",
--148=>x"8000", 149=>x"7f00", 150=>x"7e00", 151=>x"8000", 152=>x"8200", 153=>x"7f00", 154=>x"8200",
--155=>x"7f00", 156=>x"7c00", 157=>x"7d00", 158=>x"8000", 159=>x"8000", 160=>x"8300", 161=>x"8100",
--162=>x"8100", 163=>x"8000", 164=>x"7e00", 165=>x"8100", 166=>x"8200", 167=>x"8000", 168=>x"8000",
--169=>x"7d00", 170=>x"7f00", 171=>x"8000", 172=>x"7c00", 173=>x"8100", 174=>x"8000", 175=>x"7f00",
--176=>x"8000", 177=>x"7f00", 178=>x"7d00", 179=>x"7a00", 180=>x"7e00", 181=>x"8100", 182=>x"8100",
--183=>x"8000", 184=>x"8200", 185=>x"8000", 186=>x"7d00", 187=>x"7d00", 188=>x"7f00", 189=>x"8900",
--190=>x"8500", 191=>x"8000", 192=>x"8100", 193=>x"7f00", 194=>x"7e00", 195=>x"8000", 196=>x"7f00",
--197=>x"7f00", 198=>x"8000", 199=>x"8200", 200=>x"8200", 201=>x"7f00", 202=>x"7f00", 203=>x"7f00",
--204=>x"7f00", 205=>x"7f00", 206=>x"8100", 207=>x"8200", 208=>x"8200", 209=>x"8300", 210=>x"8000",
--211=>x"7f00", 212=>x"8000", 213=>x"8100", 214=>x"7f00", 215=>x"8000", 216=>x"8000", 217=>x"7e00",
--218=>x"7f00", 219=>x"7c00", 220=>x"7e00", 221=>x"7f00", 222=>x"7f00", 223=>x"7f00", 224=>x"8000",
--225=>x"7e00", 226=>x"7c00", 227=>x"7d00", 228=>x"7c00", 229=>x"7d00", 230=>x"8000", 231=>x"8200",
--232=>x"7d00", 233=>x"7a00", 234=>x"7b00", 235=>x"7a00", 236=>x"7e00", 237=>x"9100", 238=>x"9100",
--239=>x"9400", 240=>x"7900", 241=>x"7d00", 242=>x"a300", 243=>x"9900", 244=>x"9300", 245=>x"9f00",
--246=>x"9400", 247=>x"8e00", 248=>x"8600", 249=>x"8000", 250=>x"8d00", 251=>x"8d00", 252=>x"8d00",
--253=>x"8500", 254=>x"8200", 255=>x"7b00", 256=>x"9000", 257=>x"6f00", 258=>x"7b00", 259=>x"7b00",
--260=>x"7e00", 261=>x"7c00", 262=>x"7900", 263=>x"7700", 264=>x"5b00", 265=>x"6700", 266=>x"7b00",
--267=>x"7900", 268=>x"7800", 269=>x"7700", 270=>x"7b00", 271=>x"7600", 272=>x"6000", 273=>x"6e00",
--274=>x"7600", 275=>x"7600", 276=>x"7d00", 277=>x"7700", 278=>x"7900", 279=>x"7900", 280=>x"7300",
--281=>x"7000", 282=>x"7400", 283=>x"7700", 284=>x"7a00", 285=>x"7500", 286=>x"7700", 287=>x"7b00",
--288=>x"7200", 289=>x"7500", 290=>x"7600", 291=>x"7400", 292=>x"6e00", 293=>x"7000", 294=>x"7900",
--295=>x"7600", 296=>x"7500", 297=>x"7000", 298=>x"6f00", 299=>x"6d00", 300=>x"6e00", 301=>x"7200",
--302=>x"7400", 303=>x"7600", 304=>x"6c00", 305=>x"6e00", 306=>x"6900", 307=>x"6c00", 308=>x"7100",
--309=>x"7700", 310=>x"7800", 311=>x"7600", 312=>x"6a00", 313=>x"9400", 314=>x"6c00", 315=>x"7000",
--316=>x"7600", 317=>x"7800", 318=>x"7400", 319=>x"7400", 320=>x"6a00", 321=>x"6d00", 322=>x"6f00",
--323=>x"7100", 324=>x"7900", 325=>x"7500", 326=>x"7200", 327=>x"7400", 328=>x"7100", 329=>x"7100",
--330=>x"7500", 331=>x"7700", 332=>x"7a00", 333=>x"7500", 334=>x"7200", 335=>x"7c00", 336=>x"6f00",
--337=>x"8900", 338=>x"7800", 339=>x"7600", 340=>x"7400", 341=>x"7600", 342=>x"7d00", 343=>x"7800",
--344=>x"7300", 345=>x"7700", 346=>x"7200", 347=>x"7400", 348=>x"7a00", 349=>x"7b00", 350=>x"7a00",
--351=>x"7700", 352=>x"7300", 353=>x"7100", 354=>x"6f00", 355=>x"7a00", 356=>x"7b00", 357=>x"7500",
--358=>x"7200", 359=>x"7b00", 360=>x"6f00", 361=>x"7300", 362=>x"7d00", 363=>x"7500", 364=>x"7500",
--365=>x"7200", 366=>x"7200", 367=>x"7a00", 368=>x"7200", 369=>x"7900", 370=>x"7800", 371=>x"7600",
--372=>x"7700", 373=>x"7600", 374=>x"7600", 375=>x"7500", 376=>x"7700", 377=>x"7500", 378=>x"7300",
--379=>x"8700", 380=>x"7100", 381=>x"6f00", 382=>x"6e00", 383=>x"6a00", 384=>x"7800", 385=>x"7500",
--386=>x"7700", 387=>x"7000", 388=>x"6e00", 389=>x"7100", 390=>x"6e00", 391=>x"7300", 392=>x"7400",
--393=>x"7600", 394=>x"6f00", 395=>x"7400", 396=>x"7500", 397=>x"7900", 398=>x"7800", 399=>x"7b00",
--400=>x"7600", 401=>x"7700", 402=>x"7100", 403=>x"7800", 404=>x"7900", 405=>x"7a00", 406=>x"7600",
--407=>x"7600", 408=>x"7100", 409=>x"7000", 410=>x"7200", 411=>x"7400", 412=>x"7100", 413=>x"7600",
--414=>x"7700", 415=>x"7700", 416=>x"7400", 417=>x"7200", 418=>x"8d00", 419=>x"7100", 420=>x"7500",
--421=>x"7500", 422=>x"7400", 423=>x"7b00", 424=>x"7200", 425=>x"7200", 426=>x"6f00", 427=>x"6f00",
--428=>x"7300", 429=>x"8500", 430=>x"7b00", 431=>x"7b00", 432=>x"6f00", 433=>x"7100", 434=>x"7200",
--435=>x"7500", 436=>x"7800", 437=>x"7c00", 438=>x"8000", 439=>x"7600", 440=>x"7400", 441=>x"7900",
--442=>x"7700", 443=>x"7a00", 444=>x"7a00", 445=>x"7a00", 446=>x"7d00", 447=>x"7f00", 448=>x"7600",
--449=>x"7800", 450=>x"7b00", 451=>x"7600", 452=>x"7700", 453=>x"7d00", 454=>x"7f00", 455=>x"7b00",
--456=>x"6d00", 457=>x"7800", 458=>x"7700", 459=>x"7800", 460=>x"7d00", 461=>x"7c00", 462=>x"8200",
--463=>x"8000", 464=>x"7100", 465=>x"7700", 466=>x"7500", 467=>x"7500", 468=>x"7d00", 469=>x"8200",
--470=>x"8100", 471=>x"8400", 472=>x"7300", 473=>x"7c00", 474=>x"8900", 475=>x"7500", 476=>x"7d00",
--477=>x"8000", 478=>x"8400", 479=>x"7f00", 480=>x"7600", 481=>x"7800", 482=>x"7700", 483=>x"7900",
--484=>x"8200", 485=>x"7c00", 486=>x"8600", 487=>x"8300", 488=>x"7800", 489=>x"7000", 490=>x"7600",
--491=>x"7e00", 492=>x"8400", 493=>x"8500", 494=>x"8100", 495=>x"7600", 496=>x"7000", 497=>x"7700",
--498=>x"8000", 499=>x"8500"),
--11 => (0=>x"8600", 1=>x"8600", 2=>x"8500", 3=>x"8300", 4=>x"8500", 5=>x"8800", 6=>x"8400", 7=>x"7b00",
--8=>x"8600", 9=>x"8500", 10=>x"8600", 11=>x"8300", 12=>x"8500", 13=>x"8800", 14=>x"8500",
--15=>x"8400", 16=>x"8700", 17=>x"8600", 18=>x"8500", 19=>x"7c00", 20=>x"8500", 21=>x"8600",
--22=>x"8500", 23=>x"8400", 24=>x"8400", 25=>x"8500", 26=>x"8500", 27=>x"8300", 28=>x"8200",
--29=>x"8200", 30=>x"8200", 31=>x"8300", 32=>x"8200", 33=>x"8400", 34=>x"8700", 35=>x"8600",
--36=>x"8100", 37=>x"8600", 38=>x"8500", 39=>x"8400", 40=>x"7b00", 41=>x"8600", 42=>x"8600",
--43=>x"8100", 44=>x"8200", 45=>x"8500", 46=>x"8400", 47=>x"8300", 48=>x"8500", 49=>x"8400",
--50=>x"8200", 51=>x"8300", 52=>x"8500", 53=>x"8300", 54=>x"8300", 55=>x"8400", 56=>x"8300",
--57=>x"8200", 58=>x"8200", 59=>x"8500", 60=>x"8500", 61=>x"8400", 62=>x"8700", 63=>x"8200",
--64=>x"8700", 65=>x"8600", 66=>x"8500", 67=>x"8400", 68=>x"8400", 69=>x"8500", 70=>x"8600",
--71=>x"8400", 72=>x"8600", 73=>x"8700", 74=>x"8500", 75=>x"8300", 76=>x"8300", 77=>x"8300",
--78=>x"8500", 79=>x"8400", 80=>x"8400", 81=>x"8200", 82=>x"8100", 83=>x"8500", 84=>x"8200",
--85=>x"8200", 86=>x"8400", 87=>x"8200", 88=>x"8300", 89=>x"8200", 90=>x"8200", 91=>x"8200",
--92=>x"8100", 93=>x"8000", 94=>x"8500", 95=>x"8200", 96=>x"8400", 97=>x"8100", 98=>x"8200",
--99=>x"8100", 100=>x"8200", 101=>x"8000", 102=>x"8300", 103=>x"8300", 104=>x"8300", 105=>x"8300",
--106=>x"8100", 107=>x"8000", 108=>x"8100", 109=>x"8300", 110=>x"8400", 111=>x"8500", 112=>x"8300",
--113=>x"8200", 114=>x"8000", 115=>x"7d00", 116=>x"8100", 117=>x"8200", 118=>x"8100", 119=>x"8400",
--120=>x"8100", 121=>x"8200", 122=>x"8000", 123=>x"8000", 124=>x"8200", 125=>x"7c00", 126=>x"8100",
--127=>x"8400", 128=>x"7f00", 129=>x"8100", 130=>x"8400", 131=>x"8400", 132=>x"8100", 133=>x"7f00",
--134=>x"8300", 135=>x"8200", 136=>x"8000", 137=>x"8100", 138=>x"8100", 139=>x"8100", 140=>x"8000",
--141=>x"8100", 142=>x"8000", 143=>x"8100", 144=>x"8100", 145=>x"8200", 146=>x"8300", 147=>x"8200",
--148=>x"8100", 149=>x"8100", 150=>x"7f00", 151=>x"8100", 152=>x"8100", 153=>x"8100", 154=>x"8600",
--155=>x"8400", 156=>x"8300", 157=>x"8000", 158=>x"8000", 159=>x"7f00", 160=>x"8000", 161=>x"8000",
--162=>x"8200", 163=>x"7f00", 164=>x"8000", 165=>x"8100", 166=>x"7f00", 167=>x"8000", 168=>x"8300",
--169=>x"8100", 170=>x"8000", 171=>x"8000", 172=>x"8200", 173=>x"8000", 174=>x"7f00", 175=>x"8100",
--176=>x"8000", 177=>x"8100", 178=>x"8100", 179=>x"8200", 180=>x"8000", 181=>x"8100", 182=>x"7e00",
--183=>x"7e00", 184=>x"8200", 185=>x"8600", 186=>x"8200", 187=>x"7e00", 188=>x"8000", 189=>x"7f00",
--190=>x"8100", 191=>x"7f00", 192=>x"8200", 193=>x"8400", 194=>x"8100", 195=>x"8000", 196=>x"8000",
--197=>x"8000", 198=>x"8000", 199=>x"7e00", 200=>x"8700", 201=>x"7f00", 202=>x"8000", 203=>x"8100",
--204=>x"7f00", 205=>x"7f00", 206=>x"7c00", 207=>x"7a00", 208=>x"8200", 209=>x"8000", 210=>x"7f00",
--211=>x"7e00", 212=>x"7e00", 213=>x"7d00", 214=>x"8100", 215=>x"8800", 216=>x"7d00", 217=>x"7c00",
--218=>x"7d00", 219=>x"7f00", 220=>x"8000", 221=>x"8000", 222=>x"8a00", 223=>x"9500", 224=>x"8800",
--225=>x"8900", 226=>x"8800", 227=>x"8100", 228=>x"7f00", 229=>x"8600", 230=>x"9500", 231=>x"9100",
--232=>x"9400", 233=>x"8900", 234=>x"7d00", 235=>x"7500", 236=>x"7e00", 237=>x"8600", 238=>x"8b00",
--239=>x"8a00", 240=>x"8100", 241=>x"7e00", 242=>x"7900", 243=>x"7a00", 244=>x"7b00", 245=>x"7d00",
--246=>x"8400", 247=>x"8700", 248=>x"7f00", 249=>x"7d00", 250=>x"7900", 251=>x"7a00", 252=>x"7900",
--253=>x"7e00", 254=>x"8a00", 255=>x"8700", 256=>x"7c00", 257=>x"7a00", 258=>x"7d00", 259=>x"7c00",
--260=>x"7e00", 261=>x"8200", 262=>x"8800", 263=>x"8300", 264=>x"7a00", 265=>x"7900", 266=>x"7a00",
--267=>x"7600", 268=>x"7900", 269=>x"8500", 270=>x"8500", 271=>x"8400", 272=>x"8000", 273=>x"7a00",
--274=>x"7600", 275=>x"7700", 276=>x"7b00", 277=>x"7e00", 278=>x"8100", 279=>x"8500", 280=>x"7b00",
--281=>x"7c00", 282=>x"7600", 283=>x"7b00", 284=>x"8000", 285=>x"8400", 286=>x"8800", 287=>x"8600",
--288=>x"7900", 289=>x"7c00", 290=>x"8000", 291=>x"7e00", 292=>x"7900", 293=>x"8700", 294=>x"8100",
--295=>x"8200", 296=>x"7c00", 297=>x"8300", 298=>x"7d00", 299=>x"7700", 300=>x"8500", 301=>x"8100",
--302=>x"7500", 303=>x"8100", 304=>x"7b00", 305=>x"7a00", 306=>x"7a00", 307=>x"8000", 308=>x"7e00",
--309=>x"7a00", 310=>x"7f00", 311=>x"8300", 312=>x"7100", 313=>x"7b00", 314=>x"7e00", 315=>x"8100",
--316=>x"7900", 317=>x"7c00", 318=>x"8300", 319=>x"8300", 320=>x"7700", 321=>x"7e00", 322=>x"7c00",
--323=>x"7d00", 324=>x"7900", 325=>x"7f00", 326=>x"8000", 327=>x"8100", 328=>x"7c00", 329=>x"7600",
--330=>x"7d00", 331=>x"7800", 332=>x"7600", 333=>x"7d00", 334=>x"7800", 335=>x"7c00", 336=>x"7600",
--337=>x"7900", 338=>x"7a00", 339=>x"7500", 340=>x"7800", 341=>x"7800", 342=>x"7800", 343=>x"7a00",
--344=>x"7a00", 345=>x"7700", 346=>x"7800", 347=>x"7800", 348=>x"7400", 349=>x"7700", 350=>x"8000",
--351=>x"7d00", 352=>x"7800", 353=>x"7400", 354=>x"7300", 355=>x"7100", 356=>x"7400", 357=>x"7d00",
--358=>x"7d00", 359=>x"8400", 360=>x"6f00", 361=>x"7100", 362=>x"7400", 363=>x"7a00", 364=>x"7700",
--365=>x"7f00", 366=>x"8300", 367=>x"7900", 368=>x"6b00", 369=>x"6e00", 370=>x"7900", 371=>x"8000",
--372=>x"8000", 373=>x"8000", 374=>x"7d00", 375=>x"7f00", 376=>x"7100", 377=>x"7600", 378=>x"7800",
--379=>x"8000", 380=>x"8400", 381=>x"7e00", 382=>x"8100", 383=>x"8200", 384=>x"7700", 385=>x"7800",
--386=>x"7900", 387=>x"7c00", 388=>x"8100", 389=>x"8100", 390=>x"7f00", 391=>x"8500", 392=>x"7500",
--393=>x"7c00", 394=>x"7e00", 395=>x"8400", 396=>x"7f00", 397=>x"7a00", 398=>x"8100", 399=>x"8000",
--400=>x"7700", 401=>x"7c00", 402=>x"8200", 403=>x"8200", 404=>x"8000", 405=>x"7f00", 406=>x"7d00",
--407=>x"8600", 408=>x"8000", 409=>x"8900", 410=>x"8400", 411=>x"8100", 412=>x"7f00", 413=>x"8800",
--414=>x"8900", 415=>x"8b00", 416=>x"8400", 417=>x"8200", 418=>x"7f00", 419=>x"8600", 420=>x"8900",
--421=>x"8c00", 422=>x"9100", 423=>x"9000", 424=>x"7b00", 425=>x"8200", 426=>x"8900", 427=>x"8500",
--428=>x"8700", 429=>x"9000", 430=>x"9000", 431=>x"8c00", 432=>x"7d00", 433=>x"8300", 434=>x"8700",
--435=>x"8300", 436=>x"8c00", 437=>x"9400", 438=>x"8d00", 439=>x"8200", 440=>x"7e00", 441=>x"7e00",
--442=>x"8700", 443=>x"8d00", 444=>x"9200", 445=>x"8900", 446=>x"7f00", 447=>x"8200", 448=>x"8400",
--449=>x"8600", 450=>x"8f00", 451=>x"8b00", 452=>x"8500", 453=>x"8200", 454=>x"8800", 455=>x"8200",
--456=>x"8600", 457=>x"8700", 458=>x"8300", 459=>x"8600", 460=>x"8b00", 461=>x"8d00", 462=>x"8800",
--463=>x"8800", 464=>x"8b00", 465=>x"8a00", 466=>x"8400", 467=>x"8500", 468=>x"8f00", 469=>x"8d00",
--470=>x"8000", 471=>x"7f00", 472=>x"8a00", 473=>x"8d00", 474=>x"8300", 475=>x"8500", 476=>x"8500",
--477=>x"7d00", 478=>x"8100", 479=>x"8700", 480=>x"8000", 481=>x"7d00", 482=>x"8700", 483=>x"7800",
--484=>x"7300", 485=>x"8300", 486=>x"8900", 487=>x"8800", 488=>x"7c00", 489=>x"7e00", 490=>x"6c00",
--491=>x"7100", 492=>x"8700", 493=>x"8d00", 494=>x"8800", 495=>x"7b00", 496=>x"7700", 497=>x"7100",
--498=>x"8700", 499=>x"8700"),
--12 => (0=>x"8700", 1=>x"7900", 2=>x"8700", 3=>x"8700", 4=>x"8800", 5=>x"7a00", 6=>x"8800", 7=>x"8500",
--8=>x"8700", 9=>x"8600", 10=>x"8700", 11=>x"8800", 12=>x"8800", 13=>x"8600", 14=>x"8800",
--15=>x"8500", 16=>x"8700", 17=>x"8500", 18=>x"8700", 19=>x"8700", 20=>x"8700", 21=>x"8600",
--22=>x"8800", 23=>x"8500", 24=>x"8400", 25=>x"8600", 26=>x"8500", 27=>x"8400", 28=>x"8500",
--29=>x"8400", 30=>x"8400", 31=>x"8400", 32=>x"8500", 33=>x"8500", 34=>x"8300", 35=>x"8400",
--36=>x"8400", 37=>x"8200", 38=>x"8300", 39=>x"8200", 40=>x"8700", 41=>x"8400", 42=>x"8200",
--43=>x"8400", 44=>x"8300", 45=>x"8300", 46=>x"8400", 47=>x"8000", 48=>x"8200", 49=>x"8500",
--50=>x"8200", 51=>x"8300", 52=>x"8300", 53=>x"7d00", 54=>x"8400", 55=>x"8500", 56=>x"7f00",
--57=>x"8400", 58=>x"8400", 59=>x"8600", 60=>x"8400", 61=>x"8400", 62=>x"8400", 63=>x"8300",
--64=>x"8300", 65=>x"8300", 66=>x"8300", 67=>x"8600", 68=>x"8300", 69=>x"8100", 70=>x"8400",
--71=>x"8500", 72=>x"8500", 73=>x"8200", 74=>x"8200", 75=>x"8800", 76=>x"8600", 77=>x"8300",
--78=>x"8500", 79=>x"8500", 80=>x"8400", 81=>x"8100", 82=>x"8300", 83=>x"8600", 84=>x"8300",
--85=>x"8300", 86=>x"8100", 87=>x"8300", 88=>x"8200", 89=>x"8400", 90=>x"8100", 91=>x"8200",
--92=>x"8400", 93=>x"7f00", 94=>x"7f00", 95=>x"8400", 96=>x"8500", 97=>x"8400", 98=>x"8100",
--99=>x"8200", 100=>x"8200", 101=>x"8100", 102=>x"8000", 103=>x"8000", 104=>x"8a00", 105=>x"8600",
--106=>x"8500", 107=>x"8300", 108=>x"8300", 109=>x"7f00", 110=>x"7c00", 111=>x"7e00", 112=>x"8500",
--113=>x"8a00", 114=>x"8700", 115=>x"8300", 116=>x"8000", 117=>x"7b00", 118=>x"7c00", 119=>x"7e00",
--120=>x"8600", 121=>x"8400", 122=>x"7b00", 123=>x"8500", 124=>x"8200", 125=>x"8000", 126=>x"7d00",
--127=>x"7c00", 128=>x"8400", 129=>x"8300", 130=>x"8400", 131=>x"8100", 132=>x"8000", 133=>x"8200",
--134=>x"7f00", 135=>x"7c00", 136=>x"8500", 137=>x"8600", 138=>x"8400", 139=>x"8000", 140=>x"7d00",
--141=>x"7e00", 142=>x"7d00", 143=>x"7a00", 144=>x"7f00", 145=>x"8300", 146=>x"8100", 147=>x"7f00",
--148=>x"7b00", 149=>x"7f00", 150=>x"7e00", 151=>x"7c00", 152=>x"8400", 153=>x"7f00", 154=>x"7f00",
--155=>x"8100", 156=>x"7e00", 157=>x"7d00", 158=>x"7d00", 159=>x"7c00", 160=>x"8200", 161=>x"8100",
--162=>x"7d00", 163=>x"8000", 164=>x"7f00", 165=>x"7d00", 166=>x"7f00", 167=>x"7c00", 168=>x"8100",
--169=>x"8000", 170=>x"7e00", 171=>x"8000", 172=>x"7f00", 173=>x"7d00", 174=>x"8500", 175=>x"8100",
--176=>x"8200", 177=>x"8300", 178=>x"7e00", 179=>x"8000", 180=>x"7e00", 181=>x"7d00", 182=>x"7f00",
--183=>x"8100", 184=>x"8100", 185=>x"8800", 186=>x"8100", 187=>x"7b00", 188=>x"7d00", 189=>x"7b00",
--190=>x"7e00", 191=>x"7e00", 192=>x"7d00", 193=>x"7f00", 194=>x"8400", 195=>x"8600", 196=>x"8500",
--197=>x"8500", 198=>x"9200", 199=>x"7400", 200=>x"8100", 201=>x"8a00", 202=>x"8e00", 203=>x"9700",
--204=>x"9500", 205=>x"9600", 206=>x"9900", 207=>x"9b00", 208=>x"8f00", 209=>x"9500", 210=>x"9400",
--211=>x"9800", 212=>x"9500", 213=>x"8c00", 214=>x"9200", 215=>x"9400", 216=>x"8b00", 217=>x"8e00",
--218=>x"9300", 219=>x"9b00", 220=>x"8f00", 221=>x"8c00", 222=>x"8a00", 223=>x"9100", 224=>x"8a00",
--225=>x"9200", 226=>x"9400", 227=>x"9200", 228=>x"9100", 229=>x"9100", 230=>x"9000", 231=>x"9700",
--232=>x"8b00", 233=>x"9200", 234=>x"8e00", 235=>x"8e00", 236=>x"8b00", 237=>x"9300", 238=>x"9900",
--239=>x"9600", 240=>x"8900", 241=>x"8200", 242=>x"8400", 243=>x"8300", 244=>x"8d00", 245=>x"9500",
--246=>x"8d00", 247=>x"9300", 248=>x"8700", 249=>x"8100", 250=>x"7e00", 251=>x"8400", 252=>x"8f00",
--253=>x"8600", 254=>x"8600", 255=>x"8e00", 256=>x"8300", 257=>x"8200", 258=>x"7e00", 259=>x"8800",
--260=>x"7400", 261=>x"8a00", 262=>x"8900", 263=>x"8d00", 264=>x"8400", 265=>x"7e00", 266=>x"7f00",
--267=>x"8700", 268=>x"8700", 269=>x"8400", 270=>x"8b00", 271=>x"8700", 272=>x"7e00", 273=>x"8000",
--274=>x"8100", 275=>x"8200", 276=>x"8500", 277=>x"8900", 278=>x"8a00", 279=>x"8400", 280=>x"8000",
--281=>x"8600", 282=>x"8000", 283=>x"8600", 284=>x"8c00", 285=>x"8900", 286=>x"8100", 287=>x"8100",
--288=>x"8200", 289=>x"8900", 290=>x"8200", 291=>x"8b00", 292=>x"8c00", 293=>x"8200", 294=>x"7b00",
--295=>x"8700", 296=>x"8800", 297=>x"8700", 298=>x"8600", 299=>x"8c00", 300=>x"8100", 301=>x"8200",
--302=>x"8b00", 303=>x"8b00", 304=>x"8400", 305=>x"8100", 306=>x"8300", 307=>x"8800", 308=>x"8d00",
--309=>x"8b00", 310=>x"8d00", 311=>x"8800", 312=>x"8000", 313=>x"8000", 314=>x"7f00", 315=>x"8800",
--316=>x"8700", 317=>x"8400", 318=>x"8900", 319=>x"8100", 320=>x"7e00", 321=>x"7900", 322=>x"8100",
--323=>x"8500", 324=>x"8300", 325=>x"8600", 326=>x"8800", 327=>x"8a00", 328=>x"7f00", 329=>x"7e00",
--330=>x"8000", 331=>x"8700", 332=>x"8200", 333=>x"8100", 334=>x"8200", 335=>x"8400", 336=>x"8100",
--337=>x"8200", 338=>x"8600", 339=>x"8900", 340=>x"8a00", 341=>x"8700", 342=>x"7600", 343=>x"8700",
--344=>x"8500", 345=>x"8200", 346=>x"7c00", 347=>x"8e00", 348=>x"8900", 349=>x"8700", 350=>x"8c00",
--351=>x"8700", 352=>x"8000", 353=>x"8200", 354=>x"8700", 355=>x"8d00", 356=>x"8800", 357=>x"8200",
--358=>x"8900", 359=>x"8800", 360=>x"7c00", 361=>x"8700", 362=>x"8b00", 363=>x"8700", 364=>x"8100",
--365=>x"7400", 366=>x"8b00", 367=>x"8b00", 368=>x"8100", 369=>x"8c00", 370=>x"8d00", 371=>x"8900",
--372=>x"9100", 373=>x"8b00", 374=>x"8c00", 375=>x"8c00", 376=>x"8800", 377=>x"8a00", 378=>x"7200",
--379=>x"8a00", 380=>x"8a00", 381=>x"9000", 382=>x"9000", 383=>x"9000", 384=>x"8400", 385=>x"8700",
--386=>x"8200", 387=>x"8500", 388=>x"8f00", 389=>x"8c00", 390=>x"9000", 391=>x"9100", 392=>x"8d00",
--393=>x"8900", 394=>x"8700", 395=>x"8c00", 396=>x"8200", 397=>x"9000", 398=>x"8800", 399=>x"8e00",
--400=>x"8a00", 401=>x"8e00", 402=>x"8900", 403=>x"8700", 404=>x"7100", 405=>x"8f00", 406=>x"8c00",
--407=>x"8d00", 408=>x"8f00", 409=>x"8800", 410=>x"8d00", 411=>x"8c00", 412=>x"8600", 413=>x"8f00",
--414=>x"8800", 415=>x"8c00", 416=>x"8d00", 417=>x"8a00", 418=>x"8c00", 419=>x"8e00", 420=>x"8e00",
--421=>x"8700", 422=>x"8b00", 423=>x"8900", 424=>x"8600", 425=>x"8400", 426=>x"8c00", 427=>x"9000",
--428=>x"9100", 429=>x"8b00", 430=>x"9000", 431=>x"8b00", 432=>x"7b00", 433=>x"8c00", 434=>x"8700",
--435=>x"8c00", 436=>x"8f00", 437=>x"8900", 438=>x"8c00", 439=>x"8500", 440=>x"8a00", 441=>x"8200",
--442=>x"8c00", 443=>x"8c00", 444=>x"8900", 445=>x"8d00", 446=>x"8300", 447=>x"8100", 448=>x"8600",
--449=>x"8a00", 450=>x"8a00", 451=>x"8800", 452=>x"9000", 453=>x"8800", 454=>x"8600", 455=>x"7c00",
--456=>x"8400", 457=>x"8200", 458=>x"8b00", 459=>x"8e00", 460=>x"8a00", 461=>x"7700", 462=>x"7900",
--463=>x"7f00", 464=>x"8400", 465=>x"8b00", 466=>x"8d00", 467=>x"8200", 468=>x"7300", 469=>x"7100",
--470=>x"7900", 471=>x"7200", 472=>x"8b00", 473=>x"8b00", 474=>x"7f00", 475=>x"7300", 476=>x"7600",
--477=>x"7100", 478=>x"6400", 479=>x"7200", 480=>x"8800", 481=>x"7c00", 482=>x"8100", 483=>x"7e00",
--484=>x"7100", 485=>x"6500", 486=>x"7400", 487=>x"9d00", 488=>x"8000", 489=>x"7d00", 490=>x"7900",
--491=>x"6f00", 492=>x"6800", 493=>x"7e00", 494=>x"9f00", 495=>x"a300", 496=>x"7a00", 497=>x"7100",
--498=>x"6d00", 499=>x"6200"),
--13 => (0=>x"8700", 1=>x"8600", 2=>x"8700", 3=>x"8200", 4=>x"8100", 5=>x"8200", 6=>x"7b00", 7=>x"8200",
--8=>x"8700", 9=>x"8600", 10=>x"8700", 11=>x"7d00", 12=>x"8300", 13=>x"8200", 14=>x"8400",
--15=>x"8100", 16=>x"8600", 17=>x"8600", 18=>x"8500", 19=>x"7e00", 20=>x"8100", 21=>x"8200",
--22=>x"8600", 23=>x"8300", 24=>x"8600", 25=>x"8500", 26=>x"8700", 27=>x"7e00", 28=>x"8200",
--29=>x"8100", 30=>x"8200", 31=>x"8200", 32=>x"8300", 33=>x"8200", 34=>x"8500", 35=>x"8500",
--36=>x"8300", 37=>x"8000", 38=>x"7f00", 39=>x"7f00", 40=>x"8100", 41=>x"8500", 42=>x"8200",
--43=>x"8100", 44=>x"8200", 45=>x"8200", 46=>x"8000", 47=>x"8000", 48=>x"8600", 49=>x"8500",
--50=>x"8400", 51=>x"8400", 52=>x"8200", 53=>x"8100", 54=>x"8200", 55=>x"8200", 56=>x"8200",
--57=>x"8300", 58=>x"8300", 59=>x"8300", 60=>x"8200", 61=>x"8100", 62=>x"8500", 63=>x"8200",
--64=>x"8600", 65=>x"8500", 66=>x"8600", 67=>x"8200", 68=>x"8600", 69=>x"8500", 70=>x"8400",
--71=>x"7f00", 72=>x"8300", 73=>x"8300", 74=>x"8500", 75=>x"8400", 76=>x"8900", 77=>x"8200",
--78=>x"8200", 79=>x"8100", 80=>x"8700", 81=>x"8200", 82=>x"8100", 83=>x"8200", 84=>x"8300",
--85=>x"8200", 86=>x"8700", 87=>x"8300", 88=>x"8500", 89=>x"7e00", 90=>x"8100", 91=>x"8100",
--92=>x"8000", 93=>x"8200", 94=>x"8100", 95=>x"8000", 96=>x"7e00", 97=>x"7f00", 98=>x"8000",
--99=>x"7e00", 100=>x"7f00", 101=>x"7f00", 102=>x"7e00", 103=>x"8100", 104=>x"7e00", 105=>x"7d00",
--106=>x"7c00", 107=>x"7e00", 108=>x"7f00", 109=>x"8000", 110=>x"7e00", 111=>x"8000", 112=>x"7c00",
--113=>x"7900", 114=>x"7b00", 115=>x"7b00", 116=>x"7c00", 117=>x"7e00", 118=>x"8200", 119=>x"8100",
--120=>x"7b00", 121=>x"7900", 122=>x"7b00", 123=>x"8500", 124=>x"7c00", 125=>x"7c00", 126=>x"7e00",
--127=>x"8000", 128=>x"7b00", 129=>x"7a00", 130=>x"7c00", 131=>x"7900", 132=>x"7c00", 133=>x"7900",
--134=>x"7900", 135=>x"8000", 136=>x"7b00", 137=>x"7d00", 138=>x"7900", 139=>x"7600", 140=>x"7a00",
--141=>x"7900", 142=>x"7c00", 143=>x"7d00", 144=>x"7c00", 145=>x"7d00", 146=>x"7c00", 147=>x"7900",
--148=>x"7d00", 149=>x"7b00", 150=>x"7d00", 151=>x"7e00", 152=>x"7c00", 153=>x"7b00", 154=>x"7800",
--155=>x"7a00", 156=>x"7d00", 157=>x"7900", 158=>x"7a00", 159=>x"7d00", 160=>x"8100", 161=>x"7b00",
--162=>x"7a00", 163=>x"7c00", 164=>x"7d00", 165=>x"7b00", 166=>x"7600", 167=>x"7700", 168=>x"7e00",
--169=>x"7d00", 170=>x"7f00", 171=>x"7d00", 172=>x"7b00", 173=>x"7a00", 174=>x"7a00", 175=>x"7400",
--176=>x"7f00", 177=>x"7c00", 178=>x"7a00", 179=>x"7b00", 180=>x"7900", 181=>x"7b00", 182=>x"7e00",
--183=>x"8b00", 184=>x"8700", 185=>x"8a00", 186=>x"8800", 187=>x"8700", 188=>x"8500", 189=>x"9000",
--190=>x"9e00", 191=>x"ac00", 192=>x"9700", 193=>x"9100", 194=>x"9100", 195=>x"6900", 196=>x"a000",
--197=>x"a400", 198=>x"5500", 199=>x"aa00", 200=>x"9300", 201=>x"9100", 202=>x"9a00", 203=>x"a800",
--204=>x"5500", 205=>x"a300", 206=>x"a700", 207=>x"ab00", 208=>x"9200", 209=>x"9900", 210=>x"a400",
--211=>x"ac00", 212=>x"aa00", 213=>x"a700", 214=>x"a800", 215=>x"ac00", 216=>x"9600", 217=>x"9800",
--218=>x"9d00", 219=>x"a800", 220=>x"a000", 221=>x"a300", 222=>x"aa00", 223=>x"ab00", 224=>x"9600",
--225=>x"9300", 226=>x"9800", 227=>x"9900", 228=>x"a000", 229=>x"9f00", 230=>x"a000", 231=>x"a500",
--232=>x"9500", 233=>x"9300", 234=>x"9700", 235=>x"9c00", 236=>x"9c00", 237=>x"9f00", 238=>x"a600",
--239=>x"a500", 240=>x"9700", 241=>x"9500", 242=>x"9900", 243=>x"9900", 244=>x"9800", 245=>x"a100",
--246=>x"aa00", 247=>x"a500", 248=>x"9500", 249=>x"9b00", 250=>x"9800", 251=>x"9600", 252=>x"9c00",
--253=>x"a800", 254=>x"a000", 255=>x"a000", 256=>x"9300", 257=>x"9500", 258=>x"9000", 259=>x"9900",
--260=>x"9e00", 261=>x"a000", 262=>x"9e00", 263=>x"9800", 264=>x"8c00", 265=>x"9000", 266=>x"8f00",
--267=>x"9400", 268=>x"9900", 269=>x"9800", 270=>x"9800", 271=>x"9b00", 272=>x"8c00", 273=>x"8c00",
--274=>x"9200", 275=>x"8e00", 276=>x"9200", 277=>x"9a00", 278=>x"9c00", 279=>x"a200", 280=>x"8900",
--281=>x"8600", 282=>x"8200", 283=>x"8f00", 284=>x"9100", 285=>x"9900", 286=>x"9d00", 287=>x"a200",
--288=>x"8d00", 289=>x"8d00", 290=>x"8c00", 291=>x"9100", 292=>x"9300", 293=>x"9000", 294=>x"9900",
--295=>x"a000", 296=>x"8600", 297=>x"8e00", 298=>x"8a00", 299=>x"8e00", 300=>x"8c00", 301=>x"9700",
--302=>x"9500", 303=>x"9900", 304=>x"8500", 305=>x"8800", 306=>x"8500", 307=>x"8900", 308=>x"9800",
--309=>x"6800", 310=>x"9300", 311=>x"9700", 312=>x"7400", 313=>x"8f00", 314=>x"8400", 315=>x"8f00",
--316=>x"9400", 317=>x"9100", 318=>x"9200", 319=>x"9600", 320=>x"8100", 321=>x"7900", 322=>x"8700",
--323=>x"9500", 324=>x"8d00", 325=>x"9000", 326=>x"9700", 327=>x"9800", 328=>x"8700", 329=>x"8200",
--330=>x"8d00", 331=>x"8f00", 332=>x"8800", 333=>x"8800", 334=>x"9300", 335=>x"9800", 336=>x"8200",
--337=>x"8a00", 338=>x"8600", 339=>x"8c00", 340=>x"8600", 341=>x"8b00", 342=>x"9300", 343=>x"8c00",
--344=>x"8800", 345=>x"8400", 346=>x"8f00", 347=>x"8c00", 348=>x"8c00", 349=>x"8d00", 350=>x"9000",
--351=>x"9f00", 352=>x"8500", 353=>x"9100", 354=>x"8b00", 355=>x"8d00", 356=>x"8e00", 357=>x"8d00",
--358=>x"9500", 359=>x"9400", 360=>x"8d00", 361=>x"8f00", 362=>x"8d00", 363=>x"8e00", 364=>x"9300",
--365=>x"9800", 366=>x"9100", 367=>x"9100", 368=>x"8b00", 369=>x"9300", 370=>x"9300", 371=>x"9100",
--372=>x"8f00", 373=>x"8d00", 374=>x"9000", 375=>x"9000", 376=>x"9400", 377=>x"9300", 378=>x"8f00",
--379=>x"8100", 380=>x"8e00", 381=>x"8900", 382=>x"8d00", 383=>x"9400", 384=>x"9500", 385=>x"9000",
--386=>x"8600", 387=>x"8a00", 388=>x"9000", 389=>x"8800", 390=>x"9100", 391=>x"6e00", 392=>x"9200",
--393=>x"8700", 394=>x"8e00", 395=>x"8b00", 396=>x"8c00", 397=>x"8e00", 398=>x"9100", 399=>x"9200",
--400=>x"8800", 401=>x"8c00", 402=>x"8400", 403=>x"8400", 404=>x"8800", 405=>x"8800", 406=>x"8f00",
--407=>x"8d00", 408=>x"8700", 409=>x"8500", 410=>x"8700", 411=>x"8100", 412=>x"8900", 413=>x"8d00",
--414=>x"8b00", 415=>x"9100", 416=>x"8500", 417=>x"8a00", 418=>x"8900", 419=>x"8500", 420=>x"8700",
--421=>x"8d00", 422=>x"8d00", 423=>x"8200", 424=>x"8400", 425=>x"8500", 426=>x"8200", 427=>x"7d00",
--428=>x"8500", 429=>x"8200", 430=>x"7e00", 431=>x"7a00", 432=>x"8500", 433=>x"8200", 434=>x"7800",
--435=>x"8200", 436=>x"8200", 437=>x"7600", 438=>x"7e00", 439=>x"9c00", 440=>x"8300", 441=>x"8000",
--442=>x"7900", 443=>x"6f00", 444=>x"6d00", 445=>x"8100", 446=>x"a400", 447=>x"ad00", 448=>x"7e00",
--449=>x"7b00", 450=>x"6900", 451=>x"6e00", 452=>x"9000", 453=>x"b100", 454=>x"b800", 455=>x"b000",
--456=>x"7900", 457=>x"6a00", 458=>x"7500", 459=>x"9700", 460=>x"a700", 461=>x"b600", 462=>x"ba00",
--463=>x"c100", 464=>x"6e00", 465=>x"7f00", 466=>x"a600", 467=>x"b300", 468=>x"a500", 469=>x"b300",
--470=>x"c700", 471=>x"c000", 472=>x"9000", 473=>x"a500", 474=>x"a500", 475=>x"b400", 476=>x"b900",
--477=>x"b200", 478=>x"c300", 479=>x"b300", 480=>x"ad00", 481=>x"ab00", 482=>x"ae00", 483=>x"bd00",
--484=>x"b400", 485=>x"a600", 486=>x"b100", 487=>x"b400", 488=>x"af00", 489=>x"b700", 490=>x"b500",
--491=>x"b400", 492=>x"a800", 493=>x"a000", 494=>x"a100", 495=>x"a900", 496=>x"b500", 497=>x"b800",
--498=>x"a900", 499=>x"a900"),
--14 => (0=>x"8200", 1=>x"8500", 2=>x"8700", 3=>x"8400", 4=>x"8400", 5=>x"8400", 6=>x"8300", 7=>x"8400",
--8=>x"8200", 9=>x"8500", 10=>x"8600", 11=>x"8400", 12=>x"8400", 13=>x"8400", 14=>x"8300",
--15=>x"8400", 16=>x"8200", 17=>x"8100", 18=>x"8600", 19=>x"8400", 20=>x"8200", 21=>x"8300",
--22=>x"8200", 23=>x"8300", 24=>x"8100", 25=>x"8300", 26=>x"8700", 27=>x"8200", 28=>x"8100",
--29=>x"8000", 30=>x"7e00", 31=>x"8400", 32=>x"8200", 33=>x"8700", 34=>x"8500", 35=>x"8400",
--36=>x"8200", 37=>x"8000", 38=>x"8100", 39=>x"8400", 40=>x"8200", 41=>x"8100", 42=>x"8100",
--43=>x"8200", 44=>x"8000", 45=>x"8100", 46=>x"8200", 47=>x"8100", 48=>x"8200", 49=>x"8100",
--50=>x"8300", 51=>x"8400", 52=>x"8100", 53=>x"8000", 54=>x"8200", 55=>x"8300", 56=>x"8100",
--57=>x"8400", 58=>x"8200", 59=>x"8200", 60=>x"8000", 61=>x"7f00", 62=>x"8300", 63=>x"8200",
--64=>x"7e00", 65=>x"8400", 66=>x"8400", 67=>x"8400", 68=>x"8100", 69=>x"8100", 70=>x"8200",
--71=>x"8300", 72=>x"7f00", 73=>x"8400", 74=>x"8500", 75=>x"8300", 76=>x"8100", 77=>x"7f00",
--78=>x"8100", 79=>x"8400", 80=>x"8300", 81=>x"8300", 82=>x"8200", 83=>x"8300", 84=>x"8000",
--85=>x"7f00", 86=>x"8000", 87=>x"8200", 88=>x"8400", 89=>x"8200", 90=>x"8000", 91=>x"8100",
--92=>x"8000", 93=>x"7f00", 94=>x"8000", 95=>x"8000", 96=>x"7f00", 97=>x"8000", 98=>x"7f00",
--99=>x"8000", 100=>x"8000", 101=>x"7e00", 102=>x"7d00", 103=>x"8000", 104=>x"8000", 105=>x"7d00",
--106=>x"7e00", 107=>x"7e00", 108=>x"8000", 109=>x"7d00", 110=>x"7c00", 111=>x"7e00", 112=>x"7d00",
--113=>x"7d00", 114=>x"7c00", 115=>x"7c00", 116=>x"8300", 117=>x"7e00", 118=>x"7f00", 119=>x"7f00",
--120=>x"7f00", 121=>x"7e00", 122=>x"7d00", 123=>x"7f00", 124=>x"7c00", 125=>x"7b00", 126=>x"7e00",
--127=>x"7f00", 128=>x"7d00", 129=>x"7b00", 130=>x"7d00", 131=>x"7e00", 132=>x"7e00", 133=>x"7e00",
--134=>x"7c00", 135=>x"7c00", 136=>x"7d00", 137=>x"8100", 138=>x"7d00", 139=>x"7a00", 140=>x"7a00",
--141=>x"7c00", 142=>x"7a00", 143=>x"7c00", 144=>x"7c00", 145=>x"7f00", 146=>x"7b00", 147=>x"7900",
--148=>x"7a00", 149=>x"7700", 150=>x"7700", 151=>x"7c00", 152=>x"7d00", 153=>x"7900", 154=>x"7700",
--155=>x"7800", 156=>x"7800", 157=>x"7600", 158=>x"7900", 159=>x"7900", 160=>x"7900", 161=>x"7800",
--162=>x"7800", 163=>x"7900", 164=>x"7900", 165=>x"7700", 166=>x"7900", 167=>x"7800", 168=>x"7400",
--169=>x"7700", 170=>x"7500", 171=>x"7600", 172=>x"7400", 173=>x"7700", 174=>x"7500", 175=>x"7500",
--176=>x"8a00", 177=>x"8800", 178=>x"8900", 179=>x"8000", 180=>x"7d00", 181=>x"7b00", 182=>x"7400",
--183=>x"7200", 184=>x"a400", 185=>x"b100", 186=>x"ac00", 187=>x"a800", 188=>x"aa00", 189=>x"ab00",
--190=>x"a300", 191=>x"9f00", 192=>x"b000", 193=>x"ac00", 194=>x"ab00", 195=>x"b100", 196=>x"b700",
--197=>x"b800", 198=>x"bc00", 199=>x"bc00", 200=>x"b200", 201=>x"b600", 202=>x"b200", 203=>x"b100",
--204=>x"b000", 205=>x"b800", 206=>x"b100", 207=>x"b400", 208=>x"b400", 209=>x"b700", 210=>x"b500",
--211=>x"b200", 212=>x"b300", 213=>x"ae00", 214=>x"a700", 215=>x"aa00", 216=>x"b100", 217=>x"b200",
--218=>x"b500", 219=>x"b400", 220=>x"b000", 221=>x"ac00", 222=>x"ac00", 223=>x"ac00", 224=>x"a300",
--225=>x"ae00", 226=>x"b500", 227=>x"b300", 228=>x"b000", 229=>x"b300", 230=>x"b100", 231=>x"af00",
--232=>x"a600", 233=>x"a300", 234=>x"b000", 235=>x"af00", 236=>x"a700", 237=>x"af00", 238=>x"4b00",
--239=>x"b100", 240=>x"5900", 241=>x"ac00", 242=>x"a700", 243=>x"a300", 244=>x"aa00", 245=>x"b200",
--246=>x"b400", 247=>x"b100", 248=>x"a600", 249=>x"a700", 250=>x"a700", 251=>x"ab00", 252=>x"af00",
--253=>x"b500", 254=>x"b400", 255=>x"b200", 256=>x"a200", 257=>x"a000", 258=>x"ae00", 259=>x"ad00",
--260=>x"ac00", 261=>x"b000", 262=>x"b600", 263=>x"bd00", 264=>x"ab00", 265=>x"ae00", 266=>x"ab00",
--267=>x"a900", 268=>x"ae00", 269=>x"b100", 270=>x"b800", 271=>x"ba00", 272=>x"a500", 273=>x"ae00",
--274=>x"af00", 275=>x"b000", 276=>x"5000", 277=>x"b200", 278=>x"b400", 279=>x"b400", 280=>x"a300",
--281=>x"5200", 282=>x"af00", 283=>x"b200", 284=>x"ae00", 285=>x"af00", 286=>x"b500", 287=>x"ae00",
--288=>x"a400", 289=>x"a800", 290=>x"a700", 291=>x"ac00", 292=>x"ab00", 293=>x"ae00", 294=>x"b300",
--295=>x"b600", 296=>x"9f00", 297=>x"a100", 298=>x"a200", 299=>x"a500", 300=>x"a800", 301=>x"af00",
--302=>x"b600", 303=>x"b500", 304=>x"9b00", 305=>x"9e00", 306=>x"9f00", 307=>x"ac00", 308=>x"ac00",
--309=>x"b300", 310=>x"b500", 311=>x"b300", 312=>x"9b00", 313=>x"a100", 314=>x"a700", 315=>x"aa00",
--316=>x"ae00", 317=>x"4900", 318=>x"b600", 319=>x"b900", 320=>x"a200", 321=>x"9800", 322=>x"a400",
--323=>x"b000", 324=>x"b000", 325=>x"b500", 326=>x"be00", 327=>x"bc00", 328=>x"9700", 329=>x"a100",
--330=>x"a600", 331=>x"a600", 332=>x"b300", 333=>x"be00", 334=>x"b300", 335=>x"b400", 336=>x"9f00",
--337=>x"6300", 338=>x"a300", 339=>x"ab00", 340=>x"ac00", 341=>x"b600", 342=>x"ba00", 343=>x"ba00",
--344=>x"9b00", 345=>x"9d00", 346=>x"a800", 347=>x"a500", 348=>x"b000", 349=>x"bc00", 350=>x"af00",
--351=>x"b200", 352=>x"9d00", 353=>x"9800", 354=>x"a300", 355=>x"ab00", 356=>x"a700", 357=>x"ad00",
--358=>x"b700", 359=>x"b600", 360=>x"9600", 361=>x"9c00", 362=>x"a300", 363=>x"9c00", 364=>x"ab00",
--365=>x"b700", 366=>x"b100", 367=>x"b000", 368=>x"9400", 369=>x"9800", 370=>x"a200", 371=>x"ac00",
--372=>x"ae00", 373=>x"4f00", 374=>x"b500", 375=>x"b200", 376=>x"9100", 377=>x"9b00", 378=>x"a700",
--379=>x"a300", 380=>x"af00", 381=>x"af00", 382=>x"ab00", 383=>x"9a00", 384=>x"9c00", 385=>x"9b00",
--386=>x"a000", 387=>x"5300", 388=>x"b200", 389=>x"9b00", 390=>x"8800", 391=>x"9300", 392=>x"9000",
--393=>x"9900", 394=>x"ac00", 395=>x"a900", 396=>x"9100", 397=>x"7e00", 398=>x"9800", 399=>x"ba00",
--400=>x"9400", 401=>x"a100", 402=>x"a200", 403=>x"8e00", 404=>x"8500", 405=>x"a500", 406=>x"c700",
--407=>x"c100", 408=>x"8700", 409=>x"9000", 410=>x"8600", 411=>x"8c00", 412=>x"b200", 413=>x"c600",
--414=>x"c700", 415=>x"3a00", 416=>x"8000", 417=>x"8200", 418=>x"6600", 419=>x"b100", 420=>x"c200",
--421=>x"be00", 422=>x"c600", 423=>x"c600", 424=>x"8d00", 425=>x"b300", 426=>x"b900", 427=>x"b000",
--428=>x"b500", 429=>x"c500", 430=>x"c500", 431=>x"ca00", 432=>x"ae00", 433=>x"c300", 434=>x"ba00",
--435=>x"b500", 436=>x"bc00", 437=>x"c000", 438=>x"c300", 439=>x"c100", 440=>x"b500", 441=>x"b900",
--442=>x"c700", 443=>x"bf00", 444=>x"bf00", 445=>x"b700", 446=>x"bb00", 447=>x"b900", 448=>x"ba00",
--449=>x"4000", 450=>x"c200", 451=>x"3d00", 452=>x"b500", 453=>x"b900", 454=>x"b400", 455=>x"bd00",
--456=>x"b800", 457=>x"b900", 458=>x"b700", 459=>x"b700", 460=>x"bd00", 461=>x"bb00", 462=>x"c100",
--463=>x"b800", 464=>x"b900", 465=>x"ad00", 466=>x"ad00", 467=>x"ae00", 468=>x"be00", 469=>x"c400",
--470=>x"bf00", 471=>x"af00", 472=>x"b000", 473=>x"b200", 474=>x"ad00", 475=>x"b100", 476=>x"b700",
--477=>x"b100", 478=>x"ad00", 479=>x"b800", 480=>x"ab00", 481=>x"b100", 482=>x"b900", 483=>x"ae00",
--484=>x"a000", 485=>x"a300", 486=>x"b900", 487=>x"bd00", 488=>x"bb00", 489=>x"ba00", 490=>x"a900",
--491=>x"a800", 492=>x"b100", 493=>x"b700", 494=>x"b000", 495=>x"b400", 496=>x"ac00", 497=>x"a600",
--498=>x"ac00", 499=>x"bd00"),
--15 => (0=>x"8600", 1=>x"8500", 2=>x"8500", 3=>x"8700", 4=>x"8500", 5=>x"8400", 6=>x"8200", 7=>x"8500",
--8=>x"8600", 9=>x"8400", 10=>x"8600", 11=>x"8800", 12=>x"8500", 13=>x"8400", 14=>x"8100",
--15=>x"8500", 16=>x"8700", 17=>x"8500", 18=>x"8500", 19=>x"8700", 20=>x"8500", 21=>x"8400",
--22=>x"8200", 23=>x"8500", 24=>x"8400", 25=>x"8500", 26=>x"8600", 27=>x"8200", 28=>x"8400",
--29=>x"8300", 30=>x"8300", 31=>x"8400", 32=>x"8300", 33=>x"8400", 34=>x"8300", 35=>x"8300",
--36=>x"8000", 37=>x"8200", 38=>x"8300", 39=>x"8400", 40=>x"8200", 41=>x"8100", 42=>x"8400",
--43=>x"8400", 44=>x"8200", 45=>x"8200", 46=>x"8000", 47=>x"7f00", 48=>x"8500", 49=>x"8700",
--50=>x"8800", 51=>x"8500", 52=>x"8400", 53=>x"8300", 54=>x"8300", 55=>x"8100", 56=>x"8400",
--57=>x"8600", 58=>x"8600", 59=>x"8600", 60=>x"8500", 61=>x"8100", 62=>x"8400", 63=>x"8400",
--64=>x"8400", 65=>x"8800", 66=>x"8500", 67=>x"8900", 68=>x"8700", 69=>x"8100", 70=>x"8600",
--71=>x"8200", 72=>x"8600", 73=>x"8800", 74=>x"8700", 75=>x"8800", 76=>x"8700", 77=>x"8400",
--78=>x"8400", 79=>x"8300", 80=>x"8200", 81=>x"8400", 82=>x"8700", 83=>x"8900", 84=>x"8c00",
--85=>x"8700", 86=>x"8400", 87=>x"8300", 88=>x"8300", 89=>x"8300", 90=>x"8500", 91=>x"8600",
--92=>x"8800", 93=>x"8300", 94=>x"8400", 95=>x"8200", 96=>x"8400", 97=>x"8200", 98=>x"8200",
--99=>x"8200", 100=>x"8300", 101=>x"8500", 102=>x"8300", 103=>x"8200", 104=>x"7c00", 105=>x"8000",
--106=>x"8000", 107=>x"8200", 108=>x"8400", 109=>x"8300", 110=>x"8400", 111=>x"8200", 112=>x"7f00",
--113=>x"8200", 114=>x"8100", 115=>x"7e00", 116=>x"8200", 117=>x"8200", 118=>x"8200", 119=>x"8400",
--120=>x"7f00", 121=>x"8200", 122=>x"8400", 123=>x"8100", 124=>x"8000", 125=>x"8000", 126=>x"8000",
--127=>x"8300", 128=>x"7d00", 129=>x"7e00", 130=>x"8300", 131=>x"8000", 132=>x"8100", 133=>x"8100",
--134=>x"8000", 135=>x"7f00", 136=>x"7b00", 137=>x"7e00", 138=>x"8100", 139=>x"8000", 140=>x"8100",
--141=>x"8300", 142=>x"8100", 143=>x"8000", 144=>x"7c00", 145=>x"7c00", 146=>x"8200", 147=>x"8100",
--148=>x"7f00", 149=>x"8100", 150=>x"8400", 151=>x"8200", 152=>x"7d00", 153=>x"7d00", 154=>x"7d00",
--155=>x"7f00", 156=>x"8000", 157=>x"7e00", 158=>x"8100", 159=>x"8100", 160=>x"7a00", 161=>x"7900",
--162=>x"7d00", 163=>x"8000", 164=>x"7e00", 165=>x"7f00", 166=>x"8500", 167=>x"8100", 168=>x"7800",
--169=>x"7800", 170=>x"7c00", 171=>x"7d00", 172=>x"7d00", 173=>x"8000", 174=>x"8100", 175=>x"8100",
--176=>x"7500", 177=>x"7400", 178=>x"7900", 179=>x"7c00", 180=>x"7900", 181=>x"7900", 182=>x"7d00",
--183=>x"7f00", 184=>x"8b00", 185=>x"8300", 186=>x"7500", 187=>x"7300", 188=>x"7300", 189=>x"7500",
--190=>x"7700", 191=>x"7800", 192=>x"bd00", 193=>x"b100", 194=>x"a100", 195=>x"9900", 196=>x"8400",
--197=>x"7900", 198=>x"7200", 199=>x"7300", 200=>x"b200", 201=>x"b600", 202=>x"c300", 203=>x"c200",
--204=>x"ba00", 205=>x"aa00", 206=>x"9500", 207=>x"8400", 208=>x"b100", 209=>x"b700", 210=>x"b400",
--211=>x"ba00", 212=>x"ba00", 213=>x"c200", 214=>x"c500", 215=>x"b700", 216=>x"5000", 217=>x"b600",
--218=>x"b400", 219=>x"b600", 220=>x"b800", 221=>x"be00", 222=>x"bb00", 223=>x"c300", 224=>x"b200",
--225=>x"b400", 226=>x"b400", 227=>x"b400", 228=>x"b400", 229=>x"ba00", 230=>x"bf00", 231=>x"bd00",
--232=>x"ad00", 233=>x"b500", 234=>x"b700", 235=>x"ba00", 236=>x"bc00", 237=>x"b900", 238=>x"c000",
--239=>x"bf00", 240=>x"5200", 241=>x"b700", 242=>x"ba00", 243=>x"bb00", 244=>x"bb00", 245=>x"bd00",
--246=>x"bf00", 247=>x"4000", 248=>x"b700", 249=>x"b900", 250=>x"b800", 251=>x"bc00", 252=>x"4800",
--253=>x"b700", 254=>x"bf00", 255=>x"bc00", 256=>x"be00", 257=>x"ba00", 258=>x"b600", 259=>x"b700",
--260=>x"b700", 261=>x"bd00", 262=>x"c000", 263=>x"bb00", 264=>x"b300", 265=>x"b900", 266=>x"bb00",
--267=>x"b800", 268=>x"bb00", 269=>x"be00", 270=>x"bd00", 271=>x"b800", 272=>x"b500", 273=>x"b900",
--274=>x"bb00", 275=>x"b600", 276=>x"bd00", 277=>x"bb00", 278=>x"bb00", 279=>x"bf00", 280=>x"b000",
--281=>x"ba00", 282=>x"b400", 283=>x"b200", 284=>x"b800", 285=>x"bf00", 286=>x"be00", 287=>x"3f00",
--288=>x"b900", 289=>x"b500", 290=>x"b500", 291=>x"bc00", 292=>x"c000", 293=>x"bf00", 294=>x"bf00",
--295=>x"c400", 296=>x"b700", 297=>x"b700", 298=>x"bb00", 299=>x"bc00", 300=>x"c000", 301=>x"c100",
--302=>x"bf00", 303=>x"bd00", 304=>x"b800", 305=>x"b800", 306=>x"bc00", 307=>x"b900", 308=>x"ba00",
--309=>x"c000", 310=>x"c000", 311=>x"be00", 312=>x"bd00", 313=>x"be00", 314=>x"b300", 315=>x"bc00",
--316=>x"be00", 317=>x"b700", 318=>x"be00", 319=>x"be00", 320=>x"b600", 321=>x"ba00", 322=>x"bb00",
--323=>x"b700", 324=>x"b900", 325=>x"be00", 326=>x"be00", 327=>x"c000", 328=>x"bc00", 329=>x"bb00",
--330=>x"b400", 331=>x"bc00", 332=>x"be00", 333=>x"b800", 334=>x"b900", 335=>x"c100", 336=>x"bb00",
--337=>x"b800", 338=>x"3c00", 339=>x"c100", 340=>x"b800", 341=>x"bd00", 342=>x"bd00", 343=>x"b800",
--344=>x"4400", 345=>x"ba00", 346=>x"bb00", 347=>x"c000", 348=>x"c200", 349=>x"ac00", 350=>x"a300",
--351=>x"a800", 352=>x"af00", 353=>x"b700", 354=>x"bc00", 355=>x"b300", 356=>x"aa00", 357=>x"9d00",
--358=>x"ac00", 359=>x"c200", 360=>x"b600", 361=>x"bd00", 362=>x"a000", 363=>x"9700", 364=>x"a400",
--365=>x"b800", 366=>x"ce00", 367=>x"d000", 368=>x"a700", 369=>x"9d00", 370=>x"9900", 371=>x"b700",
--372=>x"ca00", 373=>x"cd00", 374=>x"cb00", 375=>x"d000", 376=>x"8d00", 377=>x"9d00", 378=>x"bf00",
--379=>x"d200", 380=>x"cf00", 381=>x"d000", 382=>x"cb00", 383=>x"c600", 384=>x"aa00", 385=>x"c700",
--386=>x"cb00", 387=>x"cb00", 388=>x"ca00", 389=>x"ca00", 390=>x"cb00", 391=>x"c800", 392=>x"c400",
--393=>x"c400", 394=>x"cb00", 395=>x"c900", 396=>x"c300", 397=>x"cb00", 398=>x"d000", 399=>x"d100",
--400=>x"c000", 401=>x"c200", 402=>x"c100", 403=>x"cc00", 404=>x"ca00", 405=>x"c500", 406=>x"cf00",
--407=>x"ce00", 408=>x"bf00", 409=>x"c200", 410=>x"c700", 411=>x"c000", 412=>x"c600", 413=>x"c300",
--414=>x"c300", 415=>x"c400", 416=>x"c800", 417=>x"be00", 418=>x"c300", 419=>x"c200", 420=>x"bb00",
--421=>x"c100", 422=>x"c100", 423=>x"be00", 424=>x"c100", 425=>x"c200", 426=>x"bb00", 427=>x"c300",
--428=>x"c100", 429=>x"b800", 430=>x"c400", 431=>x"c300", 432=>x"be00", 433=>x"bf00", 434=>x"c300",
--435=>x"b900", 436=>x"c000", 437=>x"c200", 438=>x"b800", 439=>x"b800", 440=>x"c000", 441=>x"c200",
--442=>x"c200", 443=>x"c100", 444=>x"b100", 445=>x"ba00", 446=>x"be00", 447=>x"c200", 448=>x"c100",
--449=>x"be00", 450=>x"b500", 451=>x"ac00", 452=>x"b700", 453=>x"c400", 454=>x"ca00", 455=>x"c200",
--456=>x"af00", 457=>x"a700", 458=>x"b200", 459=>x"bc00", 460=>x"c200", 461=>x"c300", 462=>x"c500",
--463=>x"c800", 464=>x"a800", 465=>x"b800", 466=>x"ba00", 467=>x"bf00", 468=>x"bc00", 469=>x"c200",
--470=>x"c200", 471=>x"3b00", 472=>x"c100", 473=>x"be00", 474=>x"bc00", 475=>x"b700", 476=>x"bd00",
--477=>x"c300", 478=>x"c600", 479=>x"c100", 480=>x"bd00", 481=>x"b600", 482=>x"b900", 483=>x"bc00",
--484=>x"b700", 485=>x"c000", 486=>x"c400", 487=>x"bf00", 488=>x"b600", 489=>x"bc00", 490=>x"bf00",
--491=>x"bc00", 492=>x"bf00", 493=>x"bf00", 494=>x"c200", 495=>x"bb00", 496=>x"bc00", 497=>x"bf00",
--498=>x"c200", 499=>x"bd00"),
--16 => (0=>x"8c00", 1=>x"8800", 2=>x"8200", 3=>x"8000", 4=>x"8400", 5=>x"8200", 6=>x"8500", 7=>x"8300",
--8=>x"8c00", 9=>x"8600", 10=>x"8200", 11=>x"8000", 12=>x"8500", 13=>x"8200", 14=>x"8500",
--15=>x"8300", 16=>x"8a00", 17=>x"8800", 18=>x"8300", 19=>x"7f00", 20=>x"8300", 21=>x"8400",
--22=>x"8300", 23=>x"8200", 24=>x"8300", 25=>x"8600", 26=>x"8400", 27=>x"8000", 28=>x"8000",
--29=>x"7f00", 30=>x"7e00", 31=>x"8300", 32=>x"8300", 33=>x"8500", 34=>x"8200", 35=>x"8200",
--36=>x"8000", 37=>x"7f00", 38=>x"8100", 39=>x"8000", 40=>x"8100", 41=>x"8300", 42=>x"8200",
--43=>x"8400", 44=>x"8200", 45=>x"8100", 46=>x"7e00", 47=>x"7f00", 48=>x"8100", 49=>x"8200",
--50=>x"8200", 51=>x"8300", 52=>x"8300", 53=>x"8400", 54=>x"8100", 55=>x"8100", 56=>x"8100",
--57=>x"8300", 58=>x"8200", 59=>x"8200", 60=>x"8100", 61=>x"8200", 62=>x"8200", 63=>x"7f00",
--64=>x"8200", 65=>x"8100", 66=>x"8300", 67=>x"8200", 68=>x"8300", 69=>x"8300", 70=>x"8200",
--71=>x"7e00", 72=>x"8300", 73=>x"8300", 74=>x"8300", 75=>x"8400", 76=>x"8600", 77=>x"8100",
--78=>x"8100", 79=>x"7f00", 80=>x"8400", 81=>x"8300", 82=>x"8200", 83=>x"8000", 84=>x"8900",
--85=>x"8000", 86=>x"8100", 87=>x"7e00", 88=>x"8200", 89=>x"8200", 90=>x"8200", 91=>x"8100",
--92=>x"8200", 93=>x"8200", 94=>x"8100", 95=>x"8100", 96=>x"8100", 97=>x"8100", 98=>x"8300",
--99=>x"8300", 100=>x"8100", 101=>x"8200", 102=>x"8000", 103=>x"7f00", 104=>x"8300", 105=>x"8400",
--106=>x"8300", 107=>x"8400", 108=>x"7f00", 109=>x"7f00", 110=>x"7f00", 111=>x"7e00", 112=>x"8200",
--113=>x"8400", 114=>x"8500", 115=>x"8400", 116=>x"8100", 117=>x"7e00", 118=>x"7f00", 119=>x"7f00",
--120=>x"8500", 121=>x"8100", 122=>x"8400", 123=>x"8200", 124=>x"7f00", 125=>x"7d00", 126=>x"8000",
--127=>x"7f00", 128=>x"8500", 129=>x"8300", 130=>x"8300", 131=>x"8100", 132=>x"8000", 133=>x"7d00",
--134=>x"7e00", 135=>x"7e00", 136=>x"8300", 137=>x"8500", 138=>x"8300", 139=>x"8100", 140=>x"7f00",
--141=>x"8100", 142=>x"8000", 143=>x"8000", 144=>x"8300", 145=>x"8400", 146=>x"8400", 147=>x"8000",
--148=>x"7f00", 149=>x"8000", 150=>x"8100", 151=>x"8000", 152=>x"8600", 153=>x"8200", 154=>x"8200",
--155=>x"8200", 156=>x"7e00", 157=>x"8100", 158=>x"7f00", 159=>x"7f00", 160=>x"8300", 161=>x"8200",
--162=>x"7f00", 163=>x"7e00", 164=>x"7d00", 165=>x"8100", 166=>x"7f00", 167=>x"7c00", 168=>x"8000",
--169=>x"8400", 170=>x"8000", 171=>x"8000", 172=>x"8300", 173=>x"8000", 174=>x"7e00", 175=>x"7f00",
--176=>x"7c00", 177=>x"7d00", 178=>x"7c00", 179=>x"7e00", 180=>x"7f00", 181=>x"7f00", 182=>x"7e00",
--183=>x"8000", 184=>x"7800", 185=>x"7d00", 186=>x"7b00", 187=>x"7c00", 188=>x"7d00", 189=>x"7d00",
--190=>x"7c00", 191=>x"7f00", 192=>x"7600", 193=>x"7800", 194=>x"7a00", 195=>x"7c00", 196=>x"7c00",
--197=>x"7c00", 198=>x"7d00", 199=>x"7d00", 200=>x"7400", 201=>x"7100", 202=>x"7100", 203=>x"7900",
--204=>x"7900", 205=>x"7a00", 206=>x"7c00", 207=>x"7a00", 208=>x"a700", 209=>x"8f00", 210=>x"7700",
--211=>x"6f00", 212=>x"7500", 213=>x"7600", 214=>x"7900", 215=>x"7800", 216=>x"c400", 217=>x"c000",
--218=>x"b100", 219=>x"8900", 220=>x"7200", 221=>x"7000", 222=>x"7700", 223=>x"7800", 224=>x"c200",
--225=>x"c600", 226=>x"c800", 227=>x"c200", 228=>x"a500", 229=>x"7c00", 230=>x"6f00", 231=>x"7300",
--232=>x"c100", 233=>x"c400", 234=>x"c200", 235=>x"c500", 236=>x"c600", 237=>x"bb00", 238=>x"8e00",
--239=>x"9100", 240=>x"c100", 241=>x"c400", 242=>x"c000", 243=>x"c100", 244=>x"c300", 245=>x"cb00",
--246=>x"c400", 247=>x"a200", 248=>x"bc00", 249=>x"c200", 250=>x"c200", 251=>x"c100", 252=>x"c600",
--253=>x"c500", 254=>x"ca00", 255=>x"c800", 256=>x"bd00", 257=>x"bb00", 258=>x"bf00", 259=>x"c100",
--260=>x"c500", 261=>x"c400", 262=>x"c400", 263=>x"c200", 264=>x"b800", 265=>x"bf00", 266=>x"c200",
--267=>x"c100", 268=>x"c500", 269=>x"c300", 270=>x"c400", 271=>x"c500", 272=>x"bd00", 273=>x"bd00",
--274=>x"c000", 275=>x"c300", 276=>x"c400", 277=>x"c300", 278=>x"c700", 279=>x"c500", 280=>x"c100",
--281=>x"be00", 282=>x"bd00", 283=>x"c300", 284=>x"c300", 285=>x"c600", 286=>x"c500", 287=>x"c400",
--288=>x"bf00", 289=>x"bf00", 290=>x"c400", 291=>x"c300", 292=>x"c400", 293=>x"c400", 294=>x"c400",
--295=>x"c400", 296=>x"c100", 297=>x"3d00", 298=>x"c100", 299=>x"c700", 300=>x"c400", 301=>x"c400",
--302=>x"c400", 303=>x"c000", 304=>x"be00", 305=>x"c100", 306=>x"c400", 307=>x"c500", 308=>x"c300",
--309=>x"c300", 310=>x"c500", 311=>x"c000", 312=>x"c400", 313=>x"b900", 314=>x"c300", 315=>x"c500",
--316=>x"c300", 317=>x"c000", 318=>x"c000", 319=>x"bc00", 320=>x"c000", 321=>x"c000", 322=>x"c400",
--323=>x"bc00", 324=>x"ba00", 325=>x"b900", 326=>x"b900", 327=>x"b900", 328=>x"c100", 329=>x"bc00",
--330=>x"b000", 331=>x"b100", 332=>x"b800", 333=>x"bc00", 334=>x"cb00", 335=>x"d300", 336=>x"ab00",
--337=>x"ab00", 338=>x"b100", 339=>x"be00", 340=>x"ce00", 341=>x"d400", 342=>x"d300", 343=>x"d500",
--344=>x"b400", 345=>x"c500", 346=>x"cf00", 347=>x"d700", 348=>x"d500", 349=>x"d200", 350=>x"cd00",
--351=>x"cd00", 352=>x"d100", 353=>x"d500", 354=>x"d500", 355=>x"d500", 356=>x"d200", 357=>x"ce00",
--358=>x"c800", 359=>x"3500", 360=>x"d200", 361=>x"d600", 362=>x"ce00", 363=>x"cb00", 364=>x"cb00",
--365=>x"cd00", 366=>x"d000", 367=>x"c900", 368=>x"ca00", 369=>x"cb00", 370=>x"c900", 371=>x"ce00",
--372=>x"d500", 373=>x"d000", 374=>x"cd00", 375=>x"cb00", 376=>x"c800", 377=>x"c900", 378=>x"cf00",
--379=>x"d700", 380=>x"d000", 381=>x"d000", 382=>x"cc00", 383=>x"c900", 384=>x"c900", 385=>x"d200",
--386=>x"ca00", 387=>x"ce00", 388=>x"cc00", 389=>x"c500", 390=>x"c500", 391=>x"c400", 392=>x"cb00",
--393=>x"c600", 394=>x"ca00", 395=>x"c700", 396=>x"c300", 397=>x"c200", 398=>x"c300", 399=>x"c700",
--400=>x"ca00", 401=>x"c300", 402=>x"3a00", 403=>x"ca00", 404=>x"c400", 405=>x"cb00", 406=>x"c600",
--407=>x"c200", 408=>x"c500", 409=>x"3a00", 410=>x"c600", 411=>x"c900", 412=>x"ca00", 413=>x"c000",
--414=>x"c400", 415=>x"c500", 416=>x"c300", 417=>x"c600", 418=>x"3b00", 419=>x"c100", 420=>x"c400",
--421=>x"c800", 422=>x"cc00", 423=>x"cb00", 424=>x"b700", 425=>x"bc00", 426=>x"bc00", 427=>x"c400",
--428=>x"cc00", 429=>x"cd00", 430=>x"ce00", 431=>x"cc00", 432=>x"b700", 433=>x"c100", 434=>x"c900",
--435=>x"3800", 436=>x"c900", 437=>x"cd00", 438=>x"cc00", 439=>x"ce00", 440=>x"c700", 441=>x"c300",
--442=>x"c400", 443=>x"ca00", 444=>x"c500", 445=>x"c900", 446=>x"cc00", 447=>x"cb00", 448=>x"c400",
--449=>x"c500", 450=>x"c000", 451=>x"c200", 452=>x"c700", 453=>x"c600", 454=>x"cd00", 455=>x"ce00",
--456=>x"c200", 457=>x"c500", 458=>x"ca00", 459=>x"c100", 460=>x"c300", 461=>x"cc00", 462=>x"c700",
--463=>x"3100", 464=>x"c900", 465=>x"c200", 466=>x"c500", 467=>x"c700", 468=>x"c400", 469=>x"c600",
--470=>x"c500", 471=>x"c400", 472=>x"c400", 473=>x"c400", 474=>x"bd00", 475=>x"c800", 476=>x"c400",
--477=>x"c000", 478=>x"c600", 479=>x"c600", 480=>x"c300", 481=>x"c400", 482=>x"c400", 483=>x"4200",
--484=>x"c400", 485=>x"c100", 486=>x"c000", 487=>x"c200", 488=>x"bf00", 489=>x"c500", 490=>x"c200",
--491=>x"c300", 492=>x"be00", 493=>x"be00", 494=>x"bb00", 495=>x"b700", 496=>x"ba00", 497=>x"c000",
--498=>x"c600", 499=>x"c200"),
--17 => (0=>x"8000", 1=>x"8200", 2=>x"8100", 3=>x"8600", 4=>x"8200", 5=>x"7f00", 6=>x"8200", 7=>x"8300",
--8=>x"8000", 9=>x"8200", 10=>x"8100", 11=>x"8600", 12=>x"8200", 13=>x"7f00", 14=>x"8200",
--15=>x"8300", 16=>x"8000", 17=>x"8200", 18=>x"8000", 19=>x"8600", 20=>x"8100", 21=>x"7e00",
--22=>x"8100", 23=>x"8200", 24=>x"7f00", 25=>x"8000", 26=>x"8000", 27=>x"8000", 28=>x"7e00",
--29=>x"7e00", 30=>x"8100", 31=>x"8300", 32=>x"7f00", 33=>x"7f00", 34=>x"7f00", 35=>x"8000",
--36=>x"7d00", 37=>x"7e00", 38=>x"7f00", 39=>x"7f00", 40=>x"8000", 41=>x"8000", 42=>x"8000",
--43=>x"8000", 44=>x"7f00", 45=>x"8000", 46=>x"7e00", 47=>x"7f00", 48=>x"8000", 49=>x"8100",
--50=>x"8200", 51=>x"8100", 52=>x"7f00", 53=>x"8100", 54=>x"8000", 55=>x"8200", 56=>x"8000",
--57=>x"8100", 58=>x"7f00", 59=>x"7f00", 60=>x"8000", 61=>x"7f00", 62=>x"7f00", 63=>x"8100",
--64=>x"8200", 65=>x"8100", 66=>x"7f00", 67=>x"7f00", 68=>x"7f00", 69=>x"7b00", 70=>x"8000",
--71=>x"8100", 72=>x"7f00", 73=>x"8300", 74=>x"8200", 75=>x"8200", 76=>x"8100", 77=>x"7e00",
--78=>x"7f00", 79=>x"7e00", 80=>x"8100", 81=>x"8000", 82=>x"8000", 83=>x"8200", 84=>x"8300",
--85=>x"7e00", 86=>x"7d00", 87=>x"7f00", 88=>x"8000", 89=>x"8200", 90=>x"7e00", 91=>x"7c00",
--92=>x"7d00", 93=>x"7f00", 94=>x"7d00", 95=>x"8000", 96=>x"7f00", 97=>x"8200", 98=>x"8000",
--99=>x"7f00", 100=>x"7e00", 101=>x"7d00", 102=>x"7c00", 103=>x"7e00", 104=>x"7d00", 105=>x"7f00",
--106=>x"8000", 107=>x"7e00", 108=>x"8000", 109=>x"7e00", 110=>x"7e00", 111=>x"7f00", 112=>x"8000",
--113=>x"8000", 114=>x"8000", 115=>x"8000", 116=>x"7d00", 117=>x"7f00", 118=>x"7f00", 119=>x"7d00",
--120=>x"7d00", 121=>x"8200", 122=>x"7f00", 123=>x"8000", 124=>x"8100", 125=>x"7e00", 126=>x"7c00",
--127=>x"7f00", 128=>x"7c00", 129=>x"8200", 130=>x"8000", 131=>x"7d00", 132=>x"8000", 133=>x"7e00",
--134=>x"7c00", 135=>x"7f00", 136=>x"8000", 137=>x"8300", 138=>x"7e00", 139=>x"7e00", 140=>x"8100",
--141=>x"7d00", 142=>x"7d00", 143=>x"7e00", 144=>x"8000", 145=>x"7f00", 146=>x"8000", 147=>x"7e00",
--148=>x"7e00", 149=>x"7e00", 150=>x"7c00", 151=>x"7d00", 152=>x"8000", 153=>x"8200", 154=>x"8100",
--155=>x"7f00", 156=>x"7e00", 157=>x"8000", 158=>x"7e00", 159=>x"7d00", 160=>x"7f00", 161=>x"8000",
--162=>x"7f00", 163=>x"7f00", 164=>x"7e00", 165=>x"7d00", 166=>x"7e00", 167=>x"7f00", 168=>x"7b00",
--169=>x"7e00", 170=>x"8200", 171=>x"7a00", 172=>x"7f00", 173=>x"7c00", 174=>x"8200", 175=>x"8200",
--176=>x"7e00", 177=>x"8100", 178=>x"8100", 179=>x"8200", 180=>x"8200", 181=>x"7e00", 182=>x"8000",
--183=>x"8000", 184=>x"7f00", 185=>x"8100", 186=>x"8200", 187=>x"8100", 188=>x"8300", 189=>x"7f00",
--190=>x"8000", 191=>x"7d00", 192=>x"7f00", 193=>x"8200", 194=>x"8200", 195=>x"8100", 196=>x"8300",
--197=>x"8300", 198=>x"8200", 199=>x"7d00", 200=>x"7e00", 201=>x"8200", 202=>x"8300", 203=>x"8200",
--204=>x"8100", 205=>x"8100", 206=>x"8000", 207=>x"7d00", 208=>x"7d00", 209=>x"7d00", 210=>x"7f00",
--211=>x"7f00", 212=>x"7d00", 213=>x"7f00", 214=>x"7f00", 215=>x"7e00", 216=>x"7800", 217=>x"7b00",
--218=>x"7c00", 219=>x"7e00", 220=>x"7d00", 221=>x"7f00", 222=>x"7f00", 223=>x"8100", 224=>x"7500",
--225=>x"7600", 226=>x"7e00", 227=>x"7c00", 228=>x"7e00", 229=>x"8100", 230=>x"7f00", 231=>x"7e00",
--232=>x"6c00", 233=>x"7600", 234=>x"7c00", 235=>x"7900", 236=>x"7a00", 237=>x"7d00", 238=>x"8000",
--239=>x"7b00", 240=>x"7800", 241=>x"6c00", 242=>x"8800", 243=>x"7300", 244=>x"7600", 245=>x"7500",
--246=>x"7700", 247=>x"7900", 248=>x"b800", 249=>x"8f00", 250=>x"7000", 251=>x"6d00", 252=>x"7100",
--253=>x"7100", 254=>x"7600", 255=>x"7800", 256=>x"c900", 257=>x"c400", 258=>x"9f00", 259=>x"7400",
--260=>x"6a00", 261=>x"6d00", 262=>x"7200", 263=>x"7200", 264=>x"c300", 265=>x"c100", 266=>x"c500",
--267=>x"b500", 268=>x"8500", 269=>x"9700", 270=>x"6700", 271=>x"6b00", 272=>x"c100", 273=>x"c300",
--274=>x"c200", 275=>x"c900", 276=>x"c300", 277=>x"9e00", 278=>x"6c00", 279=>x"6300", 280=>x"c300",
--281=>x"c500", 282=>x"c600", 283=>x"c900", 284=>x"cc00", 285=>x"ca00", 286=>x"ab00", 287=>x"7200",
--288=>x"c300", 289=>x"c300", 290=>x"c500", 291=>x"ca00", 292=>x"ca00", 293=>x"ca00", 294=>x"d000",
--295=>x"b100", 296=>x"c300", 297=>x"c600", 298=>x"c800", 299=>x"c600", 300=>x"c400", 301=>x"c100",
--302=>x"c400", 303=>x"cc00", 304=>x"c100", 305=>x"c100", 306=>x"bc00", 307=>x"b800", 308=>x"bc00",
--309=>x"c100", 310=>x"cb00", 311=>x"d500", 312=>x"b800", 313=>x"bc00", 314=>x"be00", 315=>x"cb00",
--316=>x"d300", 317=>x"d700", 318=>x"d900", 319=>x"db00", 320=>x"c500", 321=>x"d100", 322=>x"d400",
--323=>x"d400", 324=>x"d800", 325=>x"d600", 326=>x"d500", 327=>x"d700", 328=>x"d800", 329=>x"d300",
--330=>x"d300", 331=>x"d200", 332=>x"d200", 333=>x"d600", 334=>x"d200", 335=>x"d300", 336=>x"d300",
--337=>x"cf00", 338=>x"cf00", 339=>x"d300", 340=>x"d000", 341=>x"d200", 342=>x"d300", 343=>x"ce00",
--344=>x"ce00", 345=>x"d000", 346=>x"d100", 347=>x"cf00", 348=>x"cf00", 349=>x"cd00", 350=>x"d200",
--351=>x"d500", 352=>x"d000", 353=>x"ce00", 354=>x"cf00", 355=>x"d000", 356=>x"3200", 357=>x"cf00",
--358=>x"cf00", 359=>x"d200", 360=>x"ce00", 361=>x"d100", 362=>x"ce00", 363=>x"cf00", 364=>x"ce00",
--365=>x"cb00", 366=>x"cf00", 367=>x"3200", 368=>x"c900", 369=>x"cf00", 370=>x"ce00", 371=>x"cb00",
--372=>x"cc00", 373=>x"ca00", 374=>x"ca00", 375=>x"cf00", 376=>x"c500", 377=>x"c100", 378=>x"c400",
--379=>x"cb00", 380=>x"ca00", 381=>x"ce00", 382=>x"d600", 383=>x"d900", 384=>x"ca00", 385=>x"c700",
--386=>x"c700", 387=>x"cf00", 388=>x"d100", 389=>x"cb00", 390=>x"cf00", 391=>x"ce00", 392=>x"2e00",
--393=>x"d100", 394=>x"c900", 395=>x"c700", 396=>x"c800", 397=>x"c500", 398=>x"c700", 399=>x"c800",
--400=>x"c700", 401=>x"c800", 402=>x"c900", 403=>x"ca00", 404=>x"c900", 405=>x"cb00", 406=>x"d000",
--407=>x"cd00", 408=>x"cd00", 409=>x"c400", 410=>x"cb00", 411=>x"d300", 412=>x"cf00", 413=>x"ce00",
--414=>x"cd00", 415=>x"cf00", 416=>x"ce00", 417=>x"d100", 418=>x"c500", 419=>x"cd00", 420=>x"d200",
--421=>x"cf00", 422=>x"cf00", 423=>x"cf00", 424=>x"c500", 425=>x"ce00", 426=>x"d100", 427=>x"c800",
--428=>x"ce00", 429=>x"cd00", 430=>x"d000", 431=>x"cc00", 432=>x"cd00", 433=>x"c800", 434=>x"d400",
--435=>x"ce00", 436=>x"c300", 437=>x"cf00", 438=>x"d000", 439=>x"cf00", 440=>x"cf00", 441=>x"ca00",
--442=>x"c900", 443=>x"d100", 444=>x"c800", 445=>x"cc00", 446=>x"cd00", 447=>x"cc00", 448=>x"cd00",
--449=>x"cc00", 450=>x"c600", 451=>x"3300", 452=>x"ce00", 453=>x"ca00", 454=>x"cd00", 455=>x"cf00",
--456=>x"cd00", 457=>x"ca00", 458=>x"c800", 459=>x"cc00", 460=>x"ca00", 461=>x"cc00", 462=>x"c700",
--463=>x"c600", 464=>x"ca00", 465=>x"ce00", 466=>x"c700", 467=>x"c500", 468=>x"c400", 469=>x"c100",
--470=>x"ca00", 471=>x"cb00", 472=>x"c700", 473=>x"c800", 474=>x"bf00", 475=>x"be00", 476=>x"c400",
--477=>x"c800", 478=>x"ce00", 479=>x"cf00", 480=>x"bf00", 481=>x"bb00", 482=>x"c200", 483=>x"cb00",
--484=>x"cc00", 485=>x"ca00", 486=>x"ca00", 487=>x"cd00", 488=>x"be00", 489=>x"c700", 490=>x"c900",
--491=>x"cb00", 492=>x"cc00", 493=>x"c800", 494=>x"ca00", 495=>x"cc00", 496=>x"c400", 497=>x"c900",
--498=>x"c800", 499=>x"c300"),
--18 => (0=>x"8000", 1=>x"8200", 2=>x"8100", 3=>x"8100", 4=>x"7f00", 5=>x"7f00", 6=>x"7f00", 7=>x"8000",
--8=>x"8000", 9=>x"8300", 10=>x"8000", 11=>x"8000", 12=>x"7f00", 13=>x"7f00", 14=>x"7f00",
--15=>x"8000", 16=>x"7f00", 17=>x"8100", 18=>x"8200", 19=>x"8000", 20=>x"8000", 21=>x"7f00",
--22=>x"8000", 23=>x"8000", 24=>x"7f00", 25=>x"8100", 26=>x"8200", 27=>x"7f00", 28=>x"8000",
--29=>x"8100", 30=>x"7e00", 31=>x"7c00", 32=>x"8000", 33=>x"8300", 34=>x"7f00", 35=>x"7f00",
--36=>x"8100", 37=>x"7e00", 38=>x"7d00", 39=>x"7e00", 40=>x"7d00", 41=>x"8000", 42=>x"8200",
--43=>x"7f00", 44=>x"8000", 45=>x"7e00", 46=>x"7f00", 47=>x"7f00", 48=>x"7f00", 49=>x"7c00",
--50=>x"8000", 51=>x"8100", 52=>x"7e00", 53=>x"7f00", 54=>x"8100", 55=>x"7f00", 56=>x"7f00",
--57=>x"7e00", 58=>x"8000", 59=>x"8300", 60=>x"7f00", 61=>x"8100", 62=>x"8200", 63=>x"7f00",
--64=>x"8100", 65=>x"8200", 66=>x"8000", 67=>x"8100", 68=>x"8000", 69=>x"8000", 70=>x"8100",
--71=>x"8200", 72=>x"8000", 73=>x"8200", 74=>x"8300", 75=>x"8100", 76=>x"8200", 77=>x"7d00",
--78=>x"7e00", 79=>x"8200", 80=>x"7f00", 81=>x"7e00", 82=>x"8300", 83=>x"8200", 84=>x"7e00",
--85=>x"7e00", 86=>x"8000", 87=>x"7f00", 88=>x"7f00", 89=>x"7c00", 90=>x"7f00", 91=>x"7f00",
--92=>x"7e00", 93=>x"7d00", 94=>x"8300", 95=>x"7f00", 96=>x"7e00", 97=>x"8000", 98=>x"7f00",
--99=>x"7d00", 100=>x"7d00", 101=>x"7b00", 102=>x"8000", 103=>x"8100", 104=>x"7f00", 105=>x"7f00",
--106=>x"7f00", 107=>x"7e00", 108=>x"7e00", 109=>x"8000", 110=>x"8000", 111=>x"7e00", 112=>x"7d00",
--113=>x"7e00", 114=>x"7e00", 115=>x"7e00", 116=>x"7c00", 117=>x"8000", 118=>x"8100", 119=>x"7d00",
--120=>x"7c00", 121=>x"7d00", 122=>x"7c00", 123=>x"7f00", 124=>x"7e00", 125=>x"7f00", 126=>x"8000",
--127=>x"8200", 128=>x"7f00", 129=>x"7d00", 130=>x"7e00", 131=>x"7e00", 132=>x"7f00", 133=>x"8000",
--134=>x"7f00", 135=>x"8000", 136=>x"8000", 137=>x"7f00", 138=>x"7b00", 139=>x"7d00", 140=>x"8000",
--141=>x"7f00", 142=>x"8000", 143=>x"7f00", 144=>x"7a00", 145=>x"7f00", 146=>x"7f00", 147=>x"7d00",
--148=>x"7c00", 149=>x"7d00", 150=>x"7e00", 151=>x"7e00", 152=>x"7d00", 153=>x"7c00", 154=>x"7e00",
--155=>x"7d00", 156=>x"8000", 157=>x"7d00", 158=>x"7d00", 159=>x"7f00", 160=>x"8000", 161=>x"7e00",
--162=>x"7d00", 163=>x"7f00", 164=>x"7d00", 165=>x"7c00", 166=>x"8000", 167=>x"7e00", 168=>x"7c00",
--169=>x"7f00", 170=>x"7d00", 171=>x"7e00", 172=>x"7e00", 173=>x"7e00", 174=>x"8000", 175=>x"7e00",
--176=>x"7e00", 177=>x"8000", 178=>x"8200", 179=>x"7f00", 180=>x"7f00", 181=>x"7d00", 182=>x"7e00",
--183=>x"8000", 184=>x"7d00", 185=>x"7e00", 186=>x"8100", 187=>x"7e00", 188=>x"7f00", 189=>x"8000",
--190=>x"8100", 191=>x"7f00", 192=>x"8000", 193=>x"7d00", 194=>x"7e00", 195=>x"7f00", 196=>x"7e00",
--197=>x"8000", 198=>x"7d00", 199=>x"7d00", 200=>x"8000", 201=>x"7e00", 202=>x"7c00", 203=>x"8100",
--204=>x"7f00", 205=>x"7d00", 206=>x"8000", 207=>x"7c00", 208=>x"7e00", 209=>x"8000", 210=>x"7d00",
--211=>x"8000", 212=>x"7c00", 213=>x"7c00", 214=>x"7d00", 215=>x"7e00", 216=>x"7e00", 217=>x"7e00",
--218=>x"7a00", 219=>x"7e00", 220=>x"7e00", 221=>x"7b00", 222=>x"7b00", 223=>x"7a00", 224=>x"7e00",
--225=>x"7b00", 226=>x"7d00", 227=>x"8000", 228=>x"7c00", 229=>x"7a00", 230=>x"7b00", 231=>x"7900",
--232=>x"7800", 233=>x"7900", 234=>x"7e00", 235=>x"7d00", 236=>x"7900", 237=>x"7d00", 238=>x"7b00",
--239=>x"7a00", 240=>x"7900", 241=>x"7900", 242=>x"7700", 243=>x"7a00", 244=>x"7600", 245=>x"7900",
--246=>x"7a00", 247=>x"7800", 248=>x"7700", 249=>x"7600", 250=>x"7a00", 251=>x"7900", 252=>x"7800",
--253=>x"7600", 254=>x"7700", 255=>x"7800", 256=>x"7400", 257=>x"7700", 258=>x"7800", 259=>x"7800",
--260=>x"7700", 261=>x"7800", 262=>x"7700", 263=>x"7700", 264=>x"6e00", 265=>x"7500", 266=>x"7400",
--267=>x"7100", 268=>x"7300", 269=>x"7300", 270=>x"7300", 271=>x"7700", 272=>x"6c00", 273=>x"6c00",
--274=>x"6a00", 275=>x"6c00", 276=>x"6e00", 277=>x"7100", 278=>x"7100", 279=>x"7300", 280=>x"6200",
--281=>x"6500", 282=>x"6800", 283=>x"6900", 284=>x"6a00", 285=>x"6c00", 286=>x"6e00", 287=>x"7200",
--288=>x"7500", 289=>x"5900", 290=>x"5d00", 291=>x"6000", 292=>x"6400", 293=>x"6700", 294=>x"6b00",
--295=>x"6c00", 296=>x"bb00", 297=>x"7b00", 298=>x"7200", 299=>x"6400", 300=>x"a700", 301=>x"6100",
--302=>x"6300", 303=>x"6900", 304=>x"da00", 305=>x"d500", 306=>x"cf00", 307=>x"b900", 308=>x"7600",
--309=>x"5500", 310=>x"5e00", 311=>x"6500", 312=>x"dc00", 313=>x"e400", 314=>x"e600", 315=>x"e900",
--316=>x"c400", 317=>x"6500", 318=>x"5500", 319=>x"5a00", 320=>x"d600", 321=>x"da00", 322=>x"e100",
--323=>x"e300", 324=>x"e600", 325=>x"9d00", 326=>x"4e00", 327=>x"5200", 328=>x"d800", 329=>x"d700",
--330=>x"dd00", 331=>x"e200", 332=>x"e300", 333=>x"d000", 334=>x"7700", 335=>x"4b00", 336=>x"d000",
--337=>x"d600", 338=>x"d800", 339=>x"df00", 340=>x"e000", 341=>x"e300", 342=>x"c400", 343=>x"6000",
--344=>x"cd00", 345=>x"d000", 346=>x"d800", 347=>x"da00", 348=>x"e000", 349=>x"de00", 350=>x"e200",
--351=>x"a500", 352=>x"d300", 353=>x"ce00", 354=>x"d000", 355=>x"d400", 356=>x"d500", 357=>x"df00",
--358=>x"df00", 359=>x"da00", 360=>x"cd00", 361=>x"d200", 362=>x"d200", 363=>x"d600", 364=>x"d500",
--365=>x"de00", 366=>x"e100", 367=>x"de00", 368=>x"d100", 369=>x"d400", 370=>x"2600", 371=>x"d900",
--372=>x"da00", 373=>x"df00", 374=>x"e500", 375=>x"e000", 376=>x"d700", 377=>x"d200", 378=>x"d500",
--379=>x"d200", 380=>x"d400", 381=>x"d800", 382=>x"dc00", 383=>x"e100", 384=>x"cb00", 385=>x"ca00",
--386=>x"cc00", 387=>x"ce00", 388=>x"ce00", 389=>x"d100", 390=>x"d400", 391=>x"d600", 392=>x"c700",
--393=>x"ce00", 394=>x"d100", 395=>x"d100", 396=>x"d400", 397=>x"d300", 398=>x"d400", 399=>x"d400",
--400=>x"ce00", 401=>x"cf00", 402=>x"d100", 403=>x"d300", 404=>x"d000", 405=>x"d300", 406=>x"d200",
--407=>x"d400", 408=>x"d000", 409=>x"d000", 410=>x"ce00", 411=>x"d200", 412=>x"d100", 413=>x"d100",
--414=>x"d400", 415=>x"ce00", 416=>x"cf00", 417=>x"d000", 418=>x"cd00", 419=>x"cb00", 420=>x"cf00",
--421=>x"d000", 422=>x"d100", 423=>x"cc00", 424=>x"ce00", 425=>x"d100", 426=>x"cf00", 427=>x"ce00",
--428=>x"d200", 429=>x"d100", 430=>x"d300", 431=>x"d100", 432=>x"ce00", 433=>x"d200", 434=>x"cf00",
--435=>x"cf00", 436=>x"cf00", 437=>x"cc00", 438=>x"ca00", 439=>x"cd00", 440=>x"cd00", 441=>x"cb00",
--442=>x"cc00", 443=>x"cb00", 444=>x"ca00", 445=>x"cd00", 446=>x"cb00", 447=>x"cd00", 448=>x"cb00",
--449=>x"c300", 450=>x"c400", 451=>x"c900", 452=>x"ca00", 453=>x"d100", 454=>x"d400", 455=>x"d100",
--456=>x"c800", 457=>x"cb00", 458=>x"c800", 459=>x"cb00", 460=>x"ce00", 461=>x"cf00", 462=>x"d000",
--463=>x"d400", 464=>x"cb00", 465=>x"d400", 466=>x"cd00", 467=>x"c400", 468=>x"ca00", 469=>x"ce00",
--470=>x"cf00", 471=>x"d000", 472=>x"cc00", 473=>x"ca00", 474=>x"d200", 475=>x"cd00", 476=>x"c800",
--477=>x"cb00", 478=>x"ce00", 479=>x"cf00", 480=>x"ce00", 481=>x"c900", 482=>x"c900", 483=>x"cd00",
--484=>x"cf00", 485=>x"c700", 486=>x"ca00", 487=>x"d000", 488=>x"cb00", 489=>x"c800", 490=>x"c600",
--491=>x"c300", 492=>x"c900", 493=>x"c700", 494=>x"c400", 495=>x"3300", 496=>x"c500", 497=>x"c600",
--498=>x"ca00", 499=>x"c700"),
--19 => (0=>x"7d00", 1=>x"7c00", 2=>x"7800", 3=>x"7a00", 4=>x"7500", 5=>x"7100", 6=>x"7000", 7=>x"6600",
--8=>x"8300", 9=>x"7b00", 10=>x"7800", 11=>x"7900", 12=>x"7600", 13=>x"7100", 14=>x"7000",
--15=>x"6600", 16=>x"7a00", 17=>x"7a00", 18=>x"7a00", 19=>x"7800", 20=>x"7300", 21=>x"7200",
--22=>x"6f00", 23=>x"6600", 24=>x"7c00", 25=>x"7900", 26=>x"7b00", 27=>x"7800", 28=>x"7300",
--29=>x"7100", 30=>x"6c00", 31=>x"6700", 32=>x"7c00", 33=>x"7c00", 34=>x"7800", 35=>x"7700",
--36=>x"7400", 37=>x"7000", 38=>x"6f00", 39=>x"6d00", 40=>x"7c00", 41=>x"7b00", 42=>x"7600",
--43=>x"7700", 44=>x"7500", 45=>x"7200", 46=>x"6f00", 47=>x"6b00", 48=>x"7c00", 49=>x"7b00",
--50=>x"7a00", 51=>x"7a00", 52=>x"7500", 53=>x"7100", 54=>x"6f00", 55=>x"6e00", 56=>x"7b00",
--57=>x"8300", 58=>x"7c00", 59=>x"7900", 60=>x"7600", 61=>x"7200", 62=>x"6e00", 63=>x"7300",
--64=>x"8000", 65=>x"7c00", 66=>x"7900", 67=>x"7900", 68=>x"7600", 69=>x"7500", 70=>x"7200",
--71=>x"7700", 72=>x"7e00", 73=>x"7d00", 74=>x"7d00", 75=>x"7a00", 76=>x"7400", 77=>x"7200",
--78=>x"7100", 79=>x"7200", 80=>x"7e00", 81=>x"7c00", 82=>x"7b00", 83=>x"7b00", 84=>x"8000",
--85=>x"7900", 86=>x"7100", 87=>x"7100", 88=>x"7e00", 89=>x"7b00", 90=>x"7b00", 91=>x"7a00",
--92=>x"7900", 93=>x"7800", 94=>x"7200", 95=>x"7100", 96=>x"7d00", 97=>x"7c00", 98=>x"7e00",
--99=>x"7900", 100=>x"7900", 101=>x"7800", 102=>x"7300", 103=>x"6e00", 104=>x"7e00", 105=>x"7c00",
--106=>x"7a00", 107=>x"7a00", 108=>x"7e00", 109=>x"7d00", 110=>x"7400", 111=>x"6e00", 112=>x"7d00",
--113=>x"7b00", 114=>x"7b00", 115=>x"7900", 116=>x"7900", 117=>x"7900", 118=>x"7700", 119=>x"7100",
--120=>x"8000", 121=>x"8100", 122=>x"7d00", 123=>x"7700", 124=>x"7400", 125=>x"7700", 126=>x"7600",
--127=>x"7400", 128=>x"7c00", 129=>x"8000", 130=>x"7c00", 131=>x"7900", 132=>x"7700", 133=>x"7800",
--134=>x"7300", 135=>x"7000", 136=>x"7d00", 137=>x"7e00", 138=>x"7d00", 139=>x"7a00", 140=>x"7a00",
--141=>x"7700", 142=>x"7400", 143=>x"6f00", 144=>x"8000", 145=>x"7c00", 146=>x"7b00", 147=>x"7900",
--148=>x"7800", 149=>x"7500", 150=>x"7700", 151=>x"7400", 152=>x"8100", 153=>x"7d00", 154=>x"7c00",
--155=>x"7a00", 156=>x"7800", 157=>x"7500", 158=>x"7800", 159=>x"7900", 160=>x"7d00", 161=>x"7c00",
--162=>x"7c00", 163=>x"7800", 164=>x"7500", 165=>x"8c00", 166=>x"7400", 167=>x"7300", 168=>x"7d00",
--169=>x"7900", 170=>x"7a00", 171=>x"7a00", 172=>x"7500", 173=>x"7600", 174=>x"7300", 175=>x"7300",
--176=>x"7d00", 177=>x"7a00", 178=>x"7c00", 179=>x"7a00", 180=>x"7600", 181=>x"7700", 182=>x"6f00",
--183=>x"7300", 184=>x"7b00", 185=>x"7e00", 186=>x"7d00", 187=>x"7800", 188=>x"7500", 189=>x"7300",
--190=>x"7300", 191=>x"7100", 192=>x"8100", 193=>x"7d00", 194=>x"7a00", 195=>x"7700", 196=>x"7900",
--197=>x"7700", 198=>x"7200", 199=>x"7100", 200=>x"7d00", 201=>x"7c00", 202=>x"7900", 203=>x"7700",
--204=>x"7800", 205=>x"7800", 206=>x"7500", 207=>x"6f00", 208=>x"7c00", 209=>x"7600", 210=>x"7700",
--211=>x"7900", 212=>x"7500", 213=>x"7500", 214=>x"7600", 215=>x"7100", 216=>x"7b00", 217=>x"7800",
--218=>x"7900", 219=>x"7800", 220=>x"8a00", 221=>x"7000", 222=>x"7400", 223=>x"7000", 224=>x"7b00",
--225=>x"7700", 226=>x"7600", 227=>x"7500", 228=>x"7400", 229=>x"7100", 230=>x"7300", 231=>x"6f00",
--232=>x"7700", 233=>x"7400", 234=>x"7100", 235=>x"7300", 236=>x"7100", 237=>x"7000", 238=>x"7000",
--239=>x"6f00", 240=>x"7800", 241=>x"7500", 242=>x"7300", 243=>x"7400", 244=>x"7300", 245=>x"7200",
--246=>x"7000", 247=>x"6d00", 248=>x"7700", 249=>x"7600", 250=>x"7500", 251=>x"7300", 252=>x"7100",
--253=>x"7100", 254=>x"6d00", 255=>x"6b00", 256=>x"7500", 257=>x"7400", 258=>x"7500", 259=>x"7200",
--260=>x"8f00", 261=>x"7100", 262=>x"7000", 263=>x"6f00", 264=>x"7400", 265=>x"7500", 266=>x"7400",
--267=>x"7100", 268=>x"7100", 269=>x"6f00", 270=>x"6e00", 271=>x"6f00", 272=>x"7300", 273=>x"7200",
--274=>x"7200", 275=>x"7100", 276=>x"6d00", 277=>x"6d00", 278=>x"6e00", 279=>x"6a00", 280=>x"7200",
--281=>x"7100", 282=>x"8d00", 283=>x"6f00", 284=>x"6f00", 285=>x"6f00", 286=>x"6e00", 287=>x"6a00",
--288=>x"7200", 289=>x"6e00", 290=>x"7000", 291=>x"6f00", 292=>x"6c00", 293=>x"6a00", 294=>x"6a00",
--295=>x"6c00", 296=>x"6e00", 297=>x"6c00", 298=>x"6e00", 299=>x"6d00", 300=>x"6b00", 301=>x"6a00",
--302=>x"6b00", 303=>x"6900", 304=>x"6c00", 305=>x"6c00", 306=>x"6c00", 307=>x"6b00", 308=>x"6a00",
--309=>x"6800", 310=>x"6700", 311=>x"6800", 312=>x"6600", 313=>x"9700", 314=>x"9600", 315=>x"6a00",
--316=>x"6500", 317=>x"6400", 318=>x"6500", 319=>x"6800", 320=>x"5d00", 321=>x"6200", 322=>x"6700",
--323=>x"6500", 324=>x"6400", 325=>x"6600", 326=>x"6400", 327=>x"6600", 328=>x"5900", 329=>x"5b00",
--330=>x"6400", 331=>x"6500", 332=>x"6700", 333=>x"6500", 334=>x"6500", 335=>x"6400", 336=>x"b000",
--337=>x"5700", 338=>x"5c00", 339=>x"6000", 340=>x"6000", 341=>x"6400", 342=>x"6200", 343=>x"6100",
--344=>x"5400", 345=>x"4e00", 346=>x"5400", 347=>x"5c00", 348=>x"5d00", 349=>x"6300", 350=>x"6100",
--351=>x"6100", 352=>x"9a00", 353=>x"4f00", 354=>x"4e00", 355=>x"5400", 356=>x"5900", 357=>x"5e00",
--358=>x"6200", 359=>x"6000", 360=>x"d500", 361=>x"7900", 362=>x"4800", 363=>x"5100", 364=>x"5500",
--365=>x"5800", 366=>x"5900", 367=>x"5c00", 368=>x"de00", 369=>x"bf00", 370=>x"6100", 371=>x"4800",
--372=>x"5000", 373=>x"5100", 374=>x"5400", 375=>x"5700", 376=>x"df00", 377=>x"e400", 378=>x"a200",
--379=>x"4d00", 380=>x"4b00", 381=>x"4a00", 382=>x"5000", 383=>x"5300", 384=>x"d900", 385=>x"de00",
--386=>x"d300", 387=>x"9b00", 388=>x"6700", 389=>x"5000", 390=>x"4d00", 391=>x"4c00", 392=>x"d600",
--393=>x"da00", 394=>x"e000", 395=>x"e200", 396=>x"cb00", 397=>x"9000", 398=>x"4b00", 399=>x"4600",
--400=>x"d600", 401=>x"d900", 402=>x"da00", 403=>x"de00", 404=>x"e600", 405=>x"db00", 406=>x"9400",
--407=>x"5f00", 408=>x"d300", 409=>x"d600", 410=>x"d500", 411=>x"d500", 412=>x"da00", 413=>x"e200",
--414=>x"df00", 415=>x"9600", 416=>x"d200", 417=>x"d600", 418=>x"d300", 419=>x"d300", 420=>x"d400",
--421=>x"da00", 422=>x"e100", 423=>x"d600", 424=>x"cd00", 425=>x"d600", 426=>x"d900", 427=>x"d700",
--428=>x"d800", 429=>x"da00", 430=>x"d600", 431=>x"e000", 432=>x"c900", 433=>x"cf00", 434=>x"d300",
--435=>x"d700", 436=>x"d700", 437=>x"dd00", 438=>x"dc00", 439=>x"dd00", 440=>x"cc00", 441=>x"d000",
--442=>x"d400", 443=>x"d700", 444=>x"d800", 445=>x"d800", 446=>x"df00", 447=>x"e100", 448=>x"cd00",
--449=>x"ce00", 450=>x"d200", 451=>x"d400", 452=>x"d500", 453=>x"d300", 454=>x"d900", 455=>x"df00",
--456=>x"d000", 457=>x"ca00", 458=>x"cf00", 459=>x"d300", 460=>x"d100", 461=>x"d500", 462=>x"d700",
--463=>x"df00", 464=>x"d300", 465=>x"cb00", 466=>x"cd00", 467=>x"d400", 468=>x"d100", 469=>x"d200",
--470=>x"d600", 471=>x"d800", 472=>x"cf00", 473=>x"d100", 474=>x"d100", 475=>x"d000", 476=>x"d000",
--477=>x"d200", 478=>x"d200", 479=>x"d400", 480=>x"ce00", 481=>x"ce00", 482=>x"cf00", 483=>x"cd00",
--484=>x"ca00", 485=>x"cc00", 486=>x"cd00", 487=>x"d200", 488=>x"cf00", 489=>x"cc00", 490=>x"ca00",
--491=>x"cc00", 492=>x"cd00", 493=>x"cb00", 494=>x"d000", 495=>x"cf00", 496=>x"ce00", 497=>x"d000",
--498=>x"cb00", 499=>x"d000")
--);
--
--
---- 256x256 - 32 FDAs
---- constant c_PIXEL  : t_MATRIX := (
---- 0  => (0=>x"a200", 1=>x"a200", 2=>x"a000", 3=>x"a000", 4=>x"a300", 5=>x"a100", 6=>x"9f00", 7=>x"9f00",
---- 8=>x"a200", 9=>x"a200", 10=>x"a000", 11=>x"a000", 12=>x"a300", 13=>x"a100", 14=>x"9f00",
---- 15=>x"9f00", 16=>x"a300", 17=>x"a100", 18=>x"a000", 19=>x"a100", 20=>x"a200", 21=>x"9e00",
---- 22=>x"9e00", 23=>x"9d00", 24=>x"a200", 25=>x"9f00", 26=>x"9e00", 27=>x"9e00", 28=>x"9f00",
---- 29=>x"a000", 30=>x"9b00", 31=>x"9900", 32=>x"9c00", 33=>x"9d00", 34=>x"9e00", 35=>x"9d00",
---- 36=>x"9f00", 37=>x"9e00", 38=>x"9d00", 39=>x"9a00", 40=>x"9b00", 41=>x"9d00", 42=>x"9d00",
---- 43=>x"9700", 44=>x"9d00", 45=>x"9d00", 46=>x"9d00", 47=>x"9c00", 48=>x"9d00", 49=>x"9d00",
---- 50=>x"9d00", 51=>x"9a00", 52=>x"9d00", 53=>x"9d00", 54=>x"9b00", 55=>x"9c00", 56=>x"9e00",
---- 57=>x"9e00", 58=>x"9d00", 59=>x"9c00", 60=>x"6300", 61=>x"9b00", 62=>x"9c00", 63=>x"9b00",
---- 64=>x"9d00", 65=>x"6100", 66=>x"9c00", 67=>x"9a00", 68=>x"9c00", 69=>x"9d00", 70=>x"9c00",
---- 71=>x"9c00", 72=>x"9c00", 73=>x"9c00", 74=>x"9f00", 75=>x"9a00", 76=>x"9c00", 77=>x"9c00",
---- 78=>x"9c00", 79=>x"9e00", 80=>x"9b00", 81=>x"9c00", 82=>x"9d00", 83=>x"9c00", 84=>x"9b00",
---- 85=>x"9d00", 86=>x"9e00", 87=>x"9e00", 88=>x"9e00", 89=>x"9d00", 90=>x"9900", 91=>x"9c00",
---- 92=>x"9d00", 93=>x"9b00", 94=>x"9e00", 95=>x"9d00", 96=>x"9c00", 97=>x"9a00", 98=>x"9900",
---- 99=>x"9d00", 100=>x"9f00", 101=>x"9f00", 102=>x"9d00", 103=>x"9e00", 104=>x"9a00", 105=>x"9a00",
---- 106=>x"9900", 107=>x"9c00", 108=>x"9e00", 109=>x"9f00", 110=>x"9f00", 111=>x"9d00", 112=>x"9e00",
---- 113=>x"9e00", 114=>x"9d00", 115=>x"9d00", 116=>x"9d00", 117=>x"9f00", 118=>x"9f00", 119=>x"9d00",
---- 120=>x"9d00", 121=>x"6000", 122=>x"6000", 123=>x"9e00", 124=>x"9f00", 125=>x"6100", 126=>x"a100",
---- 127=>x"9f00", 128=>x"9d00", 129=>x"9f00", 130=>x"9f00", 131=>x"9c00", 132=>x"9d00", 133=>x"9e00",
---- 134=>x"a000", 135=>x"a000", 136=>x"9f00", 137=>x"9f00", 138=>x"9d00", 139=>x"9c00", 140=>x"9d00",
---- 141=>x"9e00", 142=>x"9f00", 143=>x"a100", 144=>x"a000", 145=>x"9d00", 146=>x"9e00", 147=>x"6000",
---- 148=>x"a100", 149=>x"a400", 150=>x"a300", 151=>x"a100", 152=>x"a100", 153=>x"a000", 154=>x"a100",
---- 155=>x"6100", 156=>x"a100", 157=>x"a300", 158=>x"a000", 159=>x"a100", 160=>x"a500", 161=>x"a200",
---- 162=>x"a200", 163=>x"a000", 164=>x"9f00", 165=>x"a200", 166=>x"a200", 167=>x"a100", 168=>x"a000",
---- 169=>x"a000", 170=>x"a200", 171=>x"a100", 172=>x"9f00", 173=>x"a100", 174=>x"a100", 175=>x"a400",
---- 176=>x"a100", 177=>x"9f00", 178=>x"a100", 179=>x"a200", 180=>x"a000", 181=>x"a000", 182=>x"a200",
---- 183=>x"a700", 184=>x"a300", 185=>x"a000", 186=>x"a200", 187=>x"a000", 188=>x"9e00", 189=>x"a100",
---- 190=>x"a300", 191=>x"5700", 192=>x"a300", 193=>x"a200", 194=>x"a200", 195=>x"a100", 196=>x"9f00",
---- 197=>x"a200", 198=>x"a600", 199=>x"a900", 200=>x"a200", 201=>x"a300", 202=>x"a000", 203=>x"a000",
---- 204=>x"9f00", 205=>x"a300", 206=>x"aa00", 207=>x"ac00", 208=>x"a100", 209=>x"9f00", 210=>x"9d00",
---- 211=>x"a100", 212=>x"a100", 213=>x"a600", 214=>x"aa00", 215=>x"aa00", 216=>x"a100", 217=>x"a200",
---- 218=>x"a000", 219=>x"a300", 220=>x"a600", 221=>x"a800", 222=>x"a900", 223=>x"a700", 224=>x"9e00",
---- 225=>x"a000", 226=>x"a000", 227=>x"a400", 228=>x"a800", 229=>x"ab00", 230=>x"a900", 231=>x"a500",
---- 232=>x"5f00", 233=>x"5f00", 234=>x"a200", 235=>x"a600", 236=>x"aa00", 237=>x"ad00", 238=>x"a700",
---- 239=>x"a100", 240=>x"a100", 241=>x"a200", 242=>x"a700", 243=>x"aa00", 244=>x"ac00", 245=>x"a800",
---- 246=>x"a400", 247=>x"9d00", 248=>x"a200", 249=>x"a300", 250=>x"a800", 251=>x"ab00", 252=>x"ab00",
---- 253=>x"a700", 254=>x"a000", 255=>x"9800", 256=>x"a500", 257=>x"a700", 258=>x"ac00", 259=>x"ae00",
---- 260=>x"a900", 261=>x"a300", 262=>x"9d00", 263=>x"9600", 264=>x"a700", 265=>x"ab00", 266=>x"b000",
---- 267=>x"ad00", 268=>x"a700", 269=>x"9f00", 270=>x"9900", 271=>x"9300", 272=>x"a900", 273=>x"ad00",
---- 274=>x"ae00", 275=>x"aa00", 276=>x"a300", 277=>x"9c00", 278=>x"9600", 279=>x"8b00", 280=>x"ad00",
---- 281=>x"ac00", 282=>x"ab00", 283=>x"a600", 284=>x"a000", 285=>x"9a00", 286=>x"9200", 287=>x"8300",
---- 288=>x"ad00", 289=>x"ab00", 290=>x"a900", 291=>x"a400", 292=>x"9e00", 293=>x"9400", 294=>x"8b00",
---- 295=>x"7e00", 296=>x"ad00", 297=>x"ad00", 298=>x"a700", 299=>x"9f00", 300=>x"9a00", 301=>x"8f00",
---- 302=>x"8000", 303=>x"7000", 304=>x"aa00", 305=>x"a700", 306=>x"a300", 307=>x"9e00", 308=>x"9500",
---- 309=>x"8a00", 310=>x"7700", 311=>x"6000", 312=>x"a700", 313=>x"a400", 314=>x"9f00", 315=>x"9900",
---- 316=>x"8f00", 317=>x"8100", 318=>x"6d00", 319=>x"5200", 320=>x"a200", 321=>x"a200", 322=>x"6600",
---- 323=>x"9300", 324=>x"8600", 325=>x"7600", 326=>x"6100", 327=>x"5100", 328=>x"a200", 329=>x"9f00",
---- 330=>x"9700", 331=>x"8c00", 332=>x"7b00", 333=>x"6a00", 334=>x"5500", 335=>x"5000", 336=>x"9b00",
---- 337=>x"9900", 338=>x"9200", 339=>x"8400", 340=>x"8e00", 341=>x"5e00", 342=>x"4f00", 343=>x"5200",
---- 344=>x"9700", 345=>x"9400", 346=>x"8900", 347=>x"7700", 348=>x"6200", 349=>x"5100", 350=>x"5300",
---- 351=>x"5600", 352=>x"9400", 353=>x"8d00", 354=>x"7e00", 355=>x"6a00", 356=>x"5700", 357=>x"5100",
---- 358=>x"5600", 359=>x"5900", 360=>x"8b00", 361=>x"7900", 362=>x"7300", 363=>x"5d00", 364=>x"5300",
---- 365=>x"5400", 366=>x"5800", 367=>x"5800", 368=>x"8300", 369=>x"7c00", 370=>x"6700", 371=>x"5500",
---- 372=>x"5400", 373=>x"5700", 374=>x"5d00", 375=>x"5900", 376=>x"7b00", 377=>x"6f00", 378=>x"5800",
---- 379=>x"5300", 380=>x"5500", 381=>x"5b00", 382=>x"6000", 383=>x"5c00", 384=>x"6d00", 385=>x"6100",
---- 386=>x"5100", 387=>x"5500", 388=>x"5700", 389=>x"a500", 390=>x"5b00", 391=>x"5b00", 392=>x"6100",
---- 393=>x"5700", 394=>x"5400", 395=>x"5600", 396=>x"5700", 397=>x"5b00", 398=>x"6000", 399=>x"5d00",
---- 400=>x"5800", 401=>x"5400", 402=>x"5500", 403=>x"5b00", 404=>x"5800", 405=>x"5900", 406=>x"5c00",
---- 407=>x"5800", 408=>x"5b00", 409=>x"5800", 410=>x"5600", 411=>x"5c00", 412=>x"5d00", 413=>x"5b00",
---- 414=>x"5b00", 415=>x"5d00", 416=>x"5500", 417=>x"5700", 418=>x"5900", 419=>x"5d00", 420=>x"5d00",
---- 421=>x"5b00", 422=>x"5d00", 423=>x"5d00", 424=>x"5600", 425=>x"5400", 426=>x"5500", 427=>x"5d00",
---- 428=>x"5d00", 429=>x"5c00", 430=>x"5d00", 431=>x"5f00", 432=>x"5b00", 433=>x"5900", 434=>x"5a00",
---- 435=>x"5e00", 436=>x"5c00", 437=>x"5c00", 438=>x"5b00", 439=>x"5a00", 440=>x"5b00", 441=>x"5b00",
---- 442=>x"5a00", 443=>x"5d00", 444=>x"5e00", 445=>x"5a00", 446=>x"5b00", 447=>x"5d00", 448=>x"5c00",
---- 449=>x"5f00", 450=>x"5a00", 451=>x"5b00", 452=>x"5c00", 453=>x"5c00", 454=>x"5d00", 455=>x"5d00",
---- 456=>x"5c00", 457=>x"5f00", 458=>x"5b00", 459=>x"5900", 460=>x"5b00", 461=>x"5900", 462=>x"5700",
---- 463=>x"5900", 464=>x"5700", 465=>x"5900", 466=>x"5a00", 467=>x"5a00", 468=>x"5a00", 469=>x"5900",
---- 470=>x"5600", 471=>x"5900", 472=>x"5d00", 473=>x"5a00", 474=>x"a700", 475=>x"5a00", 476=>x"5800",
---- 477=>x"5700", 478=>x"5800", 479=>x"5a00", 480=>x"5900", 481=>x"5900", 482=>x"5900", 483=>x"5900",
---- 484=>x"5a00", 485=>x"5c00", 486=>x"5b00", 487=>x"5b00", 488=>x"5700", 489=>x"5700", 490=>x"5900",
---- 491=>x"5900", 492=>x"5c00", 493=>x"5a00", 494=>x"5c00", 495=>x"5e00", 496=>x"5c00", 497=>x"5b00",
---- 498=>x"5a00", 499=>x"5d00", 500=>x"5e00", 501=>x"5c00", 502=>x"a100", 503=>x"6000", 504=>x"5d00",
---- 505=>x"5b00", 506=>x"5b00", 507=>x"5c00", 508=>x"5d00", 509=>x"5c00", 510=>x"5f00", 511=>x"6000",
---- 512=>x"5d00", 513=>x"a300", 514=>x"5d00", 515=>x"5e00", 516=>x"5e00", 517=>x"6200", 518=>x"5f00",
---- 519=>x"5e00", 520=>x"5e00", 521=>x"5f00", 522=>x"5f00", 523=>x"6000", 524=>x"6100", 525=>x"6100",
---- 526=>x"6400", 527=>x"6300", 528=>x"5e00", 529=>x"6300", 530=>x"6100", 531=>x"6000", 532=>x"6100",
---- 533=>x"6300", 534=>x"6400", 535=>x"6100", 536=>x"6300", 537=>x"6400", 538=>x"6300", 539=>x"6200",
---- 540=>x"6300", 541=>x"6400", 542=>x"6500", 543=>x"9b00", 544=>x"6400", 545=>x"6400", 546=>x"6100",
---- 547=>x"6300", 548=>x"6600", 549=>x"6200", 550=>x"6300", 551=>x"6500", 552=>x"6300", 553=>x"6500",
---- 554=>x"6400", 555=>x"6500", 556=>x"6700", 557=>x"6300", 558=>x"6300", 559=>x"6300", 560=>x"6300",
---- 561=>x"6300", 562=>x"6400", 563=>x"6400", 564=>x"6300", 565=>x"6400", 566=>x"6500", 567=>x"6300",
---- 568=>x"6500", 569=>x"6400", 570=>x"6300", 571=>x"6100", 572=>x"6200", 573=>x"6200", 574=>x"6400",
---- 575=>x"6200", 576=>x"6500", 577=>x"6500", 578=>x"6300", 579=>x"6300", 580=>x"6400", 581=>x"6300",
---- 582=>x"6200", 583=>x"6500", 584=>x"6200", 585=>x"6300", 586=>x"6400", 587=>x"6500", 588=>x"6700",
---- 589=>x"6500", 590=>x"6100", 591=>x"6200", 592=>x"6500", 593=>x"6300", 594=>x"6300", 595=>x"6400",
---- 596=>x"6500", 597=>x"5f00", 598=>x"6200", 599=>x"6300", 600=>x"6a00", 601=>x"6500", 602=>x"6000",
---- 603=>x"6400", 604=>x"6300", 605=>x"6000", 606=>x"6100", 607=>x"6000", 608=>x"6200", 609=>x"6000",
---- 610=>x"5f00", 611=>x"6300", 612=>x"6500", 613=>x"6500", 614=>x"6000", 615=>x"6000", 616=>x"6000",
---- 617=>x"6200", 618=>x"6500", 619=>x"6200", 620=>x"9f00", 621=>x"6300", 622=>x"6100", 623=>x"6000",
---- 624=>x"6100", 625=>x"6100", 626=>x"6200", 627=>x"6100", 628=>x"6100", 629=>x"6200", 630=>x"6100",
---- 631=>x"6200", 632=>x"6100", 633=>x"6100", 634=>x"5e00", 635=>x"6400", 636=>x"6000", 637=>x"5d00",
---- 638=>x"6000", 639=>x"6000", 640=>x"6300", 641=>x"6100", 642=>x"5f00", 643=>x"5e00", 644=>x"5d00",
---- 645=>x"5e00", 646=>x"5d00", 647=>x"6000", 648=>x"5d00", 649=>x"6500", 650=>x"5f00", 651=>x"5e00",
---- 652=>x"5e00", 653=>x"a000", 654=>x"6000", 655=>x"5e00", 656=>x"5f00", 657=>x"6300", 658=>x"6200",
---- 659=>x"5e00", 660=>x"5e00", 661=>x"6100", 662=>x"6000", 663=>x"5d00", 664=>x"5f00", 665=>x"6000",
---- 666=>x"6300", 667=>x"5e00", 668=>x"5b00", 669=>x"5d00", 670=>x"5f00", 671=>x"5f00", 672=>x"6000",
---- 673=>x"6000", 674=>x"6400", 675=>x"6200", 676=>x"9f00", 677=>x"5f00", 678=>x"6000", 679=>x"6000",
---- 680=>x"5e00", 681=>x"6000", 682=>x"6000", 683=>x"6000", 684=>x"6500", 685=>x"6100", 686=>x"5e00",
---- 687=>x"5e00", 688=>x"6400", 689=>x"6100", 690=>x"6200", 691=>x"6200", 692=>x"5f00", 693=>x"6100",
---- 694=>x"6100", 695=>x"6100", 696=>x"6300", 697=>x"6300", 698=>x"6200", 699=>x"6300", 700=>x"6000",
---- 701=>x"6100", 702=>x"6300", 703=>x"6200", 704=>x"6200", 705=>x"6300", 706=>x"9f00", 707=>x"6200",
---- 708=>x"6300", 709=>x"6100", 710=>x"6000", 711=>x"6200", 712=>x"6200", 713=>x"6400", 714=>x"6200",
---- 715=>x"6200", 716=>x"6100", 717=>x"6500", 718=>x"6100", 719=>x"6300", 720=>x"6300", 721=>x"6400",
---- 722=>x"6400", 723=>x"6600", 724=>x"9c00", 725=>x"6300", 726=>x"6200", 727=>x"6200", 728=>x"6000",
---- 729=>x"6200", 730=>x"6500", 731=>x"6800", 732=>x"6600", 733=>x"6200", 734=>x"6300", 735=>x"6300",
---- 736=>x"6100", 737=>x"6400", 738=>x"6500", 739=>x"6800", 740=>x"6900", 741=>x"6500", 742=>x"6200",
---- 743=>x"6000", 744=>x"6400", 745=>x"6500", 746=>x"6600", 747=>x"6600", 748=>x"6600", 749=>x"6500",
---- 750=>x"6300", 751=>x"5e00", 752=>x"6700", 753=>x"6800", 754=>x"6700", 755=>x"6800", 756=>x"6700",
---- 757=>x"6400", 758=>x"6100", 759=>x"6100", 760=>x"6a00", 761=>x"6800", 762=>x"6b00", 763=>x"9700",
---- 764=>x"6700", 765=>x"6300", 766=>x"9f00", 767=>x"6300", 768=>x"6a00", 769=>x"6900", 770=>x"6900",
---- 771=>x"6a00", 772=>x"6600", 773=>x"6600", 774=>x"6700", 775=>x"6600", 776=>x"7000", 777=>x"6900",
---- 778=>x"6600", 779=>x"6800", 780=>x"6600", 781=>x"6600", 782=>x"6900", 783=>x"6300", 784=>x"6d00",
---- 785=>x"6b00", 786=>x"6900", 787=>x"6800", 788=>x"6700", 789=>x"6700", 790=>x"6800", 791=>x"6400",
---- 792=>x"6a00", 793=>x"6b00", 794=>x"6b00", 795=>x"6800", 796=>x"6800", 797=>x"9600", 798=>x"6700",
---- 799=>x"6300", 800=>x"6800", 801=>x"6800", 802=>x"6900", 803=>x"6900", 804=>x"6800", 805=>x"6600",
---- 806=>x"6400", 807=>x"6400", 808=>x"6f00", 809=>x"6b00", 810=>x"6a00", 811=>x"6c00", 812=>x"6a00",
---- 813=>x"6800", 814=>x"6700", 815=>x"6300", 816=>x"6c00", 817=>x"6d00", 818=>x"6c00", 819=>x"6d00",
---- 820=>x"6c00", 821=>x"6b00", 822=>x"6a00", 823=>x"6400", 824=>x"6d00", 825=>x"6c00", 826=>x"6a00",
---- 827=>x"6b00", 828=>x"6900", 829=>x"6600", 830=>x"6800", 831=>x"6700", 832=>x"6b00", 833=>x"6b00",
---- 834=>x"6c00", 835=>x"6b00", 836=>x"6800", 837=>x"6700", 838=>x"6800", 839=>x"9b00", 840=>x"6b00",
---- 841=>x"6c00", 842=>x"6d00", 843=>x"6b00", 844=>x"6700", 845=>x"9a00", 846=>x"6700", 847=>x"6700",
---- 848=>x"6b00", 849=>x"6c00", 850=>x"6d00", 851=>x"6900", 852=>x"6600", 853=>x"6900", 854=>x"6600",
---- 855=>x"6500", 856=>x"6900", 857=>x"6d00", 858=>x"6b00", 859=>x"6800", 860=>x"6900", 861=>x"6800",
---- 862=>x"6700", 863=>x"6400", 864=>x"9200", 865=>x"6900", 866=>x"6900", 867=>x"6900", 868=>x"6900",
---- 869=>x"6800", 870=>x"6800", 871=>x"6100", 872=>x"6a00", 873=>x"6a00", 874=>x"6600", 875=>x"6a00",
---- 876=>x"6a00", 877=>x"6b00", 878=>x"6900", 879=>x"6500", 880=>x"6800", 881=>x"6b00", 882=>x"6900",
---- 883=>x"6a00", 884=>x"6a00", 885=>x"6800", 886=>x"6800", 887=>x"6600", 888=>x"6600", 889=>x"6800",
---- 890=>x"6a00", 891=>x"6900", 892=>x"6800", 893=>x"6400", 894=>x"6400", 895=>x"6400", 896=>x"6500",
---- 897=>x"6600", 898=>x"6700", 899=>x"6600", 900=>x"6900", 901=>x"6800", 902=>x"6700", 903=>x"6800",
---- 904=>x"6300", 905=>x"6700", 906=>x"6a00", 907=>x"6600", 908=>x"6700", 909=>x"6800", 910=>x"6700",
---- 911=>x"6500", 912=>x"6900", 913=>x"6a00", 914=>x"6900", 915=>x"6800", 916=>x"6700", 917=>x"6600",
---- 918=>x"6600", 919=>x"6600", 920=>x"6700", 921=>x"6a00", 922=>x"6b00", 923=>x"6700", 924=>x"6700",
---- 925=>x"6300", 926=>x"6300", 927=>x"6500", 928=>x"6900", 929=>x"6900", 930=>x"6a00", 931=>x"6900",
---- 932=>x"6600", 933=>x"6000", 934=>x"6200", 935=>x"6400", 936=>x"6700", 937=>x"6a00", 938=>x"6900",
---- 939=>x"9800", 940=>x"6500", 941=>x"6400", 942=>x"6400", 943=>x"6300", 944=>x"6500", 945=>x"6700",
---- 946=>x"6700", 947=>x"6500", 948=>x"6300", 949=>x"6600", 950=>x"6300", 951=>x"6300", 952=>x"6400",
---- 953=>x"6700", 954=>x"6600", 955=>x"6700", 956=>x"6700", 957=>x"6300", 958=>x"6300", 959=>x"6000",
---- 960=>x"6600", 961=>x"6700", 962=>x"6700", 963=>x"6600", 964=>x"6600", 965=>x"6300", 966=>x"6300",
---- 967=>x"5f00", 968=>x"6100", 969=>x"6700", 970=>x"6600", 971=>x"6300", 972=>x"6500", 973=>x"6200",
---- 974=>x"6200", 975=>x"6000", 976=>x"6600", 977=>x"6700", 978=>x"6600", 979=>x"6500", 980=>x"6300",
---- 981=>x"5f00", 982=>x"6400", 983=>x"6300", 984=>x"6300", 985=>x"6400", 986=>x"6300", 987=>x"6400",
---- 988=>x"6400", 989=>x"6300", 990=>x"6300", 991=>x"6300", 992=>x"6300", 993=>x"6400", 994=>x"6500",
---- 995=>x"6400", 996=>x"6500", 997=>x"9900", 998=>x"6600", 999=>x"6400", 1000=>x"9700", 1001=>x"6800",
---- 1002=>x"6800", 1003=>x"6600", 1004=>x"6600", 1005=>x"6400", 1006=>x"6300", 1007=>x"6400", 1008=>x"6500",
---- 1009=>x"9b00", 1010=>x"6500", 1011=>x"6500", 1012=>x"6700", 1013=>x"6a00", 1014=>x"6600", 1015=>x"6400",
---- 1016=>x"6200", 1017=>x"6500", 1018=>x"6600", 1019=>x"6700", 1020=>x"6800", 1021=>x"6800", 1022=>x"6800",
---- 1023=>x"6600", 1024=>x"6300", 1025=>x"6500", 1026=>x"6400", 1027=>x"6800", 1028=>x"6a00", 1029=>x"6600",
---- 1030=>x"6500", 1031=>x"6300", 1032=>x"6300", 1033=>x"6600", 1034=>x"6500", 1035=>x"6500", 1036=>x"6400",
---- 1037=>x"6400", 1038=>x"6200", 1039=>x"6300", 1040=>x"6000", 1041=>x"6500", 1042=>x"6500", 1043=>x"6000",
---- 1044=>x"6200", 1045=>x"6300", 1046=>x"6100", 1047=>x"5f00", 1048=>x"5e00", 1049=>x"5d00", 1050=>x"6000",
---- 1051=>x"5f00", 1052=>x"5d00", 1053=>x"5f00", 1054=>x"5d00", 1055=>x"5b00", 1056=>x"6000", 1057=>x"6100",
---- 1058=>x"6200", 1059=>x"5f00", 1060=>x"5e00", 1061=>x"5e00", 1062=>x"5d00", 1063=>x"5b00", 1064=>x"6100",
---- 1065=>x"6400", 1066=>x"6300", 1067=>x"5f00", 1068=>x"5f00", 1069=>x"5d00", 1070=>x"5f00", 1071=>x"5f00",
---- 1072=>x"6600", 1073=>x"6200", 1074=>x"6300", 1075=>x"6100", 1076=>x"6100", 1077=>x"6000", 1078=>x"5f00",
---- 1079=>x"5b00", 1080=>x"6600", 1081=>x"6300", 1082=>x"6300", 1083=>x"6100", 1084=>x"6100", 1085=>x"6100",
---- 1086=>x"9e00", 1087=>x"5c00", 1088=>x"6200", 1089=>x"6500", 1090=>x"6200", 1091=>x"6300", 1092=>x"6200",
---- 1093=>x"6200", 1094=>x"6100", 1095=>x"5b00", 1096=>x"6400", 1097=>x"6300", 1098=>x"6600", 1099=>x"6300",
---- 1100=>x"6000", 1101=>x"6300", 1102=>x"6100", 1103=>x"5c00", 1104=>x"6a00", 1105=>x"6800", 1106=>x"6400",
---- 1107=>x"6400", 1108=>x"6500", 1109=>x"6700", 1110=>x"6000", 1111=>x"5900", 1112=>x"6700", 1113=>x"6500",
---- 1114=>x"6800", 1115=>x"6a00", 1116=>x"6400", 1117=>x"6500", 1118=>x"5e00", 1119=>x"5a00", 1120=>x"6800",
---- 1121=>x"6600", 1122=>x"6700", 1123=>x"6700", 1124=>x"6200", 1125=>x"6300", 1126=>x"5d00", 1127=>x"5900",
---- 1128=>x"6500", 1129=>x"6600", 1130=>x"6400", 1131=>x"6200", 1132=>x"5e00", 1133=>x"6000", 1134=>x"5c00",
---- 1135=>x"5700", 1136=>x"6600", 1137=>x"6400", 1138=>x"6200", 1139=>x"6000", 1140=>x"5e00", 1141=>x"5a00",
---- 1142=>x"5800", 1143=>x"5300", 1144=>x"6500", 1145=>x"6100", 1146=>x"5d00", 1147=>x"a600", 1148=>x"5c00",
---- 1149=>x"5800", 1150=>x"5200", 1151=>x"5000", 1152=>x"5f00", 1153=>x"5d00", 1154=>x"5b00", 1155=>x"5900",
---- 1156=>x"5800", 1157=>x"5500", 1158=>x"5300", 1159=>x"5000", 1160=>x"5a00", 1161=>x"5c00", 1162=>x"5e00",
---- 1163=>x"5b00", 1164=>x"ab00", 1165=>x"5500", 1166=>x"5400", 1167=>x"5100", 1168=>x"5a00", 1169=>x"5b00",
---- 1170=>x"6300", 1171=>x"5a00", 1172=>x"5500", 1173=>x"ac00", 1174=>x"5200", 1175=>x"5200", 1176=>x"5600",
---- 1177=>x"5300", 1178=>x"5800", 1179=>x"5800", 1180=>x"5100", 1181=>x"4e00", 1182=>x"5100", 1183=>x"5000",
---- 1184=>x"5200", 1185=>x"5400", 1186=>x"5200", 1187=>x"5000", 1188=>x"4f00", 1189=>x"4c00", 1190=>x"4e00",
---- 1191=>x"5100", 1192=>x"5400", 1193=>x"5100", 1194=>x"4e00", 1195=>x"4f00", 1196=>x"4e00", 1197=>x"4c00",
---- 1198=>x"4b00", 1199=>x"4d00", 1200=>x"5100", 1201=>x"5100", 1202=>x"4c00", 1203=>x"4b00", 1204=>x"4900",
---- 1205=>x"4b00", 1206=>x"4800", 1207=>x"4600", 1208=>x"4b00", 1209=>x"4c00", 1210=>x"4a00", 1211=>x"4a00",
---- 1212=>x"4a00", 1213=>x"4c00", 1214=>x"4a00", 1215=>x"b600", 1216=>x"4c00", 1217=>x"4b00", 1218=>x"4d00",
---- 1219=>x"4b00", 1220=>x"4a00", 1221=>x"4b00", 1222=>x"4e00", 1223=>x"4900", 1224=>x"5300", 1225=>x"4d00",
---- 1226=>x"4a00", 1227=>x"4c00", 1228=>x"4b00", 1229=>x"4c00", 1230=>x"4900", 1231=>x"4800", 1232=>x"4f00",
---- 1233=>x"4d00", 1234=>x"4c00", 1235=>x"4c00", 1236=>x"5000", 1237=>x"4d00", 1238=>x"4c00", 1239=>x"4900",
---- 1240=>x"4e00", 1241=>x"4f00", 1242=>x"4d00", 1243=>x"4b00", 1244=>x"4a00", 1245=>x"4a00", 1246=>x"4b00",
---- 1247=>x"4700", 1248=>x"5000", 1249=>x"5200", 1250=>x"5200", 1251=>x"4a00", 1252=>x"4a00", 1253=>x"4700",
---- 1254=>x"4700", 1255=>x"4800", 1256=>x"5100", 1257=>x"4f00", 1258=>x"4f00", 1259=>x"4c00", 1260=>x"4d00",
---- 1261=>x"4b00", 1262=>x"4c00", 1263=>x"4a00", 1264=>x"5300", 1265=>x"5000", 1266=>x"4e00", 1267=>x"4f00",
---- 1268=>x"4f00", 1269=>x"4e00", 1270=>x"4a00", 1271=>x"4800", 1272=>x"5500", 1273=>x"5600", 1274=>x"5300",
---- 1275=>x"5100", 1276=>x"4f00", 1277=>x"4c00", 1278=>x"4900", 1279=>x"4500", 1280=>x"5900", 1281=>x"5600",
---- 1282=>x"5100", 1283=>x"5000", 1284=>x"5000", 1285=>x"4c00", 1286=>x"4c00", 1287=>x"4900", 1288=>x"5600",
---- 1289=>x"5400", 1290=>x"4f00", 1291=>x"5100", 1292=>x"5100", 1293=>x"4d00", 1294=>x"4b00", 1295=>x"4b00",
---- 1296=>x"4f00", 1297=>x"5100", 1298=>x"5000", 1299=>x"4f00", 1300=>x"4c00", 1301=>x"4e00", 1302=>x"4f00",
---- 1303=>x"4c00", 1304=>x"4f00", 1305=>x"5200", 1306=>x"4e00", 1307=>x"4d00", 1308=>x"4d00", 1309=>x"4e00",
---- 1310=>x"4d00", 1311=>x"4900", 1312=>x"4c00", 1313=>x"5200", 1314=>x"4d00", 1315=>x"4f00", 1316=>x"4e00",
---- 1317=>x"4a00", 1318=>x"4a00", 1319=>x"4900", 1320=>x"4d00", 1321=>x"4f00", 1322=>x"4f00", 1323=>x"4d00",
---- 1324=>x"4800", 1325=>x"4c00", 1326=>x"5000", 1327=>x"4b00", 1328=>x"4e00", 1329=>x"5000", 1330=>x"4e00",
---- 1331=>x"4900", 1332=>x"4e00", 1333=>x"4f00", 1334=>x"5200", 1335=>x"4c00", 1336=>x"5100", 1337=>x"5100",
---- 1338=>x"4b00", 1339=>x"4b00", 1340=>x"5000", 1341=>x"5000", 1342=>x"4c00", 1343=>x"4900", 1344=>x"4b00",
---- 1345=>x"4c00", 1346=>x"b800", 1347=>x"4800", 1348=>x"4a00", 1349=>x"4900", 1350=>x"4c00", 1351=>x"4a00",
---- 1352=>x"4800", 1353=>x"4a00", 1354=>x"4600", 1355=>x"4a00", 1356=>x"4800", 1357=>x"4700", 1358=>x"4c00",
---- 1359=>x"4700", 1360=>x"4900", 1361=>x"4b00", 1362=>x"4700", 1363=>x"4800", 1364=>x"4600", 1365=>x"4300",
---- 1366=>x"4500", 1367=>x"4500", 1368=>x"4b00", 1369=>x"4700", 1370=>x"4600", 1371=>x"4500", 1372=>x"ba00",
---- 1373=>x"4400", 1374=>x"4400", 1375=>x"4500", 1376=>x"4700", 1377=>x"4200", 1378=>x"3d00", 1379=>x"4100",
---- 1380=>x"4300", 1381=>x"4500", 1382=>x"4600", 1383=>x"4300", 1384=>x"4800", 1385=>x"4000", 1386=>x"3c00",
---- 1387=>x"3d00", 1388=>x"4100", 1389=>x"4500", 1390=>x"4600", 1391=>x"4400", 1392=>x"3d00", 1393=>x"3c00",
---- 1394=>x"3900", 1395=>x"3b00", 1396=>x"3d00", 1397=>x"3c00", 1398=>x"4200", 1399=>x"4500", 1400=>x"3800",
---- 1401=>x"3700", 1402=>x"c600", 1403=>x"3b00", 1404=>x"3c00", 1405=>x"3e00", 1406=>x"4300", 1407=>x"4000",
---- 1408=>x"3800", 1409=>x"3800", 1410=>x"3600", 1411=>x"3900", 1412=>x"3c00", 1413=>x"3e00", 1414=>x"4300",
---- 1415=>x"4000", 1416=>x"3500", 1417=>x"3700", 1418=>x"3a00", 1419=>x"3a00", 1420=>x"3b00", 1421=>x"3b00",
---- 1422=>x"4000", 1423=>x"4000", 1424=>x"3800", 1425=>x"3800", 1426=>x"3b00", 1427=>x"3900", 1428=>x"3b00",
---- 1429=>x"3d00", 1430=>x"4200", 1431=>x"4000", 1432=>x"3600", 1433=>x"3800", 1434=>x"3600", 1435=>x"3800",
---- 1436=>x"3b00", 1437=>x"3d00", 1438=>x"3e00", 1439=>x"3f00", 1440=>x"3c00", 1441=>x"3700", 1442=>x"3500",
---- 1443=>x"3700", 1444=>x"3900", 1445=>x"3600", 1446=>x"3c00", 1447=>x"3b00", 1448=>x"3600", 1449=>x"3100",
---- 1450=>x"3400", 1451=>x"3700", 1452=>x"3700", 1453=>x"3700", 1454=>x"3900", 1455=>x"3700", 1456=>x"3b00",
---- 1457=>x"3400", 1458=>x"3000", 1459=>x"3200", 1460=>x"3300", 1461=>x"3a00", 1462=>x"3900", 1463=>x"3900",
---- 1464=>x"3400", 1465=>x"3200", 1466=>x"3200", 1467=>x"3700", 1468=>x"3300", 1469=>x"3400", 1470=>x"3300",
---- 1471=>x"3100", 1472=>x"3400", 1473=>x"3100", 1474=>x"3300", 1475=>x"3600", 1476=>x"3300", 1477=>x"3200",
---- 1478=>x"3200", 1479=>x"3100", 1480=>x"3800", 1481=>x"3300", 1482=>x"3200", 1483=>x"3300", 1484=>x"3000",
---- 1485=>x"3100", 1486=>x"2f00", 1487=>x"3000", 1488=>x"3200", 1489=>x"3100", 1490=>x"3000", 1491=>x"3300",
---- 1492=>x"3200", 1493=>x"3100", 1494=>x"3000", 1495=>x"2f00", 1496=>x"2d00", 1497=>x"3000", 1498=>x"2f00",
---- 1499=>x"2f00", 1500=>x"3400", 1501=>x"3100", 1502=>x"3200", 1503=>x"3400", 1504=>x"d100", 1505=>x"2f00",
---- 1506=>x"2d00", 1507=>x"3100", 1508=>x"3000", 1509=>x"2f00", 1510=>x"3200", 1511=>x"3000", 1512=>x"2e00",
---- 1513=>x"2e00", 1514=>x"3200", 1515=>x"3600", 1516=>x"2e00", 1517=>x"2a00", 1518=>x"3000", 1519=>x"3100",
---- 1520=>x"3100", 1521=>x"2e00", 1522=>x"3200", 1523=>x"3700", 1524=>x"3100", 1525=>x"2e00", 1526=>x"3000",
---- 1527=>x"3000", 1528=>x"3400", 1529=>x"3100", 1530=>x"2f00", 1531=>x"2f00", 1532=>x"2e00", 1533=>x"2c00",
---- 1534=>x"2e00", 1535=>x"3000", 1536=>x"2b00", 1537=>x"2b00", 1538=>x"2d00", 1539=>x"2f00", 1540=>x"3000",
---- 1541=>x"2c00", 1542=>x"2900", 1543=>x"3000", 1544=>x"2e00", 1545=>x"2c00", 1546=>x"2f00", 1547=>x"3200",
---- 1548=>x"2d00", 1549=>x"2b00", 1550=>x"2c00", 1551=>x"2c00", 1552=>x"2f00", 1553=>x"2e00", 1554=>x"3000",
---- 1555=>x"3200", 1556=>x"2c00", 1557=>x"2900", 1558=>x"2c00", 1559=>x"2900", 1560=>x"3300", 1561=>x"3700",
---- 1562=>x"3600", 1563=>x"3500", 1564=>x"3100", 1565=>x"d600", 1566=>x"2700", 1567=>x"2800", 1568=>x"3800",
---- 1569=>x"c800", 1570=>x"3b00", 1571=>x"3d00", 1572=>x"3200", 1573=>x"3000", 1574=>x"2a00", 1575=>x"2800",
---- 1576=>x"3e00", 1577=>x"4000", 1578=>x"4200", 1579=>x"3e00", 1580=>x"3700", 1581=>x"3300", 1582=>x"3400",
---- 1583=>x"3000", 1584=>x"5f00", 1585=>x"5500", 1586=>x"4a00", 1587=>x"4500", 1588=>x"3d00", 1589=>x"3700",
---- 1590=>x"3400", 1591=>x"3400", 1592=>x"7b00", 1593=>x"7500", 1594=>x"6800", 1595=>x"5900", 1596=>x"4c00",
---- 1597=>x"b900", 1598=>x"3d00", 1599=>x"3600", 1600=>x"8100", 1601=>x"8100", 1602=>x"7e00", 1603=>x"7200",
---- 1604=>x"6000", 1605=>x"5500", 1606=>x"4f00", 1607=>x"4000", 1608=>x"8900", 1609=>x"8600", 1610=>x"8400",
---- 1611=>x"8300", 1612=>x"7600", 1613=>x"6800", 1614=>x"5b00", 1615=>x"5000", 1616=>x"8b00", 1617=>x"8700",
---- 1618=>x"8b00", 1619=>x"8800", 1620=>x"8200", 1621=>x"7b00", 1622=>x"6d00", 1623=>x"6100", 1624=>x"8700",
---- 1625=>x"8500", 1626=>x"8b00", 1627=>x"8e00", 1628=>x"8d00", 1629=>x"8900", 1630=>x"7e00", 1631=>x"7200",
---- 1632=>x"8000", 1633=>x"8300", 1634=>x"8b00", 1635=>x"9200", 1636=>x"9700", 1637=>x"9200", 1638=>x"8c00",
---- 1639=>x"8100", 1640=>x"7c00", 1641=>x"8300", 1642=>x"8b00", 1643=>x"9100", 1644=>x"9700", 1645=>x"9500",
---- 1646=>x"9300", 1647=>x"8e00", 1648=>x"8200", 1649=>x"7d00", 1650=>x"8200", 1651=>x"8e00", 1652=>x"9600",
---- 1653=>x"9800", 1654=>x"9800", 1655=>x"9100", 1656=>x"6700", 1657=>x"6c00", 1658=>x"7a00", 1659=>x"8800",
---- 1660=>x"8f00", 1661=>x"9500", 1662=>x"9b00", 1663=>x"9700", 1664=>x"4700", 1665=>x"5000", 1666=>x"6e00",
---- 1667=>x"7f00", 1668=>x"8a00", 1669=>x"9400", 1670=>x"9f00", 1671=>x"9f00", 1672=>x"2e00", 1673=>x"3c00",
---- 1674=>x"5f00", 1675=>x"7700", 1676=>x"8400", 1677=>x"9200", 1678=>x"a400", 1679=>x"a400", 1680=>x"2300",
---- 1681=>x"2e00", 1682=>x"4c00", 1683=>x"6c00", 1684=>x"7e00", 1685=>x"9800", 1686=>x"a400", 1687=>x"a400",
---- 1688=>x"2300", 1689=>x"2800", 1690=>x"3600", 1691=>x"5300", 1692=>x"8d00", 1693=>x"9600", 1694=>x"a500",
---- 1695=>x"a800", 1696=>x"2000", 1697=>x"2200", 1698=>x"2a00", 1699=>x"4100", 1700=>x"7200", 1701=>x"9300",
---- 1702=>x"a400", 1703=>x"a900", 1704=>x"2400", 1705=>x"2300", 1706=>x"2a00", 1707=>x"3f00", 1708=>x"6e00",
---- 1709=>x"9400", 1710=>x"a500", 1711=>x"ab00", 1712=>x"2000", 1713=>x"2700", 1714=>x"2c00", 1715=>x"3900",
---- 1716=>x"6200", 1717=>x"8c00", 1718=>x"a300", 1719=>x"ad00", 1720=>x"1f00", 1721=>x"2400", 1722=>x"2c00",
---- 1723=>x"3c00", 1724=>x"5e00", 1725=>x"8b00", 1726=>x"9e00", 1727=>x"aa00", 1728=>x"1f00", 1729=>x"2000",
---- 1730=>x"2200", 1731=>x"cd00", 1732=>x"5900", 1733=>x"8900", 1734=>x"9a00", 1735=>x"a400", 1736=>x"1e00",
---- 1737=>x"2100", 1738=>x"2100", 1739=>x"d500", 1740=>x"5300", 1741=>x"8500", 1742=>x"9a00", 1743=>x"a600",
---- 1744=>x"1f00", 1745=>x"2000", 1746=>x"1e00", 1747=>x"2800", 1748=>x"4a00", 1749=>x"7c00", 1750=>x"9c00",
---- 1751=>x"a800", 1752=>x"1e00", 1753=>x"2000", 1754=>x"2200", 1755=>x"2b00", 1756=>x"4c00", 1757=>x"7a00",
---- 1758=>x"9a00", 1759=>x"aa00", 1760=>x"1d00", 1761=>x"2000", 1762=>x"1f00", 1763=>x"2800", 1764=>x"4b00",
---- 1765=>x"7b00", 1766=>x"9700", 1767=>x"a600", 1768=>x"2000", 1769=>x"1f00", 1770=>x"2000", 1771=>x"2600",
---- 1772=>x"4600", 1773=>x"7d00", 1774=>x"9500", 1775=>x"a400", 1776=>x"1e00", 1777=>x"1d00", 1778=>x"2000",
---- 1779=>x"2500", 1780=>x"4400", 1781=>x"7200", 1782=>x"9600", 1783=>x"a500", 1784=>x"2000", 1785=>x"1e00",
---- 1786=>x"2000", 1787=>x"2600", 1788=>x"4000", 1789=>x"6c00", 1790=>x"9400", 1791=>x"a400", 1792=>x"2000",
---- 1793=>x"2000", 1794=>x"2100", 1795=>x"2500", 1796=>x"ca00", 1797=>x"6500", 1798=>x"8f00", 1799=>x"a000",
---- 1800=>x"2500", 1801=>x"2400", 1802=>x"2400", 1803=>x"2800", 1804=>x"3100", 1805=>x"6300", 1806=>x"8b00",
---- 1807=>x"9d00", 1808=>x"2200", 1809=>x"2300", 1810=>x"2200", 1811=>x"2300", 1812=>x"3100", 1813=>x"5b00",
---- 1814=>x"8900", 1815=>x"9b00", 1816=>x"2800", 1817=>x"2700", 1818=>x"2600", 1819=>x"2300", 1820=>x"2c00",
---- 1821=>x"5300", 1822=>x"8200", 1823=>x"9b00", 1824=>x"2a00", 1825=>x"2900", 1826=>x"2500", 1827=>x"2100",
---- 1828=>x"2900", 1829=>x"4c00", 1830=>x"7d00", 1831=>x"9900", 1832=>x"2600", 1833=>x"2500", 1834=>x"2400",
---- 1835=>x"2700", 1836=>x"2900", 1837=>x"4600", 1838=>x"7800", 1839=>x"9900", 1840=>x"2600", 1841=>x"2600",
---- 1842=>x"2200", 1843=>x"2400", 1844=>x"2500", 1845=>x"4b00", 1846=>x"8100", 1847=>x"6700", 1848=>x"2400",
---- 1849=>x"2400", 1850=>x"1f00", 1851=>x"2400", 1852=>x"2800", 1853=>x"4900", 1854=>x"7600", 1855=>x"9100",
---- 1856=>x"2300", 1857=>x"2500", 1858=>x"2200", 1859=>x"2300", 1860=>x"2800", 1861=>x"3d00", 1862=>x"6900",
---- 1863=>x"9800", 1864=>x"2100", 1865=>x"2100", 1866=>x"2000", 1867=>x"2400", 1868=>x"2900", 1869=>x"3200",
---- 1870=>x"6800", 1871=>x"9d00", 1872=>x"2500", 1873=>x"2300", 1874=>x"2200", 1875=>x"1e00", 1876=>x"2100",
---- 1877=>x"3100", 1878=>x"6b00", 1879=>x"9800", 1880=>x"2900", 1881=>x"2700", 1882=>x"2200", 1883=>x"2200",
---- 1884=>x"2400", 1885=>x"3100", 1886=>x"6800", 1887=>x"9a00", 1888=>x"2f00", 1889=>x"2d00", 1890=>x"2d00",
---- 1891=>x"3300", 1892=>x"3300", 1893=>x"3600", 1894=>x"6800", 1895=>x"9700", 1896=>x"2f00", 1897=>x"3b00",
---- 1898=>x"4500", 1899=>x"4400", 1900=>x"4000", 1901=>x"4300", 1902=>x"6600", 1903=>x"9200", 1904=>x"4900",
---- 1905=>x"5400", 1906=>x"5400", 1907=>x"5100", 1908=>x"4e00", 1909=>x"5200", 1910=>x"6800", 1911=>x"8a00",
---- 1912=>x"5d00", 1913=>x"5d00", 1914=>x"5a00", 1915=>x"5700", 1916=>x"5b00", 1917=>x"5c00", 1918=>x"7000",
---- 1919=>x"8800", 1920=>x"5400", 1921=>x"5a00", 1922=>x"5a00", 1923=>x"5a00", 1924=>x"6100", 1925=>x"6500",
---- 1926=>x"7700", 1927=>x"8d00", 1928=>x"5500", 1929=>x"5a00", 1930=>x"5a00", 1931=>x"6000", 1932=>x"6500",
---- 1933=>x"6f00", 1934=>x"7f00", 1935=>x"9000", 1936=>x"4900", 1937=>x"5300", 1938=>x"6000", 1939=>x"6800",
---- 1940=>x"6e00", 1941=>x"7600", 1942=>x"8200", 1943=>x"8e00", 1944=>x"3b00", 1945=>x"4f00", 1946=>x"6100",
---- 1947=>x"7000", 1948=>x"7300", 1949=>x"7300", 1950=>x"7b00", 1951=>x"8a00", 1952=>x"3100", 1953=>x"4800",
---- 1954=>x"5e00", 1955=>x"6c00", 1956=>x"9000", 1957=>x"6c00", 1958=>x"6b00", 1959=>x"8400", 1960=>x"2900",
---- 1961=>x"3b00", 1962=>x"5000", 1963=>x"5d00", 1964=>x"5f00", 1965=>x"5f00", 1966=>x"6800", 1967=>x"7f00",
---- 1968=>x"2a00", 1969=>x"3500", 1970=>x"4200", 1971=>x"5200", 1972=>x"5a00", 1973=>x"5d00", 1974=>x"6700",
---- 1975=>x"7b00", 1976=>x"2e00", 1977=>x"3300", 1978=>x"3900", 1979=>x"4600", 1980=>x"5600", 1981=>x"5700",
---- 1982=>x"5e00", 1983=>x"7400", 1984=>x"3300", 1985=>x"3800", 1986=>x"3500", 1987=>x"3c00", 1988=>x"4b00",
---- 1989=>x"aa00", 1990=>x"5600", 1991=>x"6e00", 1992=>x"3500", 1993=>x"3c00", 1994=>x"3f00", 1995=>x"c100",
---- 1996=>x"4300", 1997=>x"4c00", 1998=>x"4f00", 1999=>x"6700", 2000=>x"3200", 2001=>x"3700", 2002=>x"3b00",
---- 2003=>x"3800", 2004=>x"3f00", 2005=>x"3f00", 2006=>x"4400", 2007=>x"6000", 2008=>x"3000", 2009=>x"3700",
---- 2010=>x"3900", 2011=>x"3100", 2012=>x"3c00", 2013=>x"3e00", 2014=>x"4100", 2015=>x"6200", 2016=>x"2f00",
---- 2017=>x"3300", 2018=>x"3500", 2019=>x"3300", 2020=>x"3900", 2021=>x"3a00", 2022=>x"3b00", 2023=>x"6500",
---- 2024=>x"3200", 2025=>x"3400", 2026=>x"3500", 2027=>x"3500", 2028=>x"3900", 2029=>x"3700", 2030=>x"3a00",
---- 2031=>x"6100", 2032=>x"2f00", 2033=>x"3000", 2034=>x"3300", 2035=>x"3200", 2036=>x"3800", 2037=>x"3500",
---- 2038=>x"3800", 2039=>x"5600", 2040=>x"2a00", 2041=>x"3200", 2042=>x"3200", 2043=>x"3200", 2044=>x"3800",
---- 2045=>x"3100", 2046=>x"cd00", 2047=>x"4d00"),
---- 1  => (0=>x"9b00", 1=>x"a000", 2=>x"9d00", 3=>x"9b00", 4=>x"9c00", 5=>x"9a00", 6=>x"9a00", 7=>x"9b00",
---- 8=>x"9b00", 9=>x"a200", 10=>x"9c00", 11=>x"9a00", 12=>x"9c00", 13=>x"9900", 14=>x"9a00",
---- 15=>x"9900", 16=>x"9a00", 17=>x"9f00", 18=>x"9b00", 19=>x"9a00", 20=>x"9c00", 21=>x"9a00",
---- 22=>x"9a00", 23=>x"9a00", 24=>x"9b00", 25=>x"9b00", 26=>x"9a00", 27=>x"9700", 28=>x"9a00",
---- 29=>x"9a00", 30=>x"9800", 31=>x"9a00", 32=>x"9b00", 33=>x"9c00", 34=>x"9b00", 35=>x"9a00",
---- 36=>x"9b00", 37=>x"9a00", 38=>x"9800", 39=>x"9a00", 40=>x"9b00", 41=>x"9b00", 42=>x"9d00",
---- 43=>x"9c00", 44=>x"9800", 45=>x"9900", 46=>x"9c00", 47=>x"9a00", 48=>x"9e00", 49=>x"9d00",
---- 50=>x"9c00", 51=>x"9c00", 52=>x"9a00", 53=>x"9900", 54=>x"6400", 55=>x"6400", 56=>x"9d00",
---- 57=>x"9c00", 58=>x"9b00", 59=>x"9a00", 60=>x"9a00", 61=>x"9a00", 62=>x"9b00", 63=>x"9c00",
---- 64=>x"9a00", 65=>x"9c00", 66=>x"9c00", 67=>x"9b00", 68=>x"9900", 69=>x"9800", 70=>x"9a00",
---- 71=>x"a100", 72=>x"9d00", 73=>x"9f00", 74=>x"9c00", 75=>x"9b00", 76=>x"9b00", 77=>x"9900",
---- 78=>x"9d00", 79=>x"a100", 80=>x"9f00", 81=>x"9f00", 82=>x"9b00", 83=>x"9c00", 84=>x"9b00",
---- 85=>x"9b00", 86=>x"9e00", 87=>x"a000", 88=>x"9f00", 89=>x"9e00", 90=>x"9c00", 91=>x"9c00",
---- 92=>x"9800", 93=>x"9b00", 94=>x"9c00", 95=>x"a200", 96=>x"9f00", 97=>x"9c00", 98=>x"9c00",
---- 99=>x"9e00", 100=>x"9d00", 101=>x"9e00", 102=>x"a100", 103=>x"a400", 104=>x"9e00", 105=>x"9f00",
---- 106=>x"9e00", 107=>x"9c00", 108=>x"9d00", 109=>x"a100", 110=>x"a300", 111=>x"a600", 112=>x"9f00",
---- 113=>x"9f00", 114=>x"9f00", 115=>x"9e00", 116=>x"9e00", 117=>x"a200", 118=>x"a700", 119=>x"a800",
---- 120=>x"9e00", 121=>x"a000", 122=>x"a000", 123=>x"a100", 124=>x"a300", 125=>x"a700", 126=>x"a700",
---- 127=>x"a800", 128=>x"9f00", 129=>x"a200", 130=>x"a000", 131=>x"a300", 132=>x"a700", 133=>x"a800",
---- 134=>x"a800", 135=>x"aa00", 136=>x"a100", 137=>x"a100", 138=>x"a300", 139=>x"a500", 140=>x"a800",
---- 141=>x"a700", 142=>x"a800", 143=>x"a800", 144=>x"a300", 145=>x"a400", 146=>x"a500", 147=>x"a700",
---- 148=>x"a800", 149=>x"a800", 150=>x"a800", 151=>x"a900", 152=>x"a300", 153=>x"5900", 154=>x"a800",
---- 155=>x"a900", 156=>x"a700", 157=>x"a800", 158=>x"a700", 159=>x"a400", 160=>x"a400", 161=>x"a700",
---- 162=>x"a900", 163=>x"a700", 164=>x"a500", 165=>x"a400", 166=>x"5e00", 167=>x"a200", 168=>x"a800",
---- 169=>x"a900", 170=>x"a900", 171=>x"a200", 172=>x"a200", 173=>x"a200", 174=>x"9e00", 175=>x"a100",
---- 176=>x"ab00", 177=>x"ab00", 178=>x"a700", 179=>x"a000", 180=>x"9c00", 181=>x"9e00", 182=>x"9a00",
---- 183=>x"9d00", 184=>x"a900", 185=>x"a500", 186=>x"a000", 187=>x"9c00", 188=>x"9a00", 189=>x"9a00",
---- 190=>x"9900", 191=>x"9700", 192=>x"ab00", 193=>x"a400", 194=>x"9e00", 195=>x"6500", 196=>x"9700",
---- 197=>x"9500", 198=>x"9400", 199=>x"9500", 200=>x"a900", 201=>x"a200", 202=>x"9c00", 203=>x"9600",
---- 204=>x"9200", 205=>x"6e00", 206=>x"8e00", 207=>x"9100", 208=>x"a800", 209=>x"a000", 210=>x"9900",
---- 211=>x"6d00", 212=>x"8c00", 213=>x"8c00", 214=>x"8d00", 215=>x"8a00", 216=>x"a300", 217=>x"9f00",
---- 218=>x"9500", 219=>x"8f00", 220=>x"8700", 221=>x"8200", 222=>x"8700", 223=>x"8a00", 224=>x"9e00",
---- 225=>x"9900", 226=>x"9000", 227=>x"8700", 228=>x"8100", 229=>x"7e00", 230=>x"8000", 231=>x"8a00",
---- 232=>x"9b00", 233=>x"9300", 234=>x"8b00", 235=>x"7e00", 236=>x"7900", 237=>x"7800", 238=>x"8000",
---- 239=>x"8f00", 240=>x"9800", 241=>x"8f00", 242=>x"7f00", 243=>x"7300", 244=>x"6d00", 245=>x"6f00",
---- 246=>x"8000", 247=>x"9000", 248=>x"6a00", 249=>x"8700", 250=>x"7700", 251=>x"6800", 252=>x"6100",
---- 253=>x"7000", 254=>x"8100", 255=>x"8d00", 256=>x"8f00", 257=>x"7d00", 258=>x"6b00", 259=>x"5c00",
---- 260=>x"5a00", 261=>x"7000", 262=>x"8000", 263=>x"8e00", 264=>x"8800", 265=>x"7400", 266=>x"6100",
---- 267=>x"4f00", 268=>x"5900", 269=>x"7000", 270=>x"8100", 271=>x"8e00", 272=>x"7f00", 273=>x"6900",
---- 274=>x"5300", 275=>x"4a00", 276=>x"5700", 277=>x"6f00", 278=>x"8200", 279=>x"8e00", 280=>x"7100",
---- 281=>x"5600", 282=>x"4a00", 283=>x"4c00", 284=>x"5a00", 285=>x"7200", 286=>x"8000", 287=>x"8a00",
---- 288=>x"6600", 289=>x"5000", 290=>x"b600", 291=>x"5000", 292=>x"6000", 293=>x"6e00", 294=>x"8000",
---- 295=>x"8c00", 296=>x"5700", 297=>x"4d00", 298=>x"4d00", 299=>x"ae00", 300=>x"6000", 301=>x"7200",
---- 302=>x"8000", 303=>x"8c00", 304=>x"5300", 305=>x"5300", 306=>x"4c00", 307=>x"5100", 308=>x"5f00",
---- 309=>x"7400", 310=>x"8100", 311=>x"8b00", 312=>x"5400", 313=>x"5700", 314=>x"5100", 315=>x"4f00",
---- 316=>x"5e00", 317=>x"7100", 318=>x"8200", 319=>x"8c00", 320=>x"5200", 321=>x"5300", 322=>x"5600",
---- 323=>x"5200", 324=>x"6000", 325=>x"7400", 326=>x"8200", 327=>x"8e00", 328=>x"5300", 329=>x"5400",
---- 330=>x"5200", 331=>x"5500", 332=>x"5f00", 333=>x"7300", 334=>x"8400", 335=>x"8e00", 336=>x"5600",
---- 337=>x"5500", 338=>x"5300", 339=>x"5700", 340=>x"6000", 341=>x"7200", 342=>x"7f00", 343=>x"8d00",
---- 344=>x"5900", 345=>x"5b00", 346=>x"5400", 347=>x"5700", 348=>x"5f00", 349=>x"7000", 350=>x"8000",
---- 351=>x"8d00", 352=>x"5b00", 353=>x"5900", 354=>x"5300", 355=>x"5600", 356=>x"6300", 357=>x"8d00",
---- 358=>x"8200", 359=>x"7200", 360=>x"5800", 361=>x"5700", 362=>x"5600", 363=>x"5700", 364=>x"9f00",
---- 365=>x"7000", 366=>x"7f00", 367=>x"8e00", 368=>x"5900", 369=>x"5700", 370=>x"5800", 371=>x"5600",
---- 372=>x"5d00", 373=>x"7000", 374=>x"7e00", 375=>x"8c00", 376=>x"5900", 377=>x"5900", 378=>x"5600",
---- 379=>x"5500", 380=>x"5d00", 381=>x"6e00", 382=>x"8000", 383=>x"8c00", 384=>x"5b00", 385=>x"5800",
---- 386=>x"5400", 387=>x"5600", 388=>x"5d00", 389=>x"6f00", 390=>x"8200", 391=>x"8c00", 392=>x"5b00",
---- 393=>x"5b00", 394=>x"5500", 395=>x"5600", 396=>x"6000", 397=>x"6e00", 398=>x"7e00", 399=>x"8700",
---- 400=>x"5c00", 401=>x"5b00", 402=>x"5600", 403=>x"5500", 404=>x"5e00", 405=>x"6c00", 406=>x"7b00",
---- 407=>x"8900", 408=>x"5c00", 409=>x"5a00", 410=>x"5700", 411=>x"5800", 412=>x"5f00", 413=>x"6d00",
---- 414=>x"7d00", 415=>x"8c00", 416=>x"5a00", 417=>x"5b00", 418=>x"5700", 419=>x"5a00", 420=>x"6100",
---- 421=>x"6e00", 422=>x"8000", 423=>x"8b00", 424=>x"5d00", 425=>x"5a00", 426=>x"5900", 427=>x"5b00",
---- 428=>x"6300", 429=>x"7100", 430=>x"8000", 431=>x"8a00", 432=>x"5b00", 433=>x"5b00", 434=>x"5900",
---- 435=>x"5700", 436=>x"5f00", 437=>x"7100", 438=>x"7f00", 439=>x"8a00", 440=>x"5c00", 441=>x"5700",
---- 442=>x"5600", 443=>x"5700", 444=>x"5c00", 445=>x"6f00", 446=>x"7d00", 447=>x"8c00", 448=>x"5b00",
---- 449=>x"5a00", 450=>x"5700", 451=>x"5500", 452=>x"5c00", 453=>x"6a00", 454=>x"7d00", 455=>x"8d00",
---- 456=>x"5600", 457=>x"5500", 458=>x"5400", 459=>x"5300", 460=>x"5c00", 461=>x"6b00", 462=>x"8000",
---- 463=>x"8c00", 464=>x"a300", 465=>x"5900", 466=>x"5400", 467=>x"5400", 468=>x"a600", 469=>x"6a00",
---- 470=>x"7a00", 471=>x"8800", 472=>x"5b00", 473=>x"5800", 474=>x"5300", 475=>x"5400", 476=>x"5600",
---- 477=>x"6900", 478=>x"7b00", 479=>x"8800", 480=>x"5c00", 481=>x"5b00", 482=>x"5800", 483=>x"5400",
---- 484=>x"5b00", 485=>x"6c00", 486=>x"7d00", 487=>x"8700", 488=>x"6000", 489=>x"5c00", 490=>x"5900",
---- 491=>x"5900", 492=>x"5b00", 493=>x"6d00", 494=>x"7c00", 495=>x"8600", 496=>x"6100", 497=>x"5b00",
---- 498=>x"5a00", 499=>x"5600", 500=>x"5b00", 501=>x"6c00", 502=>x"7800", 503=>x"7700", 504=>x"6100",
---- 505=>x"5f00", 506=>x"5d00", 507=>x"5500", 508=>x"5e00", 509=>x"6a00", 510=>x"7900", 511=>x"8800",
---- 512=>x"6000", 513=>x"6000", 514=>x"6300", 515=>x"5e00", 516=>x"6000", 517=>x"6b00", 518=>x"7e00",
---- 519=>x"8500", 520=>x"6100", 521=>x"9d00", 522=>x"6000", 523=>x"5f00", 524=>x"5f00", 525=>x"6d00",
---- 526=>x"7900", 527=>x"8a00", 528=>x"6200", 529=>x"6000", 530=>x"6000", 531=>x"5d00", 532=>x"5f00",
---- 533=>x"6c00", 534=>x"7b00", 535=>x"8a00", 536=>x"6100", 537=>x"6000", 538=>x"5f00", 539=>x"5e00",
---- 540=>x"6100", 541=>x"6900", 542=>x"7b00", 543=>x"8900", 544=>x"6400", 545=>x"6300", 546=>x"6000",
---- 547=>x"6000", 548=>x"6100", 549=>x"6d00", 550=>x"7c00", 551=>x"8900", 552=>x"6400", 553=>x"6200",
---- 554=>x"6300", 555=>x"6100", 556=>x"6600", 557=>x"6e00", 558=>x"7e00", 559=>x"8a00", 560=>x"6500",
---- 561=>x"6100", 562=>x"6000", 563=>x"6200", 564=>x"6900", 565=>x"7100", 566=>x"7f00", 567=>x"8b00",
---- 568=>x"6600", 569=>x"6300", 570=>x"6100", 571=>x"6000", 572=>x"6900", 573=>x"7100", 574=>x"7e00",
---- 575=>x"8a00", 576=>x"6500", 577=>x"6400", 578=>x"6200", 579=>x"6100", 580=>x"6600", 581=>x"7200",
---- 582=>x"7d00", 583=>x"8a00", 584=>x"6400", 585=>x"6200", 586=>x"6300", 587=>x"6400", 588=>x"6600",
---- 589=>x"7200", 590=>x"7e00", 591=>x"8900", 592=>x"6500", 593=>x"6300", 594=>x"6400", 595=>x"6500",
---- 596=>x"6800", 597=>x"7200", 598=>x"7e00", 599=>x"8800", 600=>x"6100", 601=>x"6100", 602=>x"6300",
---- 603=>x"6200", 604=>x"6700", 605=>x"6f00", 606=>x"7a00", 607=>x"8800", 608=>x"6100", 609=>x"6100",
---- 610=>x"6100", 611=>x"5f00", 612=>x"6300", 613=>x"6e00", 614=>x"7900", 615=>x"8a00", 616=>x"6300",
---- 617=>x"6500", 618=>x"5e00", 619=>x"6000", 620=>x"6400", 621=>x"6c00", 622=>x"7b00", 623=>x"8900",
---- 624=>x"9e00", 625=>x"6200", 626=>x"6100", 627=>x"6000", 628=>x"6700", 629=>x"6f00", 630=>x"7c00",
---- 631=>x"8900", 632=>x"6100", 633=>x"6000", 634=>x"5f00", 635=>x"6300", 636=>x"6400", 637=>x"6c00",
---- 638=>x"7e00", 639=>x"8b00", 640=>x"5f00", 641=>x"6000", 642=>x"6000", 643=>x"6500", 644=>x"6200",
---- 645=>x"6e00", 646=>x"7f00", 647=>x"8f00", 648=>x"5e00", 649=>x"6000", 650=>x"5f00", 651=>x"6100",
---- 652=>x"6400", 653=>x"7200", 654=>x"7f00", 655=>x"8c00", 656=>x"5d00", 657=>x"6000", 658=>x"6100",
---- 659=>x"6000", 660=>x"6400", 661=>x"7100", 662=>x"7f00", 663=>x"8c00", 664=>x"5d00", 665=>x"5c00",
---- 666=>x"5f00", 667=>x"6100", 668=>x"6800", 669=>x"7300", 670=>x"8200", 671=>x"8b00", 672=>x"5f00",
---- 673=>x"6000", 674=>x"6200", 675=>x"6400", 676=>x"6800", 677=>x"7600", 678=>x"8100", 679=>x"8d00",
---- 680=>x"6100", 681=>x"6300", 682=>x"6500", 683=>x"6900", 684=>x"6900", 685=>x"7600", 686=>x"7f00",
---- 687=>x"8b00", 688=>x"6200", 689=>x"6200", 690=>x"6700", 691=>x"6a00", 692=>x"6b00", 693=>x"7400",
---- 694=>x"8100", 695=>x"8b00", 696=>x"6300", 697=>x"6300", 698=>x"6700", 699=>x"6900", 700=>x"9400",
---- 701=>x"7400", 702=>x"7f00", 703=>x"8d00", 704=>x"6600", 705=>x"5f00", 706=>x"6400", 707=>x"6700",
---- 708=>x"6d00", 709=>x"7500", 710=>x"8400", 711=>x"8d00", 712=>x"6700", 713=>x"6500", 714=>x"6700",
---- 715=>x"6900", 716=>x"7100", 717=>x"7a00", 718=>x"8400", 719=>x"8e00", 720=>x"6300", 721=>x"6600",
---- 722=>x"6a00", 723=>x"6b00", 724=>x"7000", 725=>x"7800", 726=>x"8500", 727=>x"9100", 728=>x"6400",
---- 729=>x"6400", 730=>x"6900", 731=>x"6e00", 732=>x"6f00", 733=>x"7600", 734=>x"8500", 735=>x"9000",
---- 736=>x"6200", 737=>x"6900", 738=>x"6a00", 739=>x"6c00", 740=>x"7000", 741=>x"7a00", 742=>x"8100",
---- 743=>x"8d00", 744=>x"5f00", 745=>x"6800", 746=>x"6b00", 747=>x"6b00", 748=>x"7100", 749=>x"7a00",
---- 750=>x"8700", 751=>x"8c00", 752=>x"6100", 753=>x"6500", 754=>x"6a00", 755=>x"6c00", 756=>x"6f00",
---- 757=>x"7800", 758=>x"8400", 759=>x"8e00", 760=>x"6300", 761=>x"6300", 762=>x"6700", 763=>x"6b00",
---- 764=>x"6c00", 765=>x"7900", 766=>x"8300", 767=>x"8e00", 768=>x"6500", 769=>x"6400", 770=>x"9b00",
---- 771=>x"6900", 772=>x"6c00", 773=>x"7800", 774=>x"8400", 775=>x"9000", 776=>x"6200", 777=>x"6200",
---- 778=>x"6500", 779=>x"6700", 780=>x"6e00", 781=>x"7600", 782=>x"8200", 783=>x"8f00", 784=>x"6400",
---- 785=>x"6500", 786=>x"6700", 787=>x"6800", 788=>x"6d00", 789=>x"7400", 790=>x"7f00", 791=>x"8d00",
---- 792=>x"6500", 793=>x"6600", 794=>x"6500", 795=>x"6600", 796=>x"6a00", 797=>x"7700", 798=>x"8300",
---- 799=>x"8c00", 800=>x"6600", 801=>x"6400", 802=>x"6600", 803=>x"6600", 804=>x"6700", 805=>x"7200",
---- 806=>x"7d00", 807=>x"8b00", 808=>x"6400", 809=>x"6100", 810=>x"6600", 811=>x"6500", 812=>x"6600",
---- 813=>x"7400", 814=>x"7f00", 815=>x"8a00", 816=>x"6200", 817=>x"6200", 818=>x"6200", 819=>x"6200",
---- 820=>x"6500", 821=>x"7200", 822=>x"7e00", 823=>x"8800", 824=>x"6500", 825=>x"6300", 826=>x"6100",
---- 827=>x"5f00", 828=>x"9d00", 829=>x"6d00", 830=>x"7c00", 831=>x"8900", 832=>x"6200", 833=>x"6500",
---- 834=>x"6200", 835=>x"5f00", 836=>x"6200", 837=>x"6c00", 838=>x"7800", 839=>x"8900", 840=>x"6500",
---- 841=>x"6300", 842=>x"5f00", 843=>x"5e00", 844=>x"5e00", 845=>x"6800", 846=>x"7c00", 847=>x"8800",
---- 848=>x"6500", 849=>x"6100", 850=>x"6100", 851=>x"5b00", 852=>x"5d00", 853=>x"6900", 854=>x"7900",
---- 855=>x"8700", 856=>x"6500", 857=>x"6400", 858=>x"5f00", 859=>x"5a00", 860=>x"5a00", 861=>x"6700",
---- 862=>x"7700", 863=>x"8600", 864=>x"6200", 865=>x"6200", 866=>x"5f00", 867=>x"5900", 868=>x"5c00",
---- 869=>x"6800", 870=>x"7900", 871=>x"8600", 872=>x"6300", 873=>x"6300", 874=>x"5e00", 875=>x"5900",
---- 876=>x"5900", 877=>x"6400", 878=>x"7800", 879=>x"8500", 880=>x"6200", 881=>x"6200", 882=>x"5f00",
---- 883=>x"5b00", 884=>x"5a00", 885=>x"6400", 886=>x"7700", 887=>x"8700", 888=>x"6500", 889=>x"6500",
---- 890=>x"6200", 891=>x"5c00", 892=>x"5c00", 893=>x"6900", 894=>x"7800", 895=>x"8500", 896=>x"6200",
---- 897=>x"6400", 898=>x"6200", 899=>x"5d00", 900=>x"5a00", 901=>x"6600", 902=>x"7700", 903=>x"8700",
---- 904=>x"6300", 905=>x"6000", 906=>x"5f00", 907=>x"5e00", 908=>x"5c00", 909=>x"6400", 910=>x"7500",
---- 911=>x"8800", 912=>x"6400", 913=>x"6200", 914=>x"6000", 915=>x"5e00", 916=>x"5a00", 917=>x"6600",
---- 918=>x"7700", 919=>x"8800", 920=>x"6200", 921=>x"6300", 922=>x"5f00", 923=>x"5b00", 924=>x"5e00",
---- 925=>x"6800", 926=>x"7600", 927=>x"8600", 928=>x"6200", 929=>x"6000", 930=>x"5c00", 931=>x"5c00",
---- 932=>x"5f00", 933=>x"6500", 934=>x"7300", 935=>x"8200", 936=>x"5e00", 937=>x"5c00", 938=>x"5d00",
---- 939=>x"5b00", 940=>x"5500", 941=>x"6200", 942=>x"8900", 943=>x"8300", 944=>x"6100", 945=>x"6000",
---- 946=>x"5c00", 947=>x"5c00", 948=>x"5800", 949=>x"6500", 950=>x"7800", 951=>x"8600", 952=>x"6200",
---- 953=>x"6300", 954=>x"6100", 955=>x"5b00", 956=>x"5b00", 957=>x"6400", 958=>x"7600", 959=>x"8500",
---- 960=>x"6000", 961=>x"6200", 962=>x"6200", 963=>x"5a00", 964=>x"5800", 965=>x"6400", 966=>x"7400",
---- 967=>x"8600", 968=>x"5e00", 969=>x"6100", 970=>x"5f00", 971=>x"5a00", 972=>x"5900", 973=>x"6400",
---- 974=>x"7300", 975=>x"8800", 976=>x"6100", 977=>x"6100", 978=>x"5f00", 979=>x"5e00", 980=>x"5800",
---- 981=>x"6300", 982=>x"7200", 983=>x"8700", 984=>x"6500", 985=>x"6300", 986=>x"5f00", 987=>x"5d00",
---- 988=>x"5c00", 989=>x"6100", 990=>x"7400", 991=>x"8500", 992=>x"6200", 993=>x"6400", 994=>x"6000",
---- 995=>x"5d00", 996=>x"5900", 997=>x"6000", 998=>x"7300", 999=>x"8500", 1000=>x"6500", 1001=>x"9d00",
---- 1002=>x"6100", 1003=>x"5e00", 1004=>x"5900", 1005=>x"6000", 1006=>x"7200", 1007=>x"8500", 1008=>x"6500",
---- 1009=>x"6300", 1010=>x"9c00", 1011=>x"5b00", 1012=>x"5900", 1013=>x"6000", 1014=>x"7100", 1015=>x"8200",
---- 1016=>x"6400", 1017=>x"6200", 1018=>x"5e00", 1019=>x"5700", 1020=>x"5600", 1021=>x"5f00", 1022=>x"7300",
---- 1023=>x"8300", 1024=>x"6500", 1025=>x"5f00", 1026=>x"5c00", 1027=>x"5500", 1028=>x"5500", 1029=>x"5f00",
---- 1030=>x"7300", 1031=>x"8400", 1032=>x"6300", 1033=>x"6000", 1034=>x"5c00", 1035=>x"5800", 1036=>x"5200",
---- 1037=>x"5b00", 1038=>x"7400", 1039=>x"8500", 1040=>x"5d00", 1041=>x"5f00", 1042=>x"5900", 1043=>x"5500",
---- 1044=>x"5200", 1045=>x"5700", 1046=>x"6f00", 1047=>x"8200", 1048=>x"5d00", 1049=>x"5b00", 1050=>x"5500",
---- 1051=>x"4e00", 1052=>x"4c00", 1053=>x"5500", 1054=>x"6a00", 1055=>x"7f00", 1056=>x"5a00", 1057=>x"5800",
---- 1058=>x"5300", 1059=>x"5300", 1060=>x"4a00", 1061=>x"5200", 1062=>x"6900", 1063=>x"8100", 1064=>x"5a00",
---- 1065=>x"5500", 1066=>x"5200", 1067=>x"4f00", 1068=>x"4800", 1069=>x"ac00", 1070=>x"6d00", 1071=>x"8300",
---- 1072=>x"5a00", 1073=>x"5700", 1074=>x"5600", 1075=>x"4f00", 1076=>x"4700", 1077=>x"5200", 1078=>x"6c00",
---- 1079=>x"8100", 1080=>x"5a00", 1081=>x"5a00", 1082=>x"5200", 1083=>x"4d00", 1084=>x"4600", 1085=>x"4f00",
---- 1086=>x"6800", 1087=>x"8000", 1088=>x"5900", 1089=>x"5a00", 1090=>x"5300", 1091=>x"4e00", 1092=>x"4600",
---- 1093=>x"5200", 1094=>x"6800", 1095=>x"7e00", 1096=>x"5b00", 1097=>x"5900", 1098=>x"5600", 1099=>x"4b00",
---- 1100=>x"4800", 1101=>x"4f00", 1102=>x"6900", 1103=>x"8100", 1104=>x"5b00", 1105=>x"5600", 1106=>x"5300",
---- 1107=>x"4e00", 1108=>x"4700", 1109=>x"4d00", 1110=>x"6900", 1111=>x"8000", 1112=>x"5800", 1113=>x"5600",
---- 1114=>x"4f00", 1115=>x"4e00", 1116=>x"4600", 1117=>x"4d00", 1118=>x"6600", 1119=>x"7f00", 1120=>x"5500",
---- 1121=>x"a900", 1122=>x"5200", 1123=>x"4a00", 1124=>x"4600", 1125=>x"4a00", 1126=>x"6400", 1127=>x"7e00",
---- 1128=>x"5400", 1129=>x"5300", 1130=>x"5100", 1131=>x"4b00", 1132=>x"4100", 1133=>x"4900", 1134=>x"6200",
---- 1135=>x"7b00", 1136=>x"5300", 1137=>x"5200", 1138=>x"4a00", 1139=>x"4300", 1140=>x"3800", 1141=>x"4000",
---- 1142=>x"6000", 1143=>x"7d00", 1144=>x"5100", 1145=>x"5200", 1146=>x"4900", 1147=>x"4200", 1148=>x"3c00",
---- 1149=>x"4100", 1150=>x"5a00", 1151=>x"7b00", 1152=>x"5100", 1153=>x"4f00", 1154=>x"4700", 1155=>x"4100",
---- 1156=>x"3c00", 1157=>x"4600", 1158=>x"5b00", 1159=>x"7a00", 1160=>x"4d00", 1161=>x"4c00", 1162=>x"4600",
---- 1163=>x"3e00", 1164=>x"3b00", 1165=>x"4300", 1166=>x"5900", 1167=>x"7700", 1168=>x"4c00", 1169=>x"4b00",
---- 1170=>x"4600", 1171=>x"3f00", 1172=>x"3900", 1173=>x"4200", 1174=>x"6000", 1175=>x"7900", 1176=>x"4c00",
---- 1177=>x"4900", 1178=>x"4600", 1179=>x"3f00", 1180=>x"3800", 1181=>x"4200", 1182=>x"5f00", 1183=>x"7900",
---- 1184=>x"4b00", 1185=>x"4700", 1186=>x"4300", 1187=>x"3d00", 1188=>x"3a00", 1189=>x"3e00", 1190=>x"5900",
---- 1191=>x"7900", 1192=>x"4900", 1193=>x"4a00", 1194=>x"4300", 1195=>x"4000", 1196=>x"3900", 1197=>x"3f00",
---- 1198=>x"5900", 1199=>x"7900", 1200=>x"4600", 1201=>x"4500", 1202=>x"4100", 1203=>x"3c00", 1204=>x"3700",
---- 1205=>x"4000", 1206=>x"5800", 1207=>x"7800", 1208=>x"4300", 1209=>x"4400", 1210=>x"4000", 1211=>x"3900",
---- 1212=>x"3500", 1213=>x"4100", 1214=>x"5400", 1215=>x"7600", 1216=>x"4500", 1217=>x"4400", 1218=>x"c100",
---- 1219=>x"3900", 1220=>x"3400", 1221=>x"3a00", 1222=>x"5700", 1223=>x"7700", 1224=>x"4600", 1225=>x"4200",
---- 1226=>x"3f00", 1227=>x"3500", 1228=>x"3100", 1229=>x"3d00", 1230=>x"5c00", 1231=>x"7800", 1232=>x"4100",
---- 1233=>x"4100", 1234=>x"3e00", 1235=>x"3500", 1236=>x"3200", 1237=>x"3c00", 1238=>x"5800", 1239=>x"7600",
---- 1240=>x"4300", 1241=>x"3f00", 1242=>x"3c00", 1243=>x"3700", 1244=>x"2f00", 1245=>x"3600", 1246=>x"5500",
---- 1247=>x"7900", 1248=>x"4400", 1249=>x"3f00", 1250=>x"3500", 1251=>x"3300", 1252=>x"2c00", 1253=>x"3100",
---- 1254=>x"5400", 1255=>x"7600", 1256=>x"4300", 1257=>x"3e00", 1258=>x"3600", 1259=>x"3100", 1260=>x"2c00",
---- 1261=>x"3000", 1262=>x"5400", 1263=>x"7400", 1264=>x"4000", 1265=>x"3900", 1266=>x"3700", 1267=>x"3100",
---- 1268=>x"2a00", 1269=>x"2f00", 1270=>x"4f00", 1271=>x"7300", 1272=>x"4200", 1273=>x"3e00", 1274=>x"3a00",
---- 1275=>x"3000", 1276=>x"2a00", 1277=>x"d000", 1278=>x"5200", 1279=>x"7600", 1280=>x"4500", 1281=>x"4100",
---- 1282=>x"3e00", 1283=>x"3300", 1284=>x"2900", 1285=>x"3800", 1286=>x"5900", 1287=>x"7500", 1288=>x"4200",
---- 1289=>x"4000", 1290=>x"3e00", 1291=>x"3900", 1292=>x"3000", 1293=>x"3e00", 1294=>x"5b00", 1295=>x"7800",
---- 1296=>x"4400", 1297=>x"4000", 1298=>x"4000", 1299=>x"c300", 1300=>x"3700", 1301=>x"4600", 1302=>x"6700",
---- 1303=>x"7e00", 1304=>x"4500", 1305=>x"4500", 1306=>x"4500", 1307=>x"4300", 1308=>x"4000", 1309=>x"4f00",
---- 1310=>x"9300", 1311=>x"8200", 1312=>x"4300", 1313=>x"4100", 1314=>x"4600", 1315=>x"4700", 1316=>x"4a00",
---- 1317=>x"5600", 1318=>x"7300", 1319=>x"8600", 1320=>x"4400", 1321=>x"4200", 1322=>x"4800", 1323=>x"4b00",
---- 1324=>x"4f00", 1325=>x"5a00", 1326=>x"7600", 1327=>x"8900", 1328=>x"4600", 1329=>x"4700", 1330=>x"4300",
---- 1331=>x"4a00", 1332=>x"5500", 1333=>x"6200", 1334=>x"7800", 1335=>x"8b00", 1336=>x"4900", 1337=>x"4100",
---- 1338=>x"3c00", 1339=>x"4400", 1340=>x"5700", 1341=>x"6600", 1342=>x"7800", 1343=>x"8b00", 1344=>x"4600",
---- 1345=>x"3d00", 1346=>x"3a00", 1347=>x"4400", 1348=>x"5400", 1349=>x"6600", 1350=>x"7f00", 1351=>x"8c00",
---- 1352=>x"4000", 1353=>x"3d00", 1354=>x"3c00", 1355=>x"4500", 1356=>x"5500", 1357=>x"6800", 1358=>x"7e00",
---- 1359=>x"8c00", 1360=>x"4100", 1361=>x"4100", 1362=>x"3f00", 1363=>x"4800", 1364=>x"5100", 1365=>x"6400",
---- 1366=>x"7b00", 1367=>x"8900", 1368=>x"4100", 1369=>x"3e00", 1370=>x"4200", 1371=>x"4b00", 1372=>x"5000",
---- 1373=>x"6000", 1374=>x"7700", 1375=>x"8600", 1376=>x"4000", 1377=>x"4000", 1378=>x"4500", 1379=>x"4300",
---- 1380=>x"4f00", 1381=>x"5f00", 1382=>x"7700", 1383=>x"8900", 1384=>x"4300", 1385=>x"3f00", 1386=>x"3f00",
---- 1387=>x"4800", 1388=>x"5100", 1389=>x"5e00", 1390=>x"7a00", 1391=>x"8900", 1392=>x"4200", 1393=>x"3c00",
---- 1394=>x"3d00", 1395=>x"b800", 1396=>x"4e00", 1397=>x"5a00", 1398=>x"7800", 1399=>x"8b00", 1400=>x"3e00",
---- 1401=>x"3d00", 1402=>x"4100", 1403=>x"4a00", 1404=>x"5000", 1405=>x"6100", 1406=>x"7700", 1407=>x"8d00",
---- 1408=>x"3f00", 1409=>x"4000", 1410=>x"4000", 1411=>x"5000", 1412=>x"5600", 1413=>x"6600", 1414=>x"7a00",
---- 1415=>x"8d00", 1416=>x"3c00", 1417=>x"3d00", 1418=>x"4600", 1419=>x"5700", 1420=>x"5b00", 1421=>x"6700",
---- 1422=>x"7e00", 1423=>x"8d00", 1424=>x"3d00", 1425=>x"3b00", 1426=>x"4900", 1427=>x"5100", 1428=>x"5b00",
---- 1429=>x"6600", 1430=>x"7b00", 1431=>x"8c00", 1432=>x"3b00", 1433=>x"3700", 1434=>x"4600", 1435=>x"5600",
---- 1436=>x"5b00", 1437=>x"6400", 1438=>x"7800", 1439=>x"8a00", 1440=>x"3700", 1441=>x"3800", 1442=>x"4600",
---- 1443=>x"ac00", 1444=>x"5b00", 1445=>x"5f00", 1446=>x"7600", 1447=>x"8a00", 1448=>x"3600", 1449=>x"3800",
---- 1450=>x"4700", 1451=>x"5500", 1452=>x"5d00", 1453=>x"5e00", 1454=>x"7200", 1455=>x"8900", 1456=>x"3500",
---- 1457=>x"3700", 1458=>x"4800", 1459=>x"5c00", 1460=>x"5800", 1461=>x"5700", 1462=>x"7200", 1463=>x"8600",
---- 1464=>x"3300", 1465=>x"3900", 1466=>x"5100", 1467=>x"6000", 1468=>x"5a00", 1469=>x"5800", 1470=>x"6e00",
---- 1471=>x"8400", 1472=>x"2e00", 1473=>x"3e00", 1474=>x"6200", 1475=>x"6400", 1476=>x"6100", 1477=>x"6300",
---- 1478=>x"7300", 1479=>x"8100", 1480=>x"2e00", 1481=>x"4500", 1482=>x"6400", 1483=>x"6900", 1484=>x"6500",
---- 1485=>x"6700", 1486=>x"7700", 1487=>x"8400", 1488=>x"3400", 1489=>x"4f00", 1490=>x"6500", 1491=>x"6600",
---- 1492=>x"6600", 1493=>x"6700", 1494=>x"7800", 1495=>x"8300", 1496=>x"3500", 1497=>x"4e00", 1498=>x"6500",
---- 1499=>x"6800", 1500=>x"6500", 1501=>x"6600", 1502=>x"7a00", 1503=>x"8400", 1504=>x"3500", 1505=>x"5300",
---- 1506=>x"6500", 1507=>x"6d00", 1508=>x"6700", 1509=>x"6400", 1510=>x"7800", 1511=>x"8500", 1512=>x"3900",
---- 1513=>x"5200", 1514=>x"5900", 1515=>x"6100", 1516=>x"5f00", 1517=>x"6500", 1518=>x"7700", 1519=>x"8500",
---- 1520=>x"3700", 1521=>x"4600", 1522=>x"5600", 1523=>x"5e00", 1524=>x"6200", 1525=>x"6900", 1526=>x"7c00",
---- 1527=>x"8800", 1528=>x"3100", 1529=>x"3c00", 1530=>x"5100", 1531=>x"5e00", 1532=>x"6500", 1533=>x"7000",
---- 1534=>x"8100", 1535=>x"8400", 1536=>x"3300", 1537=>x"3500", 1538=>x"4a00", 1539=>x"5e00", 1540=>x"9c00",
---- 1541=>x"6a00", 1542=>x"7a00", 1543=>x"8300", 1544=>x"2b00", 1545=>x"3800", 1546=>x"4500", 1547=>x"5c00",
---- 1548=>x"6000", 1549=>x"5c00", 1550=>x"7100", 1551=>x"8300", 1552=>x"2700", 1553=>x"3400", 1554=>x"4500",
---- 1555=>x"5700", 1556=>x"5d00", 1557=>x"5900", 1558=>x"6800", 1559=>x"7e00", 1560=>x"2a00", 1561=>x"3300",
---- 1562=>x"4500", 1563=>x"5000", 1564=>x"5200", 1565=>x"4d00", 1566=>x"6400", 1567=>x"7f00", 1568=>x"2500",
---- 1569=>x"3200", 1570=>x"3f00", 1571=>x"4900", 1572=>x"4d00", 1573=>x"4a00", 1574=>x"9e00", 1575=>x"8000",
---- 1576=>x"2800", 1577=>x"2f00", 1578=>x"3c00", 1579=>x"4700", 1580=>x"4800", 1581=>x"4700", 1582=>x"a300",
---- 1583=>x"7700", 1584=>x"2f00", 1585=>x"3500", 1586=>x"4300", 1587=>x"4200", 1588=>x"3b00", 1589=>x"3f00",
---- 1590=>x"5100", 1591=>x"6b00", 1592=>x"3300", 1593=>x"3d00", 1594=>x"3e00", 1595=>x"3900", 1596=>x"3600",
---- 1597=>x"3400", 1598=>x"4300", 1599=>x"5f00", 1600=>x"3b00", 1601=>x"4600", 1602=>x"3e00", 1603=>x"3700",
---- 1604=>x"3500", 1605=>x"cd00", 1606=>x"4000", 1607=>x"5600", 1608=>x"4700", 1609=>x"4d00", 1610=>x"4500",
---- 1611=>x"3800", 1612=>x"3500", 1613=>x"3100", 1614=>x"3e00", 1615=>x"5700", 1616=>x"5700", 1617=>x"5600",
---- 1618=>x"b100", 1619=>x"4200", 1620=>x"3200", 1621=>x"2d00", 1622=>x"3c00", 1623=>x"5700", 1624=>x"6400",
---- 1625=>x"5f00", 1626=>x"5500", 1627=>x"4800", 1628=>x"3200", 1629=>x"2b00", 1630=>x"3a00", 1631=>x"5500",
---- 1632=>x"7300", 1633=>x"6900", 1634=>x"5800", 1635=>x"4800", 1636=>x"3800", 1637=>x"2b00", 1638=>x"3500",
---- 1639=>x"5500", 1640=>x"8100", 1641=>x"7500", 1642=>x"6100", 1643=>x"4b00", 1644=>x"3c00", 1645=>x"2b00",
---- 1646=>x"3400", 1647=>x"5700", 1648=>x"8500", 1649=>x"8300", 1650=>x"7200", 1651=>x"5700", 1652=>x"4200",
---- 1653=>x"2b00", 1654=>x"3900", 1655=>x"5200", 1656=>x"9200", 1657=>x"9300", 1658=>x"7e00", 1659=>x"6200",
---- 1660=>x"4200", 1661=>x"2b00", 1662=>x"3800", 1663=>x"5600", 1664=>x"a100", 1665=>x"9900", 1666=>x"8500",
---- 1667=>x"6c00", 1668=>x"4300", 1669=>x"2b00", 1670=>x"3500", 1671=>x"5500", 1672=>x"a400", 1673=>x"9800",
---- 1674=>x"8a00", 1675=>x"7800", 1676=>x"5000", 1677=>x"2a00", 1678=>x"3300", 1679=>x"5200", 1680=>x"a700",
---- 1681=>x"9e00", 1682=>x"8e00", 1683=>x"7d00", 1684=>x"5800", 1685=>x"2c00", 1686=>x"3000", 1687=>x"5000",
---- 1688=>x"ab00", 1689=>x"a300", 1690=>x"9300", 1691=>x"8500", 1692=>x"5d00", 1693=>x"2c00", 1694=>x"2b00",
---- 1695=>x"4800", 1696=>x"ab00", 1697=>x"a400", 1698=>x"9a00", 1699=>x"8600", 1700=>x"6000", 1701=>x"2900",
---- 1702=>x"2500", 1703=>x"3f00", 1704=>x"aa00", 1705=>x"a900", 1706=>x"9c00", 1707=>x"8c00", 1708=>x"5700",
---- 1709=>x"2500", 1710=>x"2600", 1711=>x"4000", 1712=>x"af00", 1713=>x"a900", 1714=>x"a000", 1715=>x"8900",
---- 1716=>x"4f00", 1717=>x"2400", 1718=>x"2700", 1719=>x"4500", 1720=>x"ad00", 1721=>x"a800", 1722=>x"9900",
---- 1723=>x"8400", 1724=>x"5400", 1725=>x"2500", 1726=>x"2100", 1727=>x"4000", 1728=>x"aa00", 1729=>x"aa00",
---- 1730=>x"9c00", 1731=>x"8500", 1732=>x"5700", 1733=>x"2500", 1734=>x"2300", 1735=>x"3f00", 1736=>x"ad00",
---- 1737=>x"ac00", 1738=>x"a000", 1739=>x"8b00", 1740=>x"5600", 1741=>x"2300", 1742=>x"2500", 1743=>x"3b00",
---- 1744=>x"ae00", 1745=>x"aa00", 1746=>x"9e00", 1747=>x"8c00", 1748=>x"5e00", 1749=>x"2700", 1750=>x"2200",
---- 1751=>x"3800", 1752=>x"b100", 1753=>x"af00", 1754=>x"a000", 1755=>x"8d00", 1756=>x"9a00", 1757=>x"2c00",
---- 1758=>x"2300", 1759=>x"3800", 1760=>x"4f00", 1761=>x"ab00", 1762=>x"a000", 1763=>x"8c00", 1764=>x"6a00",
---- 1765=>x"3000", 1766=>x"2300", 1767=>x"3800", 1768=>x"ac00", 1769=>x"aa00", 1770=>x"a200", 1771=>x"8e00",
---- 1772=>x"7200", 1773=>x"3b00", 1774=>x"2400", 1775=>x"3b00", 1776=>x"ac00", 1777=>x"ac00", 1778=>x"a200",
---- 1779=>x"9100", 1780=>x"7500", 1781=>x"3700", 1782=>x"2300", 1783=>x"3700", 1784=>x"ad00", 1785=>x"ad00",
---- 1786=>x"a700", 1787=>x"9700", 1788=>x"7300", 1789=>x"3700", 1790=>x"2600", 1791=>x"3b00", 1792=>x"ac00",
---- 1793=>x"ac00", 1794=>x"a900", 1795=>x"9800", 1796=>x"7300", 1797=>x"3f00", 1798=>x"2500", 1799=>x"3b00",
---- 1800=>x"a800", 1801=>x"ad00", 1802=>x"a500", 1803=>x"9700", 1804=>x"7800", 1805=>x"3e00", 1806=>x"2a00",
---- 1807=>x"3e00", 1808=>x"a800", 1809=>x"ab00", 1810=>x"a400", 1811=>x"9900", 1812=>x"7a00", 1813=>x"4700",
---- 1814=>x"2e00", 1815=>x"3d00", 1816=>x"aa00", 1817=>x"ab00", 1818=>x"a700", 1819=>x"9700", 1820=>x"7e00",
---- 1821=>x"5100", 1822=>x"3100", 1823=>x"4000", 1824=>x"a400", 1825=>x"ab00", 1826=>x"a700", 1827=>x"9a00",
---- 1828=>x"8400", 1829=>x"5d00", 1830=>x"3900", 1831=>x"4000", 1832=>x"a200", 1833=>x"a600", 1834=>x"a300",
---- 1835=>x"9900", 1836=>x"8400", 1837=>x"6000", 1838=>x"3700", 1839=>x"3e00", 1840=>x"9f00", 1841=>x"a400",
---- 1842=>x"a300", 1843=>x"9700", 1844=>x"8400", 1845=>x"5e00", 1846=>x"3d00", 1847=>x"4000", 1848=>x"a200",
---- 1849=>x"ad00", 1850=>x"ac00", 1851=>x"a100", 1852=>x"8800", 1853=>x"5a00", 1854=>x"3d00", 1855=>x"4300",
---- 1856=>x"ad00", 1857=>x"af00", 1858=>x"af00", 1859=>x"a500", 1860=>x"9000", 1861=>x"6700", 1862=>x"3e00",
---- 1863=>x"3d00", 1864=>x"a800", 1865=>x"b000", 1866=>x"b000", 1867=>x"5700", 1868=>x"9200", 1869=>x"7300",
---- 1870=>x"c100", 1871=>x"3a00", 1872=>x"a700", 1873=>x"af00", 1874=>x"af00", 1875=>x"a900", 1876=>x"9500",
---- 1877=>x"7c00", 1878=>x"4700", 1879=>x"3c00", 1880=>x"a600", 1881=>x"af00", 1882=>x"b300", 1883=>x"aa00",
---- 1884=>x"9c00", 1885=>x"8300", 1886=>x"4c00", 1887=>x"3900", 1888=>x"a700", 1889=>x"b200", 1890=>x"b500",
---- 1891=>x"ac00", 1892=>x"a300", 1893=>x"8800", 1894=>x"4d00", 1895=>x"3d00", 1896=>x"aa00", 1897=>x"b200",
---- 1898=>x"b500", 1899=>x"b300", 1900=>x"ab00", 1901=>x"8600", 1902=>x"5200", 1903=>x"3e00", 1904=>x"a500",
---- 1905=>x"b400", 1906=>x"b900", 1907=>x"b600", 1908=>x"aa00", 1909=>x"8a00", 1910=>x"5d00", 1911=>x"4300",
---- 1912=>x"a400", 1913=>x"b200", 1914=>x"b800", 1915=>x"b400", 1916=>x"a800", 1917=>x"9100", 1918=>x"6600",
---- 1919=>x"4800", 1920=>x"a500", 1921=>x"b000", 1922=>x"b700", 1923=>x"b600", 1924=>x"ae00", 1925=>x"9600",
---- 1926=>x"7000", 1927=>x"4d00", 1928=>x"a600", 1929=>x"b000", 1930=>x"b500", 1931=>x"b700", 1932=>x"b000",
---- 1933=>x"9900", 1934=>x"7500", 1935=>x"4d00", 1936=>x"a800", 1937=>x"b200", 1938=>x"b400", 1939=>x"b000",
---- 1940=>x"aa00", 1941=>x"9800", 1942=>x"7800", 1943=>x"5000", 1944=>x"a300", 1945=>x"ad00", 1946=>x"b100",
---- 1947=>x"af00", 1948=>x"ab00", 1949=>x"9800", 1950=>x"7700", 1951=>x"5700", 1952=>x"9c00", 1953=>x"aa00",
---- 1954=>x"b000", 1955=>x"b000", 1956=>x"ab00", 1957=>x"9600", 1958=>x"7600", 1959=>x"5900", 1960=>x"9800",
---- 1961=>x"a800", 1962=>x"b200", 1963=>x"b400", 1964=>x"ae00", 1965=>x"9a00", 1966=>x"7d00", 1967=>x"5a00",
---- 1968=>x"9400", 1969=>x"aa00", 1970=>x"b000", 1971=>x"b000", 1972=>x"ab00", 1973=>x"9c00", 1974=>x"8200",
---- 1975=>x"6200", 1976=>x"8f00", 1977=>x"a400", 1978=>x"ac00", 1979=>x"ae00", 1980=>x"ab00", 1981=>x"9c00",
---- 1982=>x"8200", 1983=>x"9300", 1984=>x"8900", 1985=>x"a300", 1986=>x"ad00", 1987=>x"b200", 1988=>x"ad00",
---- 1989=>x"9b00", 1990=>x"8500", 1991=>x"7100", 1992=>x"8b00", 1993=>x"a600", 1994=>x"b600", 1995=>x"bc00",
---- 1996=>x"b800", 1997=>x"ab00", 1998=>x"8f00", 1999=>x"7600", 2000=>x"8d00", 2001=>x"b300", 2002=>x"c500",
---- 2003=>x"c900", 2004=>x"c600", 2005=>x"c200", 2006=>x"a500", 2007=>x"7900", 2008=>x"9200", 2009=>x"c100",
---- 2010=>x"ca00", 2011=>x"cc00", 2012=>x"c900", 2013=>x"c800", 2014=>x"4600", 2015=>x"8900", 2016=>x"9f00",
---- 2017=>x"c600", 2018=>x"c700", 2019=>x"cc00", 2020=>x"cb00", 2021=>x"c500", 2022=>x"be00", 2023=>x"9d00",
---- 2024=>x"a300", 2025=>x"c600", 2026=>x"c500", 2027=>x"ca00", 2028=>x"ca00", 2029=>x"c400", 2030=>x"bf00",
---- 2031=>x"a500", 2032=>x"9e00", 2033=>x"c600", 2034=>x"c500", 2035=>x"c700", 2036=>x"c600", 2037=>x"c300",
---- 2038=>x"4300", 2039=>x"a500", 2040=>x"9600", 2041=>x"c400", 2042=>x"c500", 2043=>x"3800", 2044=>x"c600",
---- 2045=>x"c100", 2046=>x"ba00", 2047=>x"9b00"),
---- 2  => (0=>x"9b00", 1=>x"9c00", 2=>x"a000", 3=>x"a400", 4=>x"a600", 5=>x"a700", 6=>x"ae00", 7=>x"ad00",
---- 8=>x"9b00", 9=>x"9c00", 10=>x"5d00", 11=>x"a400", 12=>x"a600", 13=>x"a700", 14=>x"ad00",
---- 15=>x"ad00", 16=>x"9c00", 17=>x"9b00", 18=>x"9f00", 19=>x"a300", 20=>x"a400", 21=>x"a700",
---- 22=>x"ac00", 23=>x"ad00", 24=>x"9d00", 25=>x"9900", 26=>x"9c00", 27=>x"a200", 28=>x"a600",
---- 29=>x"a900", 30=>x"ab00", 31=>x"ac00", 32=>x"9b00", 33=>x"9a00", 34=>x"a100", 35=>x"a400",
---- 36=>x"a800", 37=>x"ab00", 38=>x"ac00", 39=>x"ac00", 40=>x"9900", 41=>x"9d00", 42=>x"a100",
---- 43=>x"a600", 44=>x"a800", 45=>x"a800", 46=>x"ab00", 47=>x"ab00", 48=>x"9b00", 49=>x"a000",
---- 50=>x"a300", 51=>x"a600", 52=>x"a900", 53=>x"a900", 54=>x"a900", 55=>x"a800", 56=>x"9f00",
---- 57=>x"a300", 58=>x"a700", 59=>x"a800", 60=>x"a900", 61=>x"a800", 62=>x"a900", 63=>x"a800",
---- 64=>x"a200", 65=>x"a500", 66=>x"a800", 67=>x"a600", 68=>x"a700", 69=>x"a900", 70=>x"a500",
---- 71=>x"a700", 72=>x"a200", 73=>x"a700", 74=>x"a700", 75=>x"a600", 76=>x"a700", 77=>x"a400",
---- 78=>x"a600", 79=>x"a400", 80=>x"a400", 81=>x"a600", 82=>x"a400", 83=>x"a500", 84=>x"a700",
---- 85=>x"a400", 86=>x"a500", 87=>x"a200", 88=>x"a600", 89=>x"a600", 90=>x"a500", 91=>x"a200",
---- 92=>x"a600", 93=>x"a500", 94=>x"a400", 95=>x"a300", 96=>x"a700", 97=>x"a600", 98=>x"a800",
---- 99=>x"a500", 100=>x"5b00", 101=>x"a400", 102=>x"a300", 103=>x"9f00", 104=>x"a600", 105=>x"a700",
---- 106=>x"a600", 107=>x"5900", 108=>x"a100", 109=>x"a100", 110=>x"a100", 111=>x"9e00", 112=>x"a800",
---- 113=>x"a800", 114=>x"a600", 115=>x"a400", 116=>x"a000", 117=>x"9e00", 118=>x"9e00", 119=>x"9e00",
---- 120=>x"a900", 121=>x"a700", 122=>x"a600", 123=>x"a300", 124=>x"a000", 125=>x"9f00", 126=>x"9d00",
---- 127=>x"9d00", 128=>x"aa00", 129=>x"a700", 130=>x"a700", 131=>x"a200", 132=>x"9f00", 133=>x"9f00",
---- 134=>x"9e00", 135=>x"9e00", 136=>x"a700", 137=>x"a700", 138=>x"a900", 139=>x"a100", 140=>x"a000",
---- 141=>x"a100", 142=>x"9d00", 143=>x"9e00", 144=>x"a600", 145=>x"a600", 146=>x"a500", 147=>x"a000",
---- 148=>x"9c00", 149=>x"9e00", 150=>x"9e00", 151=>x"9f00", 152=>x"a500", 153=>x"a300", 154=>x"a200",
---- 155=>x"a100", 156=>x"9e00", 157=>x"9e00", 158=>x"a000", 159=>x"a100", 160=>x"a400", 161=>x"a300",
---- 162=>x"a000", 163=>x"a000", 164=>x"9f00", 165=>x"9f00", 166=>x"a100", 167=>x"a100", 168=>x"a000",
---- 169=>x"9c00", 170=>x"a000", 171=>x"a300", 172=>x"a000", 173=>x"9e00", 174=>x"a000", 175=>x"a000",
---- 176=>x"9c00", 177=>x"9c00", 178=>x"9d00", 179=>x"a200", 180=>x"a100", 181=>x"9f00", 182=>x"9f00",
---- 183=>x"9f00", 184=>x"9a00", 185=>x"9b00", 186=>x"a000", 187=>x"a400", 188=>x"a500", 189=>x"a300",
---- 190=>x"a000", 191=>x"a100", 192=>x"9500", 193=>x"9a00", 194=>x"a100", 195=>x"a200", 196=>x"a200",
---- 197=>x"a100", 198=>x"9f00", 199=>x"a100", 200=>x"9200", 201=>x"6500", 202=>x"a100", 203=>x"a600",
---- 204=>x"a300", 205=>x"a100", 206=>x"a100", 207=>x"a100", 208=>x"9000", 209=>x"9a00", 210=>x"a300",
---- 211=>x"a400", 212=>x"a400", 213=>x"a200", 214=>x"a200", 215=>x"a200", 216=>x"9100", 217=>x"9b00",
---- 218=>x"a200", 219=>x"a300", 220=>x"a400", 221=>x"a200", 222=>x"a200", 223=>x"5c00", 224=>x"9400",
---- 225=>x"9b00", 226=>x"a300", 227=>x"a600", 228=>x"a400", 229=>x"a300", 230=>x"a200", 231=>x"a600",
---- 232=>x"9700", 233=>x"9d00", 234=>x"a300", 235=>x"a400", 236=>x"a500", 237=>x"a600", 238=>x"a400",
---- 239=>x"a400", 240=>x"9700", 241=>x"9d00", 242=>x"a400", 243=>x"a800", 244=>x"a400", 245=>x"a700",
---- 246=>x"a400", 247=>x"a300", 248=>x"9800", 249=>x"9d00", 250=>x"a500", 251=>x"a800", 252=>x"a500",
---- 253=>x"a500", 254=>x"a600", 255=>x"a500", 256=>x"9900", 257=>x"9f00", 258=>x"a500", 259=>x"a700",
---- 260=>x"a600", 261=>x"a500", 262=>x"a400", 263=>x"a500", 264=>x"9900", 265=>x"a100", 266=>x"a600",
---- 267=>x"a600", 268=>x"a500", 269=>x"a600", 270=>x"a900", 271=>x"a300", 272=>x"9600", 273=>x"a200",
---- 274=>x"a400", 275=>x"a800", 276=>x"a700", 277=>x"a400", 278=>x"a500", 279=>x"a300", 280=>x"9400",
---- 281=>x"a000", 282=>x"a700", 283=>x"a600", 284=>x"a800", 285=>x"a400", 286=>x"a400", 287=>x"a600",
---- 288=>x"9600", 289=>x"9f00", 290=>x"a400", 291=>x"a800", 292=>x"ab00", 293=>x"a600", 294=>x"a600",
---- 295=>x"a500", 296=>x"9800", 297=>x"5f00", 298=>x"a600", 299=>x"a900", 300=>x"a700", 301=>x"a600",
---- 302=>x"5900", 303=>x"a400", 304=>x"9800", 305=>x"a000", 306=>x"a600", 307=>x"a700", 308=>x"a600",
---- 309=>x"a800", 310=>x"a700", 311=>x"a400", 312=>x"9700", 313=>x"9e00", 314=>x"a400", 315=>x"a800",
---- 316=>x"a800", 317=>x"a900", 318=>x"a800", 319=>x"a600", 320=>x"9700", 321=>x"9d00", 322=>x"a500",
---- 323=>x"a600", 324=>x"a800", 325=>x"a800", 326=>x"a700", 327=>x"a700", 328=>x"9700", 329=>x"9d00",
---- 330=>x"a400", 331=>x"a700", 332=>x"a700", 333=>x"a700", 334=>x"a900", 335=>x"a700", 336=>x"9700",
---- 337=>x"9c00", 338=>x"a300", 339=>x"a800", 340=>x"a800", 341=>x"a800", 342=>x"5700", 343=>x"a600",
---- 344=>x"9600", 345=>x"9f00", 346=>x"a500", 347=>x"a800", 348=>x"a700", 349=>x"a800", 350=>x"a700",
---- 351=>x"a600", 352=>x"9600", 353=>x"9f00", 354=>x"a400", 355=>x"a600", 356=>x"a800", 357=>x"a600",
---- 358=>x"a600", 359=>x"a500", 360=>x"9400", 361=>x"9b00", 362=>x"a200", 363=>x"a600", 364=>x"a700",
---- 365=>x"a800", 366=>x"a400", 367=>x"a600", 368=>x"9600", 369=>x"9c00", 370=>x"a200", 371=>x"a500",
---- 372=>x"a500", 373=>x"a800", 374=>x"a600", 375=>x"a400", 376=>x"9500", 377=>x"9c00", 378=>x"a000",
---- 379=>x"a400", 380=>x"a700", 381=>x"a700", 382=>x"a600", 383=>x"a600", 384=>x"9300", 385=>x"9b00",
---- 386=>x"a000", 387=>x"a500", 388=>x"a500", 389=>x"a700", 390=>x"a800", 391=>x"a700", 392=>x"9400",
---- 393=>x"9a00", 394=>x"a100", 395=>x"a400", 396=>x"a500", 397=>x"a700", 398=>x"a500", 399=>x"a600",
---- 400=>x"9300", 401=>x"9b00", 402=>x"a000", 403=>x"a300", 404=>x"a600", 405=>x"a600", 406=>x"a500",
---- 407=>x"a500", 408=>x"9300", 409=>x"9c00", 410=>x"a100", 411=>x"a700", 412=>x"a500", 413=>x"a500",
---- 414=>x"a800", 415=>x"a700", 416=>x"9300", 417=>x"9b00", 418=>x"9f00", 419=>x"a200", 420=>x"a600",
---- 421=>x"a600", 422=>x"a700", 423=>x"a600", 424=>x"9200", 425=>x"9b00", 426=>x"9f00", 427=>x"a400",
---- 428=>x"a400", 429=>x"a200", 430=>x"a400", 431=>x"a600", 432=>x"9400", 433=>x"9d00", 434=>x"9e00",
---- 435=>x"a200", 436=>x"a500", 437=>x"a300", 438=>x"a300", 439=>x"a300", 440=>x"9400", 441=>x"9c00",
---- 442=>x"a000", 443=>x"a200", 444=>x"a500", 445=>x"a500", 446=>x"a600", 447=>x"a300", 448=>x"9100",
---- 449=>x"9900", 450=>x"9f00", 451=>x"a400", 452=>x"a500", 453=>x"a500", 454=>x"a500", 455=>x"a400",
---- 456=>x"9500", 457=>x"9a00", 458=>x"9f00", 459=>x"a200", 460=>x"a500", 461=>x"a300", 462=>x"a300",
---- 463=>x"a200", 464=>x"9300", 465=>x"9c00", 466=>x"a000", 467=>x"a300", 468=>x"a600", 469=>x"a300",
---- 470=>x"a400", 471=>x"a400", 472=>x"9200", 473=>x"9b00", 474=>x"a000", 475=>x"a400", 476=>x"a300",
---- 477=>x"a500", 478=>x"a400", 479=>x"a200", 480=>x"9000", 481=>x"9b00", 482=>x"a000", 483=>x"a300",
---- 484=>x"a500", 485=>x"a400", 486=>x"a400", 487=>x"a300", 488=>x"9000", 489=>x"9900", 490=>x"a000",
---- 491=>x"a200", 492=>x"a500", 493=>x"a700", 494=>x"a700", 495=>x"a600", 496=>x"9300", 497=>x"9900",
---- 498=>x"9f00", 499=>x"a500", 500=>x"a600", 501=>x"a800", 502=>x"a600", 503=>x"a500", 504=>x"6c00",
---- 505=>x"9900", 506=>x"a000", 507=>x"a800", 508=>x"a900", 509=>x"a400", 510=>x"a800", 511=>x"a700",
---- 512=>x"9100", 513=>x"9900", 514=>x"a000", 515=>x"a400", 516=>x"a700", 517=>x"a700", 518=>x"a900",
---- 519=>x"a800", 520=>x"9000", 521=>x"9900", 522=>x"5e00", 523=>x"a700", 524=>x"a800", 525=>x"a800",
---- 526=>x"aa00", 527=>x"a800", 528=>x"9200", 529=>x"9900", 530=>x"9f00", 531=>x"a600", 532=>x"a600",
---- 533=>x"a500", 534=>x"a700", 535=>x"a800", 536=>x"9300", 537=>x"9a00", 538=>x"a000", 539=>x"a300",
---- 540=>x"a700", 541=>x"a600", 542=>x"a700", 543=>x"a600", 544=>x"9100", 545=>x"9900", 546=>x"9f00",
---- 547=>x"a400", 548=>x"a700", 549=>x"a600", 550=>x"a900", 551=>x"a800", 552=>x"9200", 553=>x"9800",
---- 554=>x"9b00", 555=>x"a400", 556=>x"a400", 557=>x"a700", 558=>x"aa00", 559=>x"aa00", 560=>x"9400",
---- 561=>x"9700", 562=>x"9e00", 563=>x"a600", 564=>x"a600", 565=>x"a900", 566=>x"a900", 567=>x"ac00",
---- 568=>x"9500", 569=>x"9c00", 570=>x"a100", 571=>x"a500", 572=>x"a700", 573=>x"ab00", 574=>x"ac00",
---- 575=>x"ad00", 576=>x"9300", 577=>x"9f00", 578=>x"a400", 579=>x"a500", 580=>x"a900", 581=>x"ab00",
---- 582=>x"ac00", 583=>x"ac00", 584=>x"9500", 585=>x"9b00", 586=>x"a100", 587=>x"a800", 588=>x"aa00",
---- 589=>x"ab00", 590=>x"5100", 591=>x"ad00", 592=>x"9400", 593=>x"9d00", 594=>x"a400", 595=>x"a900",
---- 596=>x"ab00", 597=>x"ac00", 598=>x"b000", 599=>x"b000", 600=>x"9400", 601=>x"9b00", 602=>x"a400",
---- 603=>x"ab00", 604=>x"ab00", 605=>x"ad00", 606=>x"af00", 607=>x"ae00", 608=>x"6a00", 609=>x"9b00",
---- 610=>x"a300", 611=>x"a800", 612=>x"ac00", 613=>x"ae00", 614=>x"ad00", 615=>x"ad00", 616=>x"9200",
---- 617=>x"9d00", 618=>x"a400", 619=>x"a800", 620=>x"ab00", 621=>x"ac00", 622=>x"ae00", 623=>x"ab00",
---- 624=>x"9400", 625=>x"9e00", 626=>x"a500", 627=>x"aa00", 628=>x"ad00", 629=>x"ac00", 630=>x"ad00",
---- 631=>x"ae00", 632=>x"9900", 633=>x"6100", 634=>x"a600", 635=>x"ab00", 636=>x"ab00", 637=>x"ad00",
---- 638=>x"ac00", 639=>x"ac00", 640=>x"9800", 641=>x"9e00", 642=>x"a400", 643=>x"aa00", 644=>x"ab00",
---- 645=>x"a900", 646=>x"ab00", 647=>x"ac00", 648=>x"9500", 649=>x"9e00", 650=>x"a400", 651=>x"a800",
---- 652=>x"aa00", 653=>x"ac00", 654=>x"ac00", 655=>x"ac00", 656=>x"9700", 657=>x"9f00", 658=>x"a400",
---- 659=>x"a900", 660=>x"ac00", 661=>x"aa00", 662=>x"ac00", 663=>x"ab00", 664=>x"9600", 665=>x"9f00",
---- 666=>x"a300", 667=>x"5500", 668=>x"a900", 669=>x"aa00", 670=>x"ab00", 671=>x"a800", 672=>x"9600",
---- 673=>x"6200", 674=>x"a400", 675=>x"a900", 676=>x"ab00", 677=>x"ad00", 678=>x"ae00", 679=>x"ad00",
---- 680=>x"9700", 681=>x"9f00", 682=>x"a400", 683=>x"a900", 684=>x"ac00", 685=>x"ac00", 686=>x"ab00",
---- 687=>x"ae00", 688=>x"9300", 689=>x"a000", 690=>x"a500", 691=>x"ab00", 692=>x"ab00", 693=>x"ac00",
---- 694=>x"ad00", 695=>x"ad00", 696=>x"9600", 697=>x"9e00", 698=>x"a500", 699=>x"ab00", 700=>x"a900",
---- 701=>x"ad00", 702=>x"ac00", 703=>x"ac00", 704=>x"9600", 705=>x"9f00", 706=>x"a500", 707=>x"ac00",
---- 708=>x"ac00", 709=>x"ad00", 710=>x"af00", 711=>x"af00", 712=>x"9700", 713=>x"9d00", 714=>x"a500",
---- 715=>x"ab00", 716=>x"ae00", 717=>x"ab00", 718=>x"ae00", 719=>x"af00", 720=>x"9900", 721=>x"9e00",
---- 722=>x"a600", 723=>x"ad00", 724=>x"ac00", 725=>x"ac00", 726=>x"ae00", 727=>x"af00", 728=>x"9800",
---- 729=>x"a100", 730=>x"a700", 731=>x"ab00", 732=>x"ac00", 733=>x"ad00", 734=>x"ac00", 735=>x"ad00",
---- 736=>x"9800", 737=>x"a000", 738=>x"a900", 739=>x"ac00", 740=>x"ac00", 741=>x"ab00", 742=>x"ad00",
---- 743=>x"ad00", 744=>x"9800", 745=>x"a000", 746=>x"a800", 747=>x"ac00", 748=>x"ac00", 749=>x"aa00",
---- 750=>x"ac00", 751=>x"ac00", 752=>x"9600", 753=>x"9d00", 754=>x"a600", 755=>x"a900", 756=>x"ac00",
---- 757=>x"ab00", 758=>x"aa00", 759=>x"b000", 760=>x"9600", 761=>x"9d00", 762=>x"a600", 763=>x"aa00",
---- 764=>x"ac00", 765=>x"ac00", 766=>x"ab00", 767=>x"ab00", 768=>x"9600", 769=>x"9d00", 770=>x"a400",
---- 771=>x"a900", 772=>x"ab00", 773=>x"aa00", 774=>x"aa00", 775=>x"aa00", 776=>x"9600", 777=>x"9d00",
---- 778=>x"a500", 779=>x"a800", 780=>x"a900", 781=>x"5400", 782=>x"aa00", 783=>x"ac00", 784=>x"9700",
---- 785=>x"9e00", 786=>x"a500", 787=>x"aa00", 788=>x"ad00", 789=>x"ac00", 790=>x"a900", 791=>x"ac00",
---- 792=>x"9500", 793=>x"9e00", 794=>x"a500", 795=>x"aa00", 796=>x"ac00", 797=>x"aa00", 798=>x"ad00",
---- 799=>x"ad00", 800=>x"9600", 801=>x"9e00", 802=>x"a600", 803=>x"aa00", 804=>x"ac00", 805=>x"aa00",
---- 806=>x"ac00", 807=>x"aa00", 808=>x"9600", 809=>x"a000", 810=>x"a800", 811=>x"ac00", 812=>x"ab00",
---- 813=>x"5400", 814=>x"ac00", 815=>x"ac00", 816=>x"9400", 817=>x"9f00", 818=>x"a500", 819=>x"aa00",
---- 820=>x"ac00", 821=>x"ab00", 822=>x"ac00", 823=>x"af00", 824=>x"9500", 825=>x"9d00", 826=>x"a500",
---- 827=>x"a700", 828=>x"ac00", 829=>x"ab00", 830=>x"ad00", 831=>x"ae00", 832=>x"9200", 833=>x"9e00",
---- 834=>x"a800", 835=>x"aa00", 836=>x"ab00", 837=>x"ad00", 838=>x"ad00", 839=>x"ac00", 840=>x"9400",
---- 841=>x"9f00", 842=>x"a400", 843=>x"5400", 844=>x"ae00", 845=>x"ac00", 846=>x"ad00", 847=>x"ad00",
---- 848=>x"9400", 849=>x"9c00", 850=>x"a200", 851=>x"a900", 852=>x"ad00", 853=>x"ae00", 854=>x"ad00",
---- 855=>x"ac00", 856=>x"9400", 857=>x"9900", 858=>x"a500", 859=>x"a900", 860=>x"ab00", 861=>x"ad00",
---- 862=>x"ab00", 863=>x"ab00", 864=>x"9000", 865=>x"9c00", 866=>x"a200", 867=>x"ab00", 868=>x"ae00",
---- 869=>x"ab00", 870=>x"ac00", 871=>x"af00", 872=>x"6d00", 873=>x"9a00", 874=>x"a400", 875=>x"a900",
---- 876=>x"aa00", 877=>x"5200", 878=>x"ad00", 879=>x"ae00", 880=>x"9200", 881=>x"9b00", 882=>x"a200",
---- 883=>x"aa00", 884=>x"ab00", 885=>x"ac00", 886=>x"ae00", 887=>x"ae00", 888=>x"9200", 889=>x"9b00",
---- 890=>x"a300", 891=>x"a900", 892=>x"ae00", 893=>x"ac00", 894=>x"aa00", 895=>x"af00", 896=>x"9200",
---- 897=>x"9b00", 898=>x"a200", 899=>x"a600", 900=>x"ab00", 901=>x"ad00", 902=>x"5200", 903=>x"ac00",
---- 904=>x"9400", 905=>x"9b00", 906=>x"a300", 907=>x"a700", 908=>x"ab00", 909=>x"af00", 910=>x"ad00",
---- 911=>x"ad00", 912=>x"9100", 913=>x"9b00", 914=>x"a400", 915=>x"a900", 916=>x"ac00", 917=>x"ac00",
---- 918=>x"ae00", 919=>x"af00", 920=>x"9100", 921=>x"9a00", 922=>x"a400", 923=>x"aa00", 924=>x"ab00",
---- 925=>x"ae00", 926=>x"ad00", 927=>x"5100", 928=>x"8f00", 929=>x"9800", 930=>x"a300", 931=>x"a800",
---- 932=>x"ab00", 933=>x"ad00", 934=>x"ae00", 935=>x"b000", 936=>x"9100", 937=>x"9b00", 938=>x"a400",
---- 939=>x"ab00", 940=>x"ad00", 941=>x"ae00", 942=>x"ae00", 943=>x"b000", 944=>x"9000", 945=>x"9800",
---- 946=>x"a100", 947=>x"5500", 948=>x"ac00", 949=>x"ad00", 950=>x"af00", 951=>x"ad00", 952=>x"9000",
---- 953=>x"9700", 954=>x"a500", 955=>x"ad00", 956=>x"ad00", 957=>x"ad00", 958=>x"b000", 959=>x"ad00",
---- 960=>x"9400", 961=>x"9d00", 962=>x"a400", 963=>x"aa00", 964=>x"aa00", 965=>x"ae00", 966=>x"b000",
---- 967=>x"af00", 968=>x"9300", 969=>x"9c00", 970=>x"a300", 971=>x"a900", 972=>x"ac00", 973=>x"ac00",
---- 974=>x"b000", 975=>x"af00", 976=>x"8f00", 977=>x"9a00", 978=>x"5c00", 979=>x"a900", 980=>x"ac00",
---- 981=>x"ae00", 982=>x"af00", 983=>x"af00", 984=>x"9000", 985=>x"9c00", 986=>x"a400", 987=>x"a800",
---- 988=>x"ad00", 989=>x"b000", 990=>x"b100", 991=>x"b200", 992=>x"9300", 993=>x"9c00", 994=>x"5d00",
---- 995=>x"a900", 996=>x"ad00", 997=>x"ad00", 998=>x"b100", 999=>x"b200", 1000=>x"9200", 1001=>x"9a00",
---- 1002=>x"a300", 1003=>x"ab00", 1004=>x"ae00", 1005=>x"ad00", 1006=>x"b000", 1007=>x"af00", 1008=>x"9100",
---- 1009=>x"9700", 1010=>x"a000", 1011=>x"aa00", 1012=>x"ae00", 1013=>x"ac00", 1014=>x"b000", 1015=>x"af00",
---- 1016=>x"9200", 1017=>x"9900", 1018=>x"a100", 1019=>x"ab00", 1020=>x"af00", 1021=>x"af00", 1022=>x"ae00",
---- 1023=>x"af00", 1024=>x"9100", 1025=>x"9a00", 1026=>x"a200", 1027=>x"ab00", 1028=>x"af00", 1029=>x"b100",
---- 1030=>x"af00", 1031=>x"b000", 1032=>x"9000", 1033=>x"9800", 1034=>x"a200", 1035=>x"aa00", 1036=>x"ae00",
---- 1037=>x"b000", 1038=>x"b000", 1039=>x"b300", 1040=>x"8f00", 1041=>x"9a00", 1042=>x"a400", 1043=>x"a900",
---- 1044=>x"ac00", 1045=>x"b100", 1046=>x"b000", 1047=>x"b100", 1048=>x"8f00", 1049=>x"9800", 1050=>x"a300",
---- 1051=>x"ab00", 1052=>x"ae00", 1053=>x"b000", 1054=>x"ae00", 1055=>x"b100", 1056=>x"8e00", 1057=>x"9800",
---- 1058=>x"a400", 1059=>x"ac00", 1060=>x"b000", 1061=>x"ae00", 1062=>x"b000", 1063=>x"b200", 1064=>x"8e00",
---- 1065=>x"9a00", 1066=>x"a400", 1067=>x"ad00", 1068=>x"b000", 1069=>x"b200", 1070=>x"af00", 1071=>x"b100",
---- 1072=>x"8d00", 1073=>x"9a00", 1074=>x"a400", 1075=>x"ac00", 1076=>x"b000", 1077=>x"b000", 1078=>x"b100",
---- 1079=>x"b200", 1080=>x"8d00", 1081=>x"9a00", 1082=>x"a400", 1083=>x"aa00", 1084=>x"b200", 1085=>x"b100",
---- 1086=>x"b100", 1087=>x"b600", 1088=>x"8f00", 1089=>x"9900", 1090=>x"a200", 1091=>x"ac00", 1092=>x"b100",
---- 1093=>x"b200", 1094=>x"b400", 1095=>x"b300", 1096=>x"9000", 1097=>x"9800", 1098=>x"a400", 1099=>x"aa00",
---- 1100=>x"b000", 1101=>x"b300", 1102=>x"b400", 1103=>x"b400", 1104=>x"8d00", 1105=>x"9b00", 1106=>x"a400",
---- 1107=>x"ab00", 1108=>x"af00", 1109=>x"b200", 1110=>x"b400", 1111=>x"b500", 1112=>x"6e00", 1113=>x"9c00",
---- 1114=>x"a300", 1115=>x"ab00", 1116=>x"ae00", 1117=>x"b100", 1118=>x"b300", 1119=>x"b600", 1120=>x"8e00",
---- 1121=>x"9900", 1122=>x"a300", 1123=>x"ab00", 1124=>x"b100", 1125=>x"b300", 1126=>x"b300", 1127=>x"b600",
---- 1128=>x"8c00", 1129=>x"9700", 1130=>x"a500", 1131=>x"ab00", 1132=>x"b000", 1133=>x"b200", 1134=>x"b300",
---- 1135=>x"b600", 1136=>x"8c00", 1137=>x"9800", 1138=>x"a200", 1139=>x"a900", 1140=>x"ae00", 1141=>x"4e00",
---- 1142=>x"b500", 1143=>x"b400", 1144=>x"8d00", 1145=>x"9700", 1146=>x"a100", 1147=>x"a900", 1148=>x"af00",
---- 1149=>x"b300", 1150=>x"b500", 1151=>x"b500", 1152=>x"8b00", 1153=>x"9600", 1154=>x"a100", 1155=>x"aa00",
---- 1156=>x"ad00", 1157=>x"b200", 1158=>x"b400", 1159=>x"b400", 1160=>x"8900", 1161=>x"9700", 1162=>x"a200",
---- 1163=>x"aa00", 1164=>x"af00", 1165=>x"b300", 1166=>x"b200", 1167=>x"b200", 1168=>x"8a00", 1169=>x"9700",
---- 1170=>x"a200", 1171=>x"a900", 1172=>x"af00", 1173=>x"b200", 1174=>x"b400", 1175=>x"b500", 1176=>x"8b00",
---- 1177=>x"9600", 1178=>x"a200", 1179=>x"aa00", 1180=>x"af00", 1181=>x"b000", 1182=>x"b200", 1183=>x"b300",
---- 1184=>x"8b00", 1185=>x"9800", 1186=>x"a200", 1187=>x"ab00", 1188=>x"af00", 1189=>x"b100", 1190=>x"b200",
---- 1191=>x"b300", 1192=>x"8800", 1193=>x"9700", 1194=>x"a100", 1195=>x"a800", 1196=>x"ae00", 1197=>x"b000",
---- 1198=>x"b200", 1199=>x"b400", 1200=>x"8a00", 1201=>x"9600", 1202=>x"5f00", 1203=>x"a900", 1204=>x"ac00",
---- 1205=>x"ae00", 1206=>x"b200", 1207=>x"b100", 1208=>x"8c00", 1209=>x"9600", 1210=>x"9f00", 1211=>x"a800",
---- 1212=>x"ab00", 1213=>x"ae00", 1214=>x"b000", 1215=>x"ae00", 1216=>x"8c00", 1217=>x"9900", 1218=>x"9f00",
---- 1219=>x"a800", 1220=>x"ad00", 1221=>x"af00", 1222=>x"ac00", 1223=>x"ac00", 1224=>x"8a00", 1225=>x"9500",
---- 1226=>x"9f00", 1227=>x"a500", 1228=>x"ac00", 1229=>x"ae00", 1230=>x"ac00", 1231=>x"ac00", 1232=>x"8900",
---- 1233=>x"9400", 1234=>x"9f00", 1235=>x"a600", 1236=>x"ac00", 1237=>x"ae00", 1238=>x"ac00", 1239=>x"ac00",
---- 1240=>x"8900", 1241=>x"9600", 1242=>x"9f00", 1243=>x"a700", 1244=>x"ab00", 1245=>x"ad00", 1246=>x"ad00",
---- 1247=>x"ab00", 1248=>x"8700", 1249=>x"9600", 1250=>x"a000", 1251=>x"a700", 1252=>x"ab00", 1253=>x"ad00",
---- 1254=>x"af00", 1255=>x"4f00", 1256=>x"8600", 1257=>x"9700", 1258=>x"9f00", 1259=>x"a700", 1260=>x"ab00",
---- 1261=>x"ad00", 1262=>x"b000", 1263=>x"b000", 1264=>x"8400", 1265=>x"9500", 1266=>x"a000", 1267=>x"a800",
---- 1268=>x"ac00", 1269=>x"ae00", 1270=>x"af00", 1271=>x"af00", 1272=>x"8600", 1273=>x"9600", 1274=>x"a100",
---- 1275=>x"a800", 1276=>x"ac00", 1277=>x"ae00", 1278=>x"af00", 1279=>x"b000", 1280=>x"8600", 1281=>x"9400",
---- 1282=>x"a200", 1283=>x"a900", 1284=>x"ad00", 1285=>x"ac00", 1286=>x"ae00", 1287=>x"ad00", 1288=>x"7500",
---- 1289=>x"6b00", 1290=>x"a100", 1291=>x"a800", 1292=>x"a900", 1293=>x"ac00", 1294=>x"ad00", 1295=>x"ae00",
---- 1296=>x"8e00", 1297=>x"9700", 1298=>x"9f00", 1299=>x"a600", 1300=>x"aa00", 1301=>x"ad00", 1302=>x"af00",
---- 1303=>x"af00", 1304=>x"9300", 1305=>x"9a00", 1306=>x"a200", 1307=>x"a800", 1308=>x"ab00", 1309=>x"ae00",
---- 1310=>x"ac00", 1311=>x"ae00", 1312=>x"9200", 1313=>x"9b00", 1314=>x"a300", 1315=>x"a500", 1316=>x"aa00",
---- 1317=>x"ab00", 1318=>x"ab00", 1319=>x"ad00", 1320=>x"9400", 1321=>x"9d00", 1322=>x"a300", 1323=>x"a700",
---- 1324=>x"a800", 1325=>x"aa00", 1326=>x"aa00", 1327=>x"ab00", 1328=>x"9800", 1329=>x"9c00", 1330=>x"a100",
---- 1331=>x"a800", 1332=>x"a700", 1333=>x"a900", 1334=>x"ab00", 1335=>x"ad00", 1336=>x"9700", 1337=>x"9d00",
---- 1338=>x"a200", 1339=>x"a600", 1340=>x"a700", 1341=>x"a900", 1342=>x"ab00", 1343=>x"b000", 1344=>x"9700",
---- 1345=>x"9e00", 1346=>x"a300", 1347=>x"a700", 1348=>x"a700", 1349=>x"ac00", 1350=>x"ab00", 1351=>x"ac00",
---- 1352=>x"9700", 1353=>x"9d00", 1354=>x"a400", 1355=>x"a700", 1356=>x"aa00", 1357=>x"a900", 1358=>x"a900",
---- 1359=>x"ac00", 1360=>x"9600", 1361=>x"9e00", 1362=>x"a300", 1363=>x"a500", 1364=>x"a800", 1365=>x"ab00",
---- 1366=>x"ab00", 1367=>x"af00", 1368=>x"9500", 1369=>x"9d00", 1370=>x"a200", 1371=>x"a600", 1372=>x"a800",
---- 1373=>x"5500", 1374=>x"ac00", 1375=>x"af00", 1376=>x"9500", 1377=>x"9b00", 1378=>x"a200", 1379=>x"a800",
---- 1380=>x"a900", 1381=>x"ab00", 1382=>x"ad00", 1383=>x"b000", 1384=>x"9700", 1385=>x"9f00", 1386=>x"a300",
---- 1387=>x"a700", 1388=>x"ab00", 1389=>x"ac00", 1390=>x"ac00", 1391=>x"ae00", 1392=>x"9700", 1393=>x"a100",
---- 1394=>x"a600", 1395=>x"a900", 1396=>x"ad00", 1397=>x"ad00", 1398=>x"ae00", 1399=>x"af00", 1400=>x"9800",
---- 1401=>x"9d00", 1402=>x"a400", 1403=>x"ad00", 1404=>x"af00", 1405=>x"ad00", 1406=>x"b000", 1407=>x"b200",
---- 1408=>x"9700", 1409=>x"9e00", 1410=>x"a500", 1411=>x"ac00", 1412=>x"af00", 1413=>x"b000", 1414=>x"b200",
---- 1415=>x"b100", 1416=>x"9700", 1417=>x"9f00", 1418=>x"a600", 1419=>x"ab00", 1420=>x"b000", 1421=>x"af00",
---- 1422=>x"b000", 1423=>x"af00", 1424=>x"9700", 1425=>x"9e00", 1426=>x"a300", 1427=>x"ab00", 1428=>x"af00",
---- 1429=>x"b000", 1430=>x"b200", 1431=>x"b200", 1432=>x"9700", 1433=>x"9c00", 1434=>x"a200", 1435=>x"aa00",
---- 1436=>x"ae00", 1437=>x"b000", 1438=>x"b200", 1439=>x"b000", 1440=>x"9600", 1441=>x"9e00", 1442=>x"a200",
---- 1443=>x"aa00", 1444=>x"ad00", 1445=>x"b100", 1446=>x"b200", 1447=>x"b300", 1448=>x"9300", 1449=>x"9e00",
---- 1450=>x"a200", 1451=>x"a800", 1452=>x"af00", 1453=>x"b200", 1454=>x"b300", 1455=>x"b300", 1456=>x"9100",
---- 1457=>x"9900", 1458=>x"a000", 1459=>x"a700", 1460=>x"b000", 1461=>x"b300", 1462=>x"b300", 1463=>x"b300",
---- 1464=>x"9000", 1465=>x"9600", 1466=>x"9d00", 1467=>x"a700", 1468=>x"af00", 1469=>x"b300", 1470=>x"b200",
---- 1471=>x"b200", 1472=>x"8c00", 1473=>x"9400", 1474=>x"9c00", 1475=>x"a600", 1476=>x"ae00", 1477=>x"af00",
---- 1478=>x"b200", 1479=>x"b100", 1480=>x"8a00", 1481=>x"9200", 1482=>x"9a00", 1483=>x"a500", 1484=>x"af00",
---- 1485=>x"b000", 1486=>x"b100", 1487=>x"b100", 1488=>x"8d00", 1489=>x"9200", 1490=>x"9a00", 1491=>x"a800",
---- 1492=>x"ad00", 1493=>x"af00", 1494=>x"b200", 1495=>x"b000", 1496=>x"8a00", 1497=>x"9500", 1498=>x"9c00",
---- 1499=>x"a500", 1500=>x"ae00", 1501=>x"af00", 1502=>x"b000", 1503=>x"b000", 1504=>x"8a00", 1505=>x"9300",
---- 1506=>x"9e00", 1507=>x"a600", 1508=>x"af00", 1509=>x"b000", 1510=>x"af00", 1511=>x"b000", 1512=>x"8a00",
---- 1513=>x"9300", 1514=>x"9c00", 1515=>x"a700", 1516=>x"ae00", 1517=>x"b000", 1518=>x"af00", 1519=>x"af00",
---- 1520=>x"8b00", 1521=>x"9500", 1522=>x"9f00", 1523=>x"a800", 1524=>x"ac00", 1525=>x"af00", 1526=>x"ad00",
---- 1527=>x"af00", 1528=>x"8b00", 1529=>x"9600", 1530=>x"9e00", 1531=>x"a700", 1532=>x"ad00", 1533=>x"ae00",
---- 1534=>x"ac00", 1535=>x"af00", 1536=>x"8f00", 1537=>x"9900", 1538=>x"a000", 1539=>x"a600", 1540=>x"ac00",
---- 1541=>x"ad00", 1542=>x"ac00", 1543=>x"ae00", 1544=>x"8d00", 1545=>x"9900", 1546=>x"a000", 1547=>x"a600",
---- 1548=>x"ad00", 1549=>x"ac00", 1550=>x"ad00", 1551=>x"ad00", 1552=>x"8b00", 1553=>x"9600", 1554=>x"a000",
---- 1555=>x"a600", 1556=>x"ab00", 1557=>x"ae00", 1558=>x"ac00", 1559=>x"ac00", 1560=>x"8c00", 1561=>x"9600",
---- 1562=>x"9e00", 1563=>x"a600", 1564=>x"ab00", 1565=>x"ad00", 1566=>x"ad00", 1567=>x"ad00", 1568=>x"8900",
---- 1569=>x"9400", 1570=>x"9d00", 1571=>x"a800", 1572=>x"ab00", 1573=>x"ad00", 1574=>x"ac00", 1575=>x"ae00",
---- 1576=>x"8500", 1577=>x"8f00", 1578=>x"9c00", 1579=>x"a400", 1580=>x"aa00", 1581=>x"ac00", 1582=>x"ab00",
---- 1583=>x"aa00", 1584=>x"7e00", 1585=>x"8d00", 1586=>x"9c00", 1587=>x"a500", 1588=>x"ab00", 1589=>x"ab00",
---- 1590=>x"aa00", 1591=>x"a900", 1592=>x"7700", 1593=>x"8900", 1594=>x"9a00", 1595=>x"a400", 1596=>x"aa00",
---- 1597=>x"a900", 1598=>x"ac00", 1599=>x"aa00", 1600=>x"7100", 1601=>x"8700", 1602=>x"9800", 1603=>x"a300",
---- 1604=>x"aa00", 1605=>x"a900", 1606=>x"ad00", 1607=>x"ad00", 1608=>x"7100", 1609=>x"8900", 1610=>x"9900",
---- 1611=>x"a200", 1612=>x"a800", 1613=>x"aa00", 1614=>x"a900", 1615=>x"ac00", 1616=>x"6f00", 1617=>x"8500",
---- 1618=>x"9a00", 1619=>x"a300", 1620=>x"a700", 1621=>x"a800", 1622=>x"5400", 1623=>x"aa00", 1624=>x"7200",
---- 1625=>x"8800", 1626=>x"9900", 1627=>x"a400", 1628=>x"a800", 1629=>x"a900", 1630=>x"ab00", 1631=>x"aa00",
---- 1632=>x"7500", 1633=>x"8a00", 1634=>x"9900", 1635=>x"a700", 1636=>x"5600", 1637=>x"ad00", 1638=>x"ad00",
---- 1639=>x"ab00", 1640=>x"7000", 1641=>x"8800", 1642=>x"9b00", 1643=>x"a500", 1644=>x"ac00", 1645=>x"ae00",
---- 1646=>x"ae00", 1647=>x"ad00", 1648=>x"6f00", 1649=>x"8800", 1650=>x"6500", 1651=>x"a400", 1652=>x"ab00",
---- 1653=>x"b100", 1654=>x"af00", 1655=>x"ad00", 1656=>x"7000", 1657=>x"8900", 1658=>x"9900", 1659=>x"a500",
---- 1660=>x"ae00", 1661=>x"b100", 1662=>x"b000", 1663=>x"af00", 1664=>x"7100", 1665=>x"8a00", 1666=>x"9d00",
---- 1667=>x"a600", 1668=>x"ae00", 1669=>x"b100", 1670=>x"b100", 1671=>x"b000", 1672=>x"7100", 1673=>x"8c00",
---- 1674=>x"9c00", 1675=>x"a500", 1676=>x"af00", 1677=>x"b300", 1678=>x"b000", 1679=>x"af00", 1680=>x"7200",
---- 1681=>x"8d00", 1682=>x"9c00", 1683=>x"a600", 1684=>x"ae00", 1685=>x"b200", 1686=>x"b200", 1687=>x"b200",
---- 1688=>x"7100", 1689=>x"8e00", 1690=>x"9c00", 1691=>x"a600", 1692=>x"b000", 1693=>x"af00", 1694=>x"b000",
---- 1695=>x"b000", 1696=>x"6f00", 1697=>x"8c00", 1698=>x"9a00", 1699=>x"a500", 1700=>x"ad00", 1701=>x"b100",
---- 1702=>x"b100", 1703=>x"ae00", 1704=>x"7000", 1705=>x"8d00", 1706=>x"9a00", 1707=>x"a500", 1708=>x"ae00",
---- 1709=>x"b300", 1710=>x"b300", 1711=>x"b000", 1712=>x"6f00", 1713=>x"8e00", 1714=>x"9a00", 1715=>x"a500",
---- 1716=>x"b000", 1717=>x"b500", 1718=>x"b400", 1719=>x"b200", 1720=>x"6f00", 1721=>x"8b00", 1722=>x"9a00",
---- 1723=>x"a800", 1724=>x"b000", 1725=>x"b200", 1726=>x"b100", 1727=>x"b000", 1728=>x"6c00", 1729=>x"8a00",
---- 1730=>x"9c00", 1731=>x"a700", 1732=>x"af00", 1733=>x"b300", 1734=>x"b100", 1735=>x"b300", 1736=>x"6b00",
---- 1737=>x"8b00", 1738=>x"9d00", 1739=>x"a800", 1740=>x"af00", 1741=>x"b400", 1742=>x"b300", 1743=>x"b200",
---- 1744=>x"6c00", 1745=>x"8a00", 1746=>x"9c00", 1747=>x"a800", 1748=>x"b300", 1749=>x"b500", 1750=>x"b300",
---- 1751=>x"b100", 1752=>x"6700", 1753=>x"8900", 1754=>x"9a00", 1755=>x"a700", 1756=>x"af00", 1757=>x"b200",
---- 1758=>x"b300", 1759=>x"b100", 1760=>x"6400", 1761=>x"8a00", 1762=>x"9d00", 1763=>x"a800", 1764=>x"b000",
---- 1765=>x"b100", 1766=>x"b100", 1767=>x"b100", 1768=>x"6300", 1769=>x"8800", 1770=>x"9b00", 1771=>x"a800",
---- 1772=>x"af00", 1773=>x"b000", 1774=>x"ad00", 1775=>x"ac00", 1776=>x"5f00", 1777=>x"8500", 1778=>x"9c00",
---- 1779=>x"a700", 1780=>x"b000", 1781=>x"b300", 1782=>x"b000", 1783=>x"af00", 1784=>x"6300", 1785=>x"8600",
---- 1786=>x"9b00", 1787=>x"a800", 1788=>x"af00", 1789=>x"b000", 1790=>x"b100", 1791=>x"b100", 1792=>x"9e00",
---- 1793=>x"8500", 1794=>x"9800", 1795=>x"a700", 1796=>x"ae00", 1797=>x"4d00", 1798=>x"b200", 1799=>x"b100",
---- 1800=>x"6100", 1801=>x"8500", 1802=>x"9600", 1803=>x"a600", 1804=>x"ae00", 1805=>x"b100", 1806=>x"b200",
---- 1807=>x"b100", 1808=>x"5d00", 1809=>x"8400", 1810=>x"9800", 1811=>x"a300", 1812=>x"ac00", 1813=>x"b000",
---- 1814=>x"b100", 1815=>x"b100", 1816=>x"5e00", 1817=>x"8400", 1818=>x"9600", 1819=>x"a500", 1820=>x"ae00",
---- 1821=>x"b100", 1822=>x"b100", 1823=>x"b100", 1824=>x"5d00", 1825=>x"8300", 1826=>x"9600", 1827=>x"a600",
---- 1828=>x"ad00", 1829=>x"b100", 1830=>x"b000", 1831=>x"af00", 1832=>x"5c00", 1833=>x"8000", 1834=>x"9500",
---- 1835=>x"a200", 1836=>x"aa00", 1837=>x"b100", 1838=>x"af00", 1839=>x"ad00", 1840=>x"5b00", 1841=>x"7e00",
---- 1842=>x"9200", 1843=>x"a000", 1844=>x"a900", 1845=>x"af00", 1846=>x"b000", 1847=>x"b000", 1848=>x"5c00",
---- 1849=>x"7e00", 1850=>x"9500", 1851=>x"a100", 1852=>x"aa00", 1853=>x"ac00", 1854=>x"af00", 1855=>x"af00",
---- 1856=>x"5500", 1857=>x"7d00", 1858=>x"9100", 1859=>x"9e00", 1860=>x"a800", 1861=>x"ab00", 1862=>x"ae00",
---- 1863=>x"ae00", 1864=>x"5800", 1865=>x"7b00", 1866=>x"8e00", 1867=>x"9e00", 1868=>x"a700", 1869=>x"ad00",
---- 1870=>x"ae00", 1871=>x"af00", 1872=>x"5700", 1873=>x"7800", 1874=>x"8f00", 1875=>x"9e00", 1876=>x"a700",
---- 1877=>x"ac00", 1878=>x"ad00", 1879=>x"af00", 1880=>x"5500", 1881=>x"7600", 1882=>x"9000", 1883=>x"9f00",
---- 1884=>x"a600", 1885=>x"ab00", 1886=>x"ae00", 1887=>x"b100", 1888=>x"5900", 1889=>x"7a00", 1890=>x"9200",
---- 1891=>x"9f00", 1892=>x"a700", 1893=>x"ac00", 1894=>x"b000", 1895=>x"af00", 1896=>x"5a00", 1897=>x"7700",
---- 1898=>x"8f00", 1899=>x"9d00", 1900=>x"a500", 1901=>x"ab00", 1902=>x"b000", 1903=>x"b000", 1904=>x"5900",
---- 1905=>x"7600", 1906=>x"8e00", 1907=>x"9d00", 1908=>x"a600", 1909=>x"ae00", 1910=>x"b100", 1911=>x"b100",
---- 1912=>x"5b00", 1913=>x"8a00", 1914=>x"8e00", 1915=>x"9d00", 1916=>x"a700", 1917=>x"ad00", 1918=>x"b000",
---- 1919=>x"b100", 1920=>x"5e00", 1921=>x"7300", 1922=>x"8d00", 1923=>x"9c00", 1924=>x"a800", 1925=>x"ad00",
---- 1926=>x"b100", 1927=>x"b400", 1928=>x"5c00", 1929=>x"7400", 1930=>x"8a00", 1931=>x"9d00", 1932=>x"a800",
---- 1933=>x"ac00", 1934=>x"b000", 1935=>x"b200", 1936=>x"5c00", 1937=>x"7500", 1938=>x"8b00", 1939=>x"9c00",
---- 1940=>x"a600", 1941=>x"ab00", 1942=>x"b000", 1943=>x"b000", 1944=>x"5c00", 1945=>x"7500", 1946=>x"8c00",
---- 1947=>x"9b00", 1948=>x"a700", 1949=>x"ad00", 1950=>x"ad00", 1951=>x"af00", 1952=>x"6000", 1953=>x"7100",
---- 1954=>x"8b00", 1955=>x"9a00", 1956=>x"a600", 1957=>x"ad00", 1958=>x"af00", 1959=>x"b100", 1960=>x"5c00",
---- 1961=>x"7200", 1962=>x"8800", 1963=>x"9900", 1964=>x"a500", 1965=>x"ae00", 1966=>x"b200", 1967=>x"b200",
---- 1968=>x"5d00", 1969=>x"7100", 1970=>x"8800", 1971=>x"9900", 1972=>x"a300", 1973=>x"ab00", 1974=>x"b000",
---- 1975=>x"b200", 1976=>x"6100", 1977=>x"7300", 1978=>x"8500", 1979=>x"9700", 1980=>x"a500", 1981=>x"ad00",
---- 1982=>x"b000", 1983=>x"b300", 1984=>x"6300", 1985=>x"7300", 1986=>x"8300", 1987=>x"9600", 1988=>x"a400",
---- 1989=>x"ac00", 1990=>x"b000", 1991=>x"b300", 1992=>x"6400", 1993=>x"7100", 1994=>x"8600", 1995=>x"9800",
---- 1996=>x"a500", 1997=>x"ae00", 1998=>x"4d00", 1999=>x"b300", 2000=>x"6600", 2001=>x"7600", 2002=>x"8700",
---- 2003=>x"9a00", 2004=>x"a500", 2005=>x"ae00", 2006=>x"b200", 2007=>x"b200", 2008=>x"6900", 2009=>x"7700",
---- 2010=>x"8500", 2011=>x"9800", 2012=>x"a400", 2013=>x"ad00", 2014=>x"b300", 2015=>x"b200", 2016=>x"6a00",
---- 2017=>x"7500", 2018=>x"8500", 2019=>x"9700", 2020=>x"a200", 2021=>x"ad00", 2022=>x"af00", 2023=>x"b000",
---- 2024=>x"6c00", 2025=>x"7400", 2026=>x"8600", 2027=>x"9800", 2028=>x"a200", 2029=>x"ae00", 2030=>x"b300",
---- 2031=>x"b000", 2032=>x"6e00", 2033=>x"7300", 2034=>x"8800", 2035=>x"9a00", 2036=>x"a300", 2037=>x"ac00",
---- 2038=>x"b200", 2039=>x"b200", 2040=>x"6a00", 2041=>x"7800", 2042=>x"8900", 2043=>x"9900", 2044=>x"a200",
---- 2045=>x"a900", 2046=>x"b200", 2047=>x"b400"),
---- 3  => (0=>x"ab00", 1=>x"ab00", 2=>x"a900", 3=>x"a200", 4=>x"9700", 5=>x"9600", 6=>x"8200", 7=>x"7300",
---- 8=>x"5400", 9=>x"ab00", 10=>x"a900", 11=>x"a300", 12=>x"9700", 13=>x"9700", 14=>x"8300",
---- 15=>x"7200", 16=>x"ab00", 17=>x"ac00", 18=>x"a900", 19=>x"a200", 20=>x"9800", 21=>x"9500",
---- 22=>x"8000", 23=>x"7000", 24=>x"ad00", 25=>x"ab00", 26=>x"a600", 27=>x"a000", 28=>x"9700",
---- 29=>x"8b00", 30=>x"7c00", 31=>x"7100", 32=>x"ac00", 33=>x"a900", 34=>x"a600", 35=>x"9e00",
---- 36=>x"9500", 37=>x"8b00", 38=>x"7d00", 39=>x"7300", 40=>x"aa00", 41=>x"a900", 42=>x"a700",
---- 43=>x"9d00", 44=>x"9100", 45=>x"8800", 46=>x"8000", 47=>x"7000", 48=>x"a800", 49=>x"a700",
---- 50=>x"a600", 51=>x"9d00", 52=>x"8e00", 53=>x"8900", 54=>x"7d00", 55=>x"6c00", 56=>x"a700",
---- 57=>x"a500", 58=>x"9f00", 59=>x"9b00", 60=>x"9300", 61=>x"8800", 62=>x"7d00", 63=>x"7200",
---- 64=>x"a600", 65=>x"a300", 66=>x"9f00", 67=>x"9b00", 68=>x"9000", 69=>x"8800", 70=>x"7c00",
---- 71=>x"6d00", 72=>x"a500", 73=>x"a300", 74=>x"9e00", 75=>x"9800", 76=>x"9000", 77=>x"8a00",
---- 78=>x"7f00", 79=>x"6f00", 80=>x"a200", 81=>x"a300", 82=>x"9d00", 83=>x"9a00", 84=>x"9100",
---- 85=>x"8b00", 86=>x"8400", 87=>x"7900", 88=>x"9f00", 89=>x"a100", 90=>x"9f00", 91=>x"9a00",
---- 92=>x"9300", 93=>x"8900", 94=>x"8200", 95=>x"7100", 96=>x"9f00", 97=>x"a200", 98=>x"9f00",
---- 99=>x"9900", 100=>x"9500", 101=>x"8b00", 102=>x"8000", 103=>x"7200", 104=>x"a000", 105=>x"a100",
---- 106=>x"a000", 107=>x"9900", 108=>x"9400", 109=>x"8b00", 110=>x"7b00", 111=>x"6c00", 112=>x"a000",
---- 113=>x"a200", 114=>x"a100", 115=>x"9c00", 116=>x"9400", 117=>x"8a00", 118=>x"7b00", 119=>x"6d00",
---- 120=>x"a000", 121=>x"a400", 122=>x"a300", 123=>x"a000", 124=>x"9400", 125=>x"8900", 126=>x"7e00",
---- 127=>x"6e00", 128=>x"a000", 129=>x"a100", 130=>x"a100", 131=>x"9d00", 132=>x"9600", 133=>x"8c00",
---- 134=>x"8000", 135=>x"6f00", 136=>x"a000", 137=>x"a300", 138=>x"a200", 139=>x"9b00", 140=>x"9300",
---- 141=>x"8800", 142=>x"7c00", 143=>x"6c00", 144=>x"9f00", 145=>x"a100", 146=>x"a100", 147=>x"9c00",
---- 148=>x"9200", 149=>x"8700", 150=>x"7f00", 151=>x"6d00", 152=>x"5d00", 153=>x"a100", 154=>x"a000",
---- 155=>x"9a00", 156=>x"9100", 157=>x"8900", 158=>x"7f00", 159=>x"6d00", 160=>x"a100", 161=>x"a100",
---- 162=>x"9f00", 163=>x"9b00", 164=>x"9400", 165=>x"8700", 166=>x"7b00", 167=>x"6900", 168=>x"5f00",
---- 169=>x"a100", 170=>x"a000", 171=>x"9a00", 172=>x"9100", 173=>x"8900", 174=>x"7b00", 175=>x"6900",
---- 176=>x"a000", 177=>x"a200", 178=>x"a000", 179=>x"9900", 180=>x"9400", 181=>x"8900", 182=>x"7c00",
---- 183=>x"6a00", 184=>x"a200", 185=>x"a400", 186=>x"a100", 187=>x"9a00", 188=>x"9500", 189=>x"8b00",
---- 190=>x"7d00", 191=>x"6b00", 192=>x"a400", 193=>x"5d00", 194=>x"a000", 195=>x"9c00", 196=>x"9500",
---- 197=>x"8a00", 198=>x"8200", 199=>x"7000", 200=>x"a400", 201=>x"a400", 202=>x"a100", 203=>x"9c00",
---- 204=>x"9500", 205=>x"8900", 206=>x"8100", 207=>x"6c00", 208=>x"a500", 209=>x"a400", 210=>x"a200",
---- 211=>x"9b00", 212=>x"9300", 213=>x"8a00", 214=>x"7f00", 215=>x"6c00", 216=>x"a600", 217=>x"a400",
---- 218=>x"a200", 219=>x"9d00", 220=>x"9100", 221=>x"8d00", 222=>x"7e00", 223=>x"6c00", 224=>x"a600",
---- 225=>x"a500", 226=>x"a400", 227=>x"9f00", 228=>x"9500", 229=>x"8b00", 230=>x"8000", 231=>x"6c00",
---- 232=>x"a500", 233=>x"a400", 234=>x"a000", 235=>x"9c00", 236=>x"6900", 237=>x"8b00", 238=>x"7e00",
---- 239=>x"6800", 240=>x"a400", 241=>x"a500", 242=>x"a100", 243=>x"9f00", 244=>x"9600", 245=>x"8d00",
---- 246=>x"8000", 247=>x"6b00", 248=>x"a600", 249=>x"a500", 250=>x"a300", 251=>x"9d00", 252=>x"9600",
---- 253=>x"8b00", 254=>x"8000", 255=>x"6e00", 256=>x"a600", 257=>x"a600", 258=>x"a400", 259=>x"9d00",
---- 260=>x"9600", 261=>x"8b00", 262=>x"7d00", 263=>x"6a00", 264=>x"a300", 265=>x"a300", 266=>x"a200",
---- 267=>x"9b00", 268=>x"9400", 269=>x"8b00", 270=>x"7e00", 271=>x"6d00", 272=>x"a300", 273=>x"a300",
---- 274=>x"a100", 275=>x"9a00", 276=>x"9100", 277=>x"8800", 278=>x"7f00", 279=>x"6b00", 280=>x"a600",
---- 281=>x"a500", 282=>x"a000", 283=>x"9b00", 284=>x"8f00", 285=>x"8800", 286=>x"7d00", 287=>x"6b00",
---- 288=>x"a200", 289=>x"a200", 290=>x"a000", 291=>x"9a00", 292=>x"9100", 293=>x"8900", 294=>x"7c00",
---- 295=>x"6a00", 296=>x"a500", 297=>x"a300", 298=>x"a000", 299=>x"9900", 300=>x"9200", 301=>x"8700",
---- 302=>x"8200", 303=>x"6c00", 304=>x"a400", 305=>x"a300", 306=>x"a000", 307=>x"9900", 308=>x"9300",
---- 309=>x"8900", 310=>x"7a00", 311=>x"6700", 312=>x"a300", 313=>x"a100", 314=>x"a000", 315=>x"9c00",
---- 316=>x"9400", 317=>x"8a00", 318=>x"7b00", 319=>x"6b00", 320=>x"a400", 321=>x"a300", 322=>x"5f00",
---- 323=>x"9a00", 324=>x"9300", 325=>x"8900", 326=>x"7900", 327=>x"6800", 328=>x"a600", 329=>x"a300",
---- 330=>x"9f00", 331=>x"9a00", 332=>x"9100", 333=>x"8600", 334=>x"7900", 335=>x"6700", 336=>x"a600",
---- 337=>x"a200", 338=>x"9d00", 339=>x"9800", 340=>x"8f00", 341=>x"8600", 342=>x"7500", 343=>x"6b00",
---- 344=>x"a600", 345=>x"a500", 346=>x"9e00", 347=>x"9800", 348=>x"9000", 349=>x"8600", 350=>x"7900",
---- 351=>x"6a00", 352=>x"a800", 353=>x"a500", 354=>x"9e00", 355=>x"9800", 356=>x"9000", 357=>x"8300",
---- 358=>x"7c00", 359=>x"6b00", 360=>x"a700", 361=>x"a400", 362=>x"9f00", 363=>x"9800", 364=>x"9000",
---- 365=>x"8400", 366=>x"7700", 367=>x"6a00", 368=>x"a400", 369=>x"a300", 370=>x"a000", 371=>x"9a00",
---- 372=>x"9000", 373=>x"8500", 374=>x"7900", 375=>x"6800", 376=>x"a600", 377=>x"a200", 378=>x"9f00",
---- 379=>x"9b00", 380=>x"9100", 381=>x"8400", 382=>x"7600", 383=>x"6700", 384=>x"a300", 385=>x"a400",
---- 386=>x"9e00", 387=>x"9a00", 388=>x"9200", 389=>x"8800", 390=>x"7800", 391=>x"6c00", 392=>x"a200",
---- 393=>x"a200", 394=>x"a000", 395=>x"9900", 396=>x"8e00", 397=>x"8500", 398=>x"7a00", 399=>x"6800",
---- 400=>x"a600", 401=>x"a300", 402=>x"a100", 403=>x"9800", 404=>x"9000", 405=>x"8600", 406=>x"7800",
---- 407=>x"6a00", 408=>x"a600", 409=>x"a300", 410=>x"a000", 411=>x"9a00", 412=>x"9100", 413=>x"8500",
---- 414=>x"7a00", 415=>x"6b00", 416=>x"a400", 417=>x"a300", 418=>x"9f00", 419=>x"6500", 420=>x"9200",
---- 421=>x"8600", 422=>x"7a00", 423=>x"6800", 424=>x"a000", 425=>x"a200", 426=>x"9f00", 427=>x"9a00",
---- 428=>x"9200", 429=>x"8900", 430=>x"7900", 431=>x"6900", 432=>x"a300", 433=>x"a300", 434=>x"a100",
---- 435=>x"9c00", 436=>x"6f00", 437=>x"8800", 438=>x"7900", 439=>x"6a00", 440=>x"a200", 441=>x"a400",
---- 442=>x"a400", 443=>x"9b00", 444=>x"9300", 445=>x"8800", 446=>x"7b00", 447=>x"6a00", 448=>x"a300",
---- 449=>x"a500", 450=>x"a400", 451=>x"9d00", 452=>x"9200", 453=>x"8700", 454=>x"7800", 455=>x"6c00",
---- 456=>x"a300", 457=>x"a300", 458=>x"a400", 459=>x"9b00", 460=>x"9200", 461=>x"8900", 462=>x"7d00",
---- 463=>x"7000", 464=>x"a300", 465=>x"a200", 466=>x"a100", 467=>x"9900", 468=>x"9300", 469=>x"8600",
---- 470=>x"7b00", 471=>x"6c00", 472=>x"a200", 473=>x"a400", 474=>x"a100", 475=>x"9a00", 476=>x"9100",
---- 477=>x"8800", 478=>x"7800", 479=>x"6800", 480=>x"a400", 481=>x"a500", 482=>x"a200", 483=>x"9a00",
---- 484=>x"9100", 485=>x"8600", 486=>x"7a00", 487=>x"6a00", 488=>x"a300", 489=>x"a200", 490=>x"a000",
---- 491=>x"9c00", 492=>x"9300", 493=>x"8600", 494=>x"7b00", 495=>x"6500", 496=>x"a400", 497=>x"a400",
---- 498=>x"a100", 499=>x"9a00", 500=>x"9300", 501=>x"8600", 502=>x"7700", 503=>x"6600", 504=>x"a600",
---- 505=>x"a700", 506=>x"a000", 507=>x"9900", 508=>x"9300", 509=>x"8600", 510=>x"7a00", 511=>x"6900",
---- 512=>x"a700", 513=>x"a700", 514=>x"a100", 515=>x"9b00", 516=>x"9500", 517=>x"8a00", 518=>x"7700",
---- 519=>x"6800", 520=>x"a500", 521=>x"a500", 522=>x"a400", 523=>x"9e00", 524=>x"9600", 525=>x"8b00",
---- 526=>x"7a00", 527=>x"6b00", 528=>x"a700", 529=>x"a700", 530=>x"a700", 531=>x"9e00", 532=>x"9800",
---- 533=>x"8d00", 534=>x"7a00", 535=>x"6a00", 536=>x"a800", 537=>x"aa00", 538=>x"a600", 539=>x"9e00",
---- 540=>x"9600", 541=>x"8c00", 542=>x"7900", 543=>x"6900", 544=>x"a800", 545=>x"a800", 546=>x"a500",
---- 547=>x"a100", 548=>x"9800", 549=>x"8c00", 550=>x"7b00", 551=>x"6e00", 552=>x"a900", 553=>x"a900",
---- 554=>x"aa00", 555=>x"a000", 556=>x"9800", 557=>x"8b00", 558=>x"7b00", 559=>x"6f00", 560=>x"ab00",
---- 561=>x"ac00", 562=>x"aa00", 563=>x"a300", 564=>x"9900", 565=>x"8d00", 566=>x"7e00", 567=>x"6c00",
---- 568=>x"ab00", 569=>x"ad00", 570=>x"aa00", 571=>x"a300", 572=>x"6400", 573=>x"8e00", 574=>x"7e00",
---- 575=>x"6900", 576=>x"ae00", 577=>x"af00", 578=>x"ac00", 579=>x"a600", 580=>x"9b00", 581=>x"8e00",
---- 582=>x"7e00", 583=>x"6a00", 584=>x"ad00", 585=>x"ad00", 586=>x"ac00", 587=>x"a600", 588=>x"9a00",
---- 589=>x"9000", 590=>x"7d00", 591=>x"6e00", 592=>x"ad00", 593=>x"af00", 594=>x"aa00", 595=>x"a500",
---- 596=>x"9b00", 597=>x"8f00", 598=>x"7c00", 599=>x"6e00", 600=>x"ab00", 601=>x"ae00", 602=>x"ab00",
---- 603=>x"a500", 604=>x"9a00", 605=>x"8d00", 606=>x"7c00", 607=>x"6e00", 608=>x"ae00", 609=>x"b000",
---- 610=>x"ab00", 611=>x"a500", 612=>x"9800", 613=>x"8d00", 614=>x"7f00", 615=>x"7000", 616=>x"ac00",
---- 617=>x"ae00", 618=>x"aa00", 619=>x"a400", 620=>x"9a00", 621=>x"8e00", 622=>x"8100", 623=>x"6f00",
---- 624=>x"5300", 625=>x"ad00", 626=>x"ac00", 627=>x"a300", 628=>x"9a00", 629=>x"8f00", 630=>x"7e00",
---- 631=>x"6c00", 632=>x"aa00", 633=>x"ab00", 634=>x"a900", 635=>x"a400", 636=>x"9b00", 637=>x"8f00",
---- 638=>x"8100", 639=>x"6c00", 640=>x"aa00", 641=>x"ab00", 642=>x"a700", 643=>x"a300", 644=>x"9a00",
---- 645=>x"8f00", 646=>x"7f00", 647=>x"6c00", 648=>x"ac00", 649=>x"ac00", 650=>x"aa00", 651=>x"a400",
---- 652=>x"9b00", 653=>x"9300", 654=>x"8000", 655=>x"6c00", 656=>x"ad00", 657=>x"ab00", 658=>x"ab00",
---- 659=>x"a500", 660=>x"9a00", 661=>x"9100", 662=>x"8300", 663=>x"6c00", 664=>x"ad00", 665=>x"ab00",
---- 666=>x"aa00", 667=>x"a600", 668=>x"9a00", 669=>x"9200", 670=>x"8300", 671=>x"6d00", 672=>x"ad00",
---- 673=>x"ad00", 674=>x"a900", 675=>x"a400", 676=>x"9c00", 677=>x"9400", 678=>x"8400", 679=>x"7200",
---- 680=>x"ab00", 681=>x"ab00", 682=>x"a800", 683=>x"a300", 684=>x"9d00", 685=>x"9400", 686=>x"8600",
---- 687=>x"6d00", 688=>x"aa00", 689=>x"ab00", 690=>x"aa00", 691=>x"a700", 692=>x"9d00", 693=>x"9100",
---- 694=>x"8300", 695=>x"6c00", 696=>x"ae00", 697=>x"ad00", 698=>x"ab00", 699=>x"a800", 700=>x"9f00",
---- 701=>x"9400", 702=>x"8500", 703=>x"6e00", 704=>x"ad00", 705=>x"ac00", 706=>x"ab00", 707=>x"a600",
---- 708=>x"9f00", 709=>x"9400", 710=>x"8300", 711=>x"6f00", 712=>x"ac00", 713=>x"ad00", 714=>x"ac00",
---- 715=>x"a500", 716=>x"9f00", 717=>x"9300", 718=>x"8300", 719=>x"6e00", 720=>x"ae00", 721=>x"ae00",
---- 722=>x"ac00", 723=>x"a700", 724=>x"9e00", 725=>x"9200", 726=>x"8500", 727=>x"7000", 728=>x"ac00",
---- 729=>x"ad00", 730=>x"ad00", 731=>x"a600", 732=>x"9e00", 733=>x"9500", 734=>x"8500", 735=>x"7200",
---- 736=>x"ae00", 737=>x"ad00", 738=>x"ad00", 739=>x"a600", 740=>x"9f00", 741=>x"9400", 742=>x"8700",
---- 743=>x"6e00", 744=>x"ad00", 745=>x"ac00", 746=>x"aa00", 747=>x"a700", 748=>x"a100", 749=>x"9300",
---- 750=>x"8400", 751=>x"6f00", 752=>x"ac00", 753=>x"ac00", 754=>x"ac00", 755=>x"a600", 756=>x"a000",
---- 757=>x"9400", 758=>x"8600", 759=>x"6f00", 760=>x"ac00", 761=>x"ac00", 762=>x"ab00", 763=>x"a700",
---- 764=>x"a000", 765=>x"9400", 766=>x"8500", 767=>x"6f00", 768=>x"aa00", 769=>x"aa00", 770=>x"aa00",
---- 771=>x"a600", 772=>x"9e00", 773=>x"9600", 774=>x"8600", 775=>x"7200", 776=>x"ab00", 777=>x"ab00",
---- 778=>x"ab00", 779=>x"a700", 780=>x"9f00", 781=>x"9400", 782=>x"8700", 783=>x"7100", 784=>x"ab00",
---- 785=>x"ac00", 786=>x"ab00", 787=>x"a800", 788=>x"9e00", 789=>x"9200", 790=>x"8700", 791=>x"7100",
---- 792=>x"ac00", 793=>x"ab00", 794=>x"aa00", 795=>x"a600", 796=>x"9d00", 797=>x"9400", 798=>x"8600",
---- 799=>x"8b00", 800=>x"aa00", 801=>x"ab00", 802=>x"ad00", 803=>x"a800", 804=>x"a000", 805=>x"9500",
---- 806=>x"8b00", 807=>x"7600", 808=>x"ac00", 809=>x"ab00", 810=>x"ae00", 811=>x"a500", 812=>x"9f00",
---- 813=>x"6b00", 814=>x"8800", 815=>x"7600", 816=>x"ae00", 817=>x"ad00", 818=>x"ac00", 819=>x"a500",
---- 820=>x"9f00", 821=>x"9600", 822=>x"8800", 823=>x"7400", 824=>x"ae00", 825=>x"ad00", 826=>x"ab00",
---- 827=>x"a800", 828=>x"9f00", 829=>x"6900", 830=>x"8800", 831=>x"7500", 832=>x"af00", 833=>x"b100",
---- 834=>x"ae00", 835=>x"a900", 836=>x"9f00", 837=>x"6b00", 838=>x"8700", 839=>x"7400", 840=>x"ae00",
---- 841=>x"ae00", 842=>x"ae00", 843=>x"aa00", 844=>x"9e00", 845=>x"9600", 846=>x"8b00", 847=>x"7400",
---- 848=>x"af00", 849=>x"ae00", 850=>x"ac00", 851=>x"a800", 852=>x"a000", 853=>x"9600", 854=>x"8900",
---- 855=>x"7700", 856=>x"ae00", 857=>x"ae00", 858=>x"ad00", 859=>x"a900", 860=>x"a100", 861=>x"9500",
---- 862=>x"8900", 863=>x"7800", 864=>x"af00", 865=>x"ae00", 866=>x"af00", 867=>x"aa00", 868=>x"9f00",
---- 869=>x"9700", 870=>x"8a00", 871=>x"7800", 872=>x"ac00", 873=>x"ae00", 874=>x"ae00", 875=>x"a800",
---- 876=>x"9e00", 877=>x"9800", 878=>x"8900", 879=>x"7400", 880=>x"ad00", 881=>x"ac00", 882=>x"ac00",
---- 883=>x"a800", 884=>x"a100", 885=>x"9500", 886=>x"8a00", 887=>x"7500", 888=>x"ae00", 889=>x"ad00",
---- 890=>x"ad00", 891=>x"a700", 892=>x"a000", 893=>x"9a00", 894=>x"8b00", 895=>x"7600", 896=>x"ae00",
---- 897=>x"ad00", 898=>x"ad00", 899=>x"aa00", 900=>x"a100", 901=>x"6600", 902=>x"8c00", 903=>x"7a00",
---- 904=>x"b000", 905=>x"ad00", 906=>x"ad00", 907=>x"ad00", 908=>x"a100", 909=>x"9600", 910=>x"8a00",
---- 911=>x"7900", 912=>x"ae00", 913=>x"ae00", 914=>x"ad00", 915=>x"ab00", 916=>x"a200", 917=>x"9700",
---- 918=>x"8900", 919=>x"7700", 920=>x"ad00", 921=>x"b000", 922=>x"ae00", 923=>x"aa00", 924=>x"a000",
---- 925=>x"9600", 926=>x"8a00", 927=>x"7800", 928=>x"af00", 929=>x"5100", 930=>x"af00", 931=>x"ab00",
---- 932=>x"a100", 933=>x"9600", 934=>x"8b00", 935=>x"7600", 936=>x"b000", 937=>x"ad00", 938=>x"ad00",
---- 939=>x"aa00", 940=>x"a100", 941=>x"9400", 942=>x"8b00", 943=>x"7700", 944=>x"4e00", 945=>x"ae00",
---- 946=>x"ac00", 947=>x"a700", 948=>x"a100", 949=>x"9900", 950=>x"8e00", 951=>x"7700", 952=>x"b100",
---- 953=>x"b000", 954=>x"af00", 955=>x"ab00", 956=>x"a000", 957=>x"9800", 958=>x"8b00", 959=>x"7500",
---- 960=>x"b100", 961=>x"af00", 962=>x"ad00", 963=>x"ab00", 964=>x"a100", 965=>x"9500", 966=>x"8900",
---- 967=>x"7500", 968=>x"af00", 969=>x"b000", 970=>x"b100", 971=>x"ac00", 972=>x"a100", 973=>x"9700",
---- 974=>x"8b00", 975=>x"7600", 976=>x"b100", 977=>x"af00", 978=>x"ae00", 979=>x"aa00", 980=>x"a300",
---- 981=>x"9900", 982=>x"8b00", 983=>x"7700", 984=>x"b100", 985=>x"b000", 986=>x"ad00", 987=>x"ab00",
---- 988=>x"a200", 989=>x"9800", 990=>x"8a00", 991=>x"7700", 992=>x"b100", 993=>x"b100", 994=>x"b100",
---- 995=>x"ac00", 996=>x"a200", 997=>x"6500", 998=>x"8c00", 999=>x"7500", 1000=>x"b100", 1001=>x"b400",
---- 1002=>x"b000", 1003=>x"ab00", 1004=>x"a300", 1005=>x"9800", 1006=>x"8e00", 1007=>x"7a00", 1008=>x"b000",
---- 1009=>x"b200", 1010=>x"b200", 1011=>x"ac00", 1012=>x"a200", 1013=>x"9600", 1014=>x"8c00", 1015=>x"7a00",
---- 1016=>x"b000", 1017=>x"b100", 1018=>x"b300", 1019=>x"ae00", 1020=>x"a200", 1021=>x"9b00", 1022=>x"8e00",
---- 1023=>x"7a00", 1024=>x"b000", 1025=>x"af00", 1026=>x"af00", 1027=>x"aa00", 1028=>x"a400", 1029=>x"9c00",
---- 1030=>x"9200", 1031=>x"7c00", 1032=>x"b100", 1033=>x"b100", 1034=>x"b000", 1035=>x"ab00", 1036=>x"a300",
---- 1037=>x"9a00", 1038=>x"8d00", 1039=>x"7c00", 1040=>x"b300", 1041=>x"b000", 1042=>x"b000", 1043=>x"aa00",
---- 1044=>x"a000", 1045=>x"9700", 1046=>x"8e00", 1047=>x"7b00", 1048=>x"b100", 1049=>x"b000", 1050=>x"b000",
---- 1051=>x"aa00", 1052=>x"a000", 1053=>x"9a00", 1054=>x"8c00", 1055=>x"7a00", 1056=>x"b100", 1057=>x"b000",
---- 1058=>x"b100", 1059=>x"aa00", 1060=>x"a000", 1061=>x"9700", 1062=>x"8b00", 1063=>x"7800", 1064=>x"b200",
---- 1065=>x"b300", 1066=>x"b400", 1067=>x"b000", 1068=>x"a100", 1069=>x"9700", 1070=>x"8b00", 1071=>x"7900",
---- 1072=>x"b300", 1073=>x"b400", 1074=>x"b400", 1075=>x"ae00", 1076=>x"a400", 1077=>x"9700", 1078=>x"8a00",
---- 1079=>x"7b00", 1080=>x"4900", 1081=>x"b400", 1082=>x"b200", 1083=>x"ae00", 1084=>x"a500", 1085=>x"9600",
---- 1086=>x"8900", 1087=>x"7b00", 1088=>x"b500", 1089=>x"b300", 1090=>x"b300", 1091=>x"af00", 1092=>x"a500",
---- 1093=>x"9a00", 1094=>x"8900", 1095=>x"7800", 1096=>x"b500", 1097=>x"b400", 1098=>x"b400", 1099=>x"4f00",
---- 1100=>x"a400", 1101=>x"9b00", 1102=>x"8a00", 1103=>x"7e00", 1104=>x"b500", 1105=>x"b600", 1106=>x"b500",
---- 1107=>x"b100", 1108=>x"a500", 1109=>x"9d00", 1110=>x"8e00", 1111=>x"7e00", 1112=>x"b800", 1113=>x"b700",
---- 1114=>x"b700", 1115=>x"b100", 1116=>x"a900", 1117=>x"9f00", 1118=>x"8e00", 1119=>x"7e00", 1120=>x"b700",
---- 1121=>x"b700", 1122=>x"b900", 1123=>x"b000", 1124=>x"aa00", 1125=>x"9f00", 1126=>x"8f00", 1127=>x"7e00",
---- 1128=>x"b800", 1129=>x"b800", 1130=>x"b500", 1131=>x"b200", 1132=>x"aa00", 1133=>x"9e00", 1134=>x"9000",
---- 1135=>x"8000", 1136=>x"b500", 1137=>x"b700", 1138=>x"b700", 1139=>x"b400", 1140=>x"a700", 1141=>x"9d00",
---- 1142=>x"9000", 1143=>x"8200", 1144=>x"b700", 1145=>x"b600", 1146=>x"b700", 1147=>x"b300", 1148=>x"a800",
---- 1149=>x"9f00", 1150=>x"8f00", 1151=>x"7f00", 1152=>x"b700", 1153=>x"b600", 1154=>x"b600", 1155=>x"b200",
---- 1156=>x"a800", 1157=>x"9f00", 1158=>x"9000", 1159=>x"8000", 1160=>x"b600", 1161=>x"b600", 1162=>x"b500",
---- 1163=>x"b000", 1164=>x"a800", 1165=>x"9e00", 1166=>x"9000", 1167=>x"7e00", 1168=>x"b400", 1169=>x"b600",
---- 1170=>x"b600", 1171=>x"b200", 1172=>x"a600", 1173=>x"9e00", 1174=>x"8d00", 1175=>x"8000", 1176=>x"b300",
---- 1177=>x"b700", 1178=>x"b600", 1179=>x"b100", 1180=>x"a700", 1181=>x"9e00", 1182=>x"9100", 1183=>x"7f00",
---- 1184=>x"b600", 1185=>x"b600", 1186=>x"b400", 1187=>x"af00", 1188=>x"a800", 1189=>x"9b00", 1190=>x"9100",
---- 1191=>x"7e00", 1192=>x"b500", 1193=>x"b300", 1194=>x"b400", 1195=>x"b000", 1196=>x"a700", 1197=>x"9900",
---- 1198=>x"9200", 1199=>x"7f00", 1200=>x"4d00", 1201=>x"b100", 1202=>x"b100", 1203=>x"ae00", 1204=>x"a400",
---- 1205=>x"9d00", 1206=>x"9000", 1207=>x"8000", 1208=>x"af00", 1209=>x"b200", 1210=>x"b000", 1211=>x"ad00",
---- 1212=>x"a600", 1213=>x"9c00", 1214=>x"9000", 1215=>x"8100", 1216=>x"af00", 1217=>x"af00", 1218=>x"b200",
---- 1219=>x"ac00", 1220=>x"a400", 1221=>x"9900", 1222=>x"9100", 1223=>x"8100", 1224=>x"b000", 1225=>x"b300",
---- 1226=>x"b100", 1227=>x"ac00", 1228=>x"a300", 1229=>x"9a00", 1230=>x"9000", 1231=>x"7f00", 1232=>x"ad00",
---- 1233=>x"b000", 1234=>x"b000", 1235=>x"ab00", 1236=>x"a400", 1237=>x"9a00", 1238=>x"8f00", 1239=>x"7f00",
---- 1240=>x"ac00", 1241=>x"b000", 1242=>x"b100", 1243=>x"ac00", 1244=>x"a400", 1245=>x"9a00", 1246=>x"9000",
---- 1247=>x"8000", 1248=>x"ae00", 1249=>x"b000", 1250=>x"b200", 1251=>x"ae00", 1252=>x"a500", 1253=>x"9d00",
---- 1254=>x"9100", 1255=>x"7e00", 1256=>x"b000", 1257=>x"b200", 1258=>x"b400", 1259=>x"ad00", 1260=>x"a600",
---- 1261=>x"9d00", 1262=>x"9100", 1263=>x"7f00", 1264=>x"b000", 1265=>x"b100", 1266=>x"b500", 1267=>x"b000",
---- 1268=>x"a900", 1269=>x"9e00", 1270=>x"9000", 1271=>x"7f00", 1272=>x"4f00", 1273=>x"b200", 1274=>x"b400",
---- 1275=>x"af00", 1276=>x"a800", 1277=>x"9d00", 1278=>x"9200", 1279=>x"7f00", 1280=>x"b100", 1281=>x"b200",
---- 1282=>x"b300", 1283=>x"af00", 1284=>x"a900", 1285=>x"9e00", 1286=>x"8f00", 1287=>x"7f00", 1288=>x"af00",
---- 1289=>x"b100", 1290=>x"b300", 1291=>x"b100", 1292=>x"a800", 1293=>x"9b00", 1294=>x"9000", 1295=>x"8300",
---- 1296=>x"5000", 1297=>x"b100", 1298=>x"b400", 1299=>x"af00", 1300=>x"aa00", 1301=>x"9e00", 1302=>x"9000",
---- 1303=>x"8500", 1304=>x"b000", 1305=>x"b200", 1306=>x"b300", 1307=>x"b000", 1308=>x"aa00", 1309=>x"a000",
---- 1310=>x"9100", 1311=>x"8300", 1312=>x"ae00", 1313=>x"b100", 1314=>x"b400", 1315=>x"b300", 1316=>x"a900",
---- 1317=>x"9e00", 1318=>x"9200", 1319=>x"8400", 1320=>x"af00", 1321=>x"b000", 1322=>x"b400", 1323=>x"b300",
---- 1324=>x"ab00", 1325=>x"9e00", 1326=>x"9200", 1327=>x"8400", 1328=>x"ad00", 1329=>x"b100", 1330=>x"b100",
---- 1331=>x"b200", 1332=>x"ab00", 1333=>x"a000", 1334=>x"9400", 1335=>x"8200", 1336=>x"b000", 1337=>x"b300",
---- 1338=>x"b600", 1339=>x"b200", 1340=>x"ab00", 1341=>x"a100", 1342=>x"9400", 1343=>x"8700", 1344=>x"af00",
---- 1345=>x"b400", 1346=>x"b200", 1347=>x"b000", 1348=>x"aa00", 1349=>x"a000", 1350=>x"9400", 1351=>x"8400",
---- 1352=>x"af00", 1353=>x"b300", 1354=>x"b600", 1355=>x"b100", 1356=>x"ab00", 1357=>x"a100", 1358=>x"9400",
---- 1359=>x"8500", 1360=>x"ae00", 1361=>x"b000", 1362=>x"b400", 1363=>x"b300", 1364=>x"aa00", 1365=>x"a200",
---- 1366=>x"9400", 1367=>x"8400", 1368=>x"b000", 1369=>x"b100", 1370=>x"b400", 1371=>x"b200", 1372=>x"ad00",
---- 1373=>x"5c00", 1374=>x"9700", 1375=>x"8600", 1376=>x"b100", 1377=>x"b300", 1378=>x"b600", 1379=>x"b200",
---- 1380=>x"ae00", 1381=>x"a400", 1382=>x"9400", 1383=>x"8600", 1384=>x"b000", 1385=>x"b400", 1386=>x"b500",
---- 1387=>x"b300", 1388=>x"ae00", 1389=>x"a400", 1390=>x"9700", 1391=>x"8400", 1392=>x"b100", 1393=>x"b500",
---- 1394=>x"b500", 1395=>x"b300", 1396=>x"ad00", 1397=>x"a100", 1398=>x"9500", 1399=>x"8300", 1400=>x"b300",
---- 1401=>x"b300", 1402=>x"b200", 1403=>x"b300", 1404=>x"ac00", 1405=>x"a300", 1406=>x"9400", 1407=>x"8000",
---- 1408=>x"b200", 1409=>x"b300", 1410=>x"b500", 1411=>x"4c00", 1412=>x"aa00", 1413=>x"a100", 1414=>x"9200",
---- 1415=>x"8100", 1416=>x"b300", 1417=>x"b600", 1418=>x"b600", 1419=>x"b300", 1420=>x"a800", 1421=>x"9f00",
---- 1422=>x"9400", 1423=>x"8200", 1424=>x"b500", 1425=>x"b600", 1426=>x"b600", 1427=>x"b200", 1428=>x"a900",
---- 1429=>x"5e00", 1430=>x"9500", 1431=>x"7d00", 1432=>x"b200", 1433=>x"b400", 1434=>x"b400", 1435=>x"b000",
---- 1436=>x"a900", 1437=>x"a800", 1438=>x"9b00", 1439=>x"8300", 1440=>x"b600", 1441=>x"b600", 1442=>x"b700",
---- 1443=>x"b300", 1444=>x"aa00", 1445=>x"a800", 1446=>x"ae00", 1447=>x"9900", 1448=>x"b400", 1449=>x"b400",
---- 1450=>x"b600", 1451=>x"4b00", 1452=>x"ac00", 1453=>x"a100", 1454=>x"9900", 1455=>x"8400", 1456=>x"b300",
---- 1457=>x"b500", 1458=>x"b500", 1459=>x"b300", 1460=>x"ac00", 1461=>x"9f00", 1462=>x"9300", 1463=>x"8000",
---- 1464=>x"b300", 1465=>x"b600", 1466=>x"b600", 1467=>x"b200", 1468=>x"aa00", 1469=>x"a000", 1470=>x"9400",
---- 1471=>x"8200", 1472=>x"b200", 1473=>x"b400", 1474=>x"b500", 1475=>x"b200", 1476=>x"ab00", 1477=>x"a200",
---- 1478=>x"6900", 1479=>x"8600", 1480=>x"b100", 1481=>x"b300", 1482=>x"b500", 1483=>x"b200", 1484=>x"aa00",
---- 1485=>x"a300", 1486=>x"9800", 1487=>x"8500", 1488=>x"b000", 1489=>x"b300", 1490=>x"b500", 1491=>x"b000",
---- 1492=>x"a900", 1493=>x"a000", 1494=>x"9500", 1495=>x"8400", 1496=>x"b000", 1497=>x"b200", 1498=>x"b300",
---- 1499=>x"b200", 1500=>x"aa00", 1501=>x"a200", 1502=>x"9600", 1503=>x"7b00", 1504=>x"4e00", 1505=>x"b100",
---- 1506=>x"b100", 1507=>x"b200", 1508=>x"a900", 1509=>x"a100", 1510=>x"9400", 1511=>x"8100", 1512=>x"b100",
---- 1513=>x"b000", 1514=>x"b300", 1515=>x"b200", 1516=>x"aa00", 1517=>x"a200", 1518=>x"9400", 1519=>x"8500",
---- 1520=>x"b300", 1521=>x"b100", 1522=>x"b300", 1523=>x"b200", 1524=>x"aa00", 1525=>x"a300", 1526=>x"9800",
---- 1527=>x"8300", 1528=>x"b000", 1529=>x"b200", 1530=>x"b300", 1531=>x"b200", 1532=>x"ae00", 1533=>x"a300",
---- 1534=>x"9700", 1535=>x"8600", 1536=>x"b100", 1537=>x"b200", 1538=>x"4d00", 1539=>x"b000", 1540=>x"ab00",
---- 1541=>x"a300", 1542=>x"9400", 1543=>x"8400", 1544=>x"b000", 1545=>x"b000", 1546=>x"b400", 1547=>x"b200",
---- 1548=>x"a800", 1549=>x"a000", 1550=>x"9200", 1551=>x"7f00", 1552=>x"af00", 1553=>x"af00", 1554=>x"b100",
---- 1555=>x"af00", 1556=>x"a800", 1557=>x"9e00", 1558=>x"9100", 1559=>x"7a00", 1560=>x"ad00", 1561=>x"ac00",
---- 1562=>x"ae00", 1563=>x"b000", 1564=>x"a800", 1565=>x"9d00", 1566=>x"8d00", 1567=>x"7800", 1568=>x"ad00",
---- 1569=>x"ae00", 1570=>x"af00", 1571=>x"af00", 1572=>x"a800", 1573=>x"9900", 1574=>x"8c00", 1575=>x"7b00",
---- 1576=>x"ab00", 1577=>x"ad00", 1578=>x"af00", 1579=>x"ad00", 1580=>x"a600", 1581=>x"9b00", 1582=>x"9000",
---- 1583=>x"a800", 1584=>x"ab00", 1585=>x"ac00", 1586=>x"ae00", 1587=>x"ad00", 1588=>x"a600", 1589=>x"a000",
---- 1590=>x"b600", 1591=>x"c300", 1592=>x"ab00", 1593=>x"ab00", 1594=>x"ac00", 1595=>x"b200", 1596=>x"b900",
---- 1597=>x"b600", 1598=>x"ac00", 1599=>x"8600", 1600=>x"ac00", 1601=>x"ab00", 1602=>x"b000", 1603=>x"bb00",
---- 1604=>x"bd00", 1605=>x"a800", 1606=>x"9500", 1607=>x"8100", 1608=>x"ac00", 1609=>x"a800", 1610=>x"b000",
---- 1611=>x"b100", 1612=>x"a900", 1613=>x"a200", 1614=>x"9700", 1615=>x"8500", 1616=>x"ab00", 1617=>x"ab00",
---- 1618=>x"ab00", 1619=>x"ac00", 1620=>x"a900", 1621=>x"a200", 1622=>x"9600", 1623=>x"7f00", 1624=>x"ab00",
---- 1625=>x"ae00", 1626=>x"ae00", 1627=>x"ae00", 1628=>x"a800", 1629=>x"9f00", 1630=>x"9300", 1631=>x"7d00",
---- 1632=>x"ac00", 1633=>x"ac00", 1634=>x"af00", 1635=>x"af00", 1636=>x"a800", 1637=>x"a000", 1638=>x"8f00",
---- 1639=>x"8800", 1640=>x"ad00", 1641=>x"ac00", 1642=>x"b100", 1643=>x"b000", 1644=>x"a800", 1645=>x"a100",
---- 1646=>x"8d00", 1647=>x"9800", 1648=>x"ad00", 1649=>x"af00", 1650=>x"b100", 1651=>x"ae00", 1652=>x"a700",
---- 1653=>x"9e00", 1654=>x"8f00", 1655=>x"a300", 1656=>x"af00", 1657=>x"ae00", 1658=>x"4d00", 1659=>x"b000",
---- 1660=>x"a900", 1661=>x"a100", 1662=>x"9100", 1663=>x"9400", 1664=>x"ae00", 1665=>x"b100", 1666=>x"b400",
---- 1667=>x"b100", 1668=>x"a900", 1669=>x"a200", 1670=>x"9200", 1671=>x"9400", 1672=>x"b000", 1673=>x"b300",
---- 1674=>x"b400", 1675=>x"b000", 1676=>x"aa00", 1677=>x"9e00", 1678=>x"9400", 1679=>x"9e00", 1680=>x"b100",
---- 1681=>x"b200", 1682=>x"b300", 1683=>x"b000", 1684=>x"a900", 1685=>x"a200", 1686=>x"9400", 1687=>x"9300",
---- 1688=>x"b200", 1689=>x"b100", 1690=>x"b300", 1691=>x"b100", 1692=>x"a900", 1693=>x"a200", 1694=>x"9800",
---- 1695=>x"8800", 1696=>x"af00", 1697=>x"b200", 1698=>x"b200", 1699=>x"b200", 1700=>x"ac00", 1701=>x"a400",
---- 1702=>x"9a00", 1703=>x"8a00", 1704=>x"af00", 1705=>x"b300", 1706=>x"b300", 1707=>x"b200", 1708=>x"ac00",
---- 1709=>x"a500", 1710=>x"9b00", 1711=>x"8a00", 1712=>x"b200", 1713=>x"b300", 1714=>x"b500", 1715=>x"b200",
---- 1716=>x"ad00", 1717=>x"a600", 1718=>x"9c00", 1719=>x"8d00", 1720=>x"b100", 1721=>x"b200", 1722=>x"b600",
---- 1723=>x"b500", 1724=>x"af00", 1725=>x"a700", 1726=>x"9c00", 1727=>x"8800", 1728=>x"b300", 1729=>x"b100",
---- 1730=>x"b500", 1731=>x"b600", 1732=>x"af00", 1733=>x"a600", 1734=>x"9c00", 1735=>x"8700", 1736=>x"b200",
---- 1737=>x"b400", 1738=>x"b600", 1739=>x"b300", 1740=>x"ac00", 1741=>x"a500", 1742=>x"9b00", 1743=>x"8900",
---- 1744=>x"b300", 1745=>x"4b00", 1746=>x"b500", 1747=>x"b400", 1748=>x"ad00", 1749=>x"a600", 1750=>x"9c00",
---- 1751=>x"8900", 1752=>x"b300", 1753=>x"b300", 1754=>x"b400", 1755=>x"b400", 1756=>x"b000", 1757=>x"a700",
---- 1758=>x"9e00", 1759=>x"8c00", 1760=>x"b100", 1761=>x"b200", 1762=>x"b100", 1763=>x"b200", 1764=>x"ac00",
---- 1765=>x"a300", 1766=>x"9c00", 1767=>x"9200", 1768=>x"ac00", 1769=>x"a900", 1770=>x"a900", 1771=>x"ad00",
---- 1772=>x"a800", 1773=>x"a000", 1774=>x"9900", 1775=>x"8f00", 1776=>x"ad00", 1777=>x"ab00", 1778=>x"af00",
---- 1779=>x"b100", 1780=>x"aa00", 1781=>x"a300", 1782=>x"9900", 1783=>x"8b00", 1784=>x"b200", 1785=>x"b100",
---- 1786=>x"b300", 1787=>x"b200", 1788=>x"ac00", 1789=>x"a600", 1790=>x"9900", 1791=>x"9200", 1792=>x"b200",
---- 1793=>x"b200", 1794=>x"b500", 1795=>x"b300", 1796=>x"ae00", 1797=>x"a600", 1798=>x"9c00", 1799=>x"8d00",
---- 1800=>x"b200", 1801=>x"b200", 1802=>x"b300", 1803=>x"b300", 1804=>x"b000", 1805=>x"a600", 1806=>x"9800",
---- 1807=>x"8f00", 1808=>x"b200", 1809=>x"b100", 1810=>x"b200", 1811=>x"b300", 1812=>x"ae00", 1813=>x"a800",
---- 1814=>x"9500", 1815=>x"9800", 1816=>x"b000", 1817=>x"b100", 1818=>x"b100", 1819=>x"b200", 1820=>x"aa00",
---- 1821=>x"a500", 1822=>x"9800", 1823=>x"9000", 1824=>x"b000", 1825=>x"b100", 1826=>x"b200", 1827=>x"b200",
---- 1828=>x"ad00", 1829=>x"a400", 1830=>x"9800", 1831=>x"8c00", 1832=>x"b100", 1833=>x"b100", 1834=>x"b200",
---- 1835=>x"b300", 1836=>x"ad00", 1837=>x"a700", 1838=>x"9c00", 1839=>x"8700", 1840=>x"b000", 1841=>x"b000",
---- 1842=>x"b100", 1843=>x"b100", 1844=>x"ad00", 1845=>x"a700", 1846=>x"9d00", 1847=>x"8500", 1848=>x"b000",
---- 1849=>x"b200", 1850=>x"b300", 1851=>x"b300", 1852=>x"ae00", 1853=>x"5a00", 1854=>x"9e00", 1855=>x"8a00",
---- 1856=>x"b000", 1857=>x"b200", 1858=>x"b300", 1859=>x"b500", 1860=>x"af00", 1861=>x"a900", 1862=>x"9e00",
---- 1863=>x"8e00", 1864=>x"b200", 1865=>x"b000", 1866=>x"b100", 1867=>x"b200", 1868=>x"af00", 1869=>x"a800",
---- 1870=>x"9d00", 1871=>x"6d00", 1872=>x"b100", 1873=>x"af00", 1874=>x"b100", 1875=>x"b500", 1876=>x"b100",
---- 1877=>x"a600", 1878=>x"9e00", 1879=>x"9500", 1880=>x"b000", 1881=>x"b000", 1882=>x"b200", 1883=>x"b500",
---- 1884=>x"b200", 1885=>x"ab00", 1886=>x"a100", 1887=>x"8e00", 1888=>x"af00", 1889=>x"ae00", 1890=>x"b300",
---- 1891=>x"b600", 1892=>x"b300", 1893=>x"ac00", 1894=>x"a400", 1895=>x"8500", 1896=>x"ac00", 1897=>x"ae00",
---- 1898=>x"b400", 1899=>x"b700", 1900=>x"b100", 1901=>x"aa00", 1902=>x"a500", 1903=>x"7e00", 1904=>x"ae00",
---- 1905=>x"ad00", 1906=>x"b300", 1907=>x"b700", 1908=>x"b100", 1909=>x"ab00", 1910=>x"a000", 1911=>x"7600",
---- 1912=>x"b100", 1913=>x"b000", 1914=>x"b500", 1915=>x"ba00", 1916=>x"b100", 1917=>x"ae00", 1918=>x"9d00",
---- 1919=>x"7700", 1920=>x"b100", 1921=>x"b000", 1922=>x"b500", 1923=>x"b900", 1924=>x"b300", 1925=>x"ac00",
---- 1926=>x"9d00", 1927=>x"7000", 1928=>x"b200", 1929=>x"b300", 1930=>x"b600", 1931=>x"b800", 1932=>x"b200",
---- 1933=>x"af00", 1934=>x"a100", 1935=>x"6400", 1936=>x"b200", 1937=>x"b500", 1938=>x"b700", 1939=>x"b800",
---- 1940=>x"b100", 1941=>x"ac00", 1942=>x"a400", 1943=>x"6100", 1944=>x"b100", 1945=>x"b300", 1946=>x"b600",
---- 1947=>x"b800", 1948=>x"b200", 1949=>x"ab00", 1950=>x"a400", 1951=>x"6900", 1952=>x"b200", 1953=>x"b300",
---- 1954=>x"b600", 1955=>x"b700", 1956=>x"b300", 1957=>x"ab00", 1958=>x"a700", 1959=>x"6c00", 1960=>x"b400",
---- 1961=>x"b400", 1962=>x"b600", 1963=>x"b700", 1964=>x"b100", 1965=>x"aa00", 1966=>x"a700", 1967=>x"7a00",
---- 1968=>x"b500", 1969=>x"b400", 1970=>x"4800", 1971=>x"b900", 1972=>x"4900", 1973=>x"ad00", 1974=>x"a800",
---- 1975=>x"8700", 1976=>x"b400", 1977=>x"b400", 1978=>x"b600", 1979=>x"b900", 1980=>x"b500", 1981=>x"a800",
---- 1982=>x"a600", 1983=>x"9000", 1984=>x"b400", 1985=>x"b500", 1986=>x"b500", 1987=>x"b800", 1988=>x"b300",
---- 1989=>x"a900", 1990=>x"5900", 1991=>x"8f00", 1992=>x"b500", 1993=>x"b500", 1994=>x"b900", 1995=>x"b900",
---- 1996=>x"b400", 1997=>x"ad00", 1998=>x"a300", 1999=>x"7200", 2000=>x"b500", 2001=>x"b600", 2002=>x"ba00",
---- 2003=>x"bb00", 2004=>x"b600", 2005=>x"ac00", 2006=>x"8100", 2007=>x"4900", 2008=>x"b600", 2009=>x"b400",
---- 2010=>x"b700", 2011=>x"b800", 2012=>x"b400", 2013=>x"aa00", 2014=>x"8700", 2015=>x"6500", 2016=>x"b300",
---- 2017=>x"b200", 2018=>x"b500", 2019=>x"b500", 2020=>x"b200", 2021=>x"ae00", 2022=>x"9600", 2023=>x"8000",
---- 2024=>x"b300", 2025=>x"b300", 2026=>x"b400", 2027=>x"b700", 2028=>x"b300", 2029=>x"ac00", 2030=>x"8800",
---- 2031=>x"7500", 2032=>x"b400", 2033=>x"b400", 2034=>x"b400", 2035=>x"b700", 2036=>x"b400", 2037=>x"ad00",
---- 2038=>x"7700", 2039=>x"5a00", 2040=>x"b400", 2041=>x"b400", 2042=>x"b500", 2043=>x"b600", 2044=>x"b200",
---- 2045=>x"b200", 2046=>x"7800", 2047=>x"5500"),
---- 4  => (0=>x"6300", 1=>x"5d00", 2=>x"5b00", 3=>x"6400", 4=>x"6400", 5=>x"6700", 6=>x"6900", 7=>x"6900",
---- 8=>x"6300", 9=>x"5e00", 10=>x"5b00", 11=>x"6500", 12=>x"6400", 13=>x"6700", 14=>x"6900",
---- 15=>x"6900", 16=>x"6400", 17=>x"5e00", 18=>x"5c00", 19=>x"6300", 20=>x"9c00", 21=>x"6600",
---- 22=>x"6900", 23=>x"6900", 24=>x"6300", 25=>x"5b00", 26=>x"5a00", 27=>x"5e00", 28=>x"6100",
---- 29=>x"6000", 30=>x"6900", 31=>x"6c00", 32=>x"6300", 33=>x"5a00", 34=>x"5800", 35=>x"5a00",
---- 36=>x"5f00", 37=>x"6400", 38=>x"6600", 39=>x"6800", 40=>x"6000", 41=>x"5b00", 42=>x"5900",
---- 43=>x"5b00", 44=>x"6200", 45=>x"6100", 46=>x"6300", 47=>x"6700", 48=>x"6300", 49=>x"5900",
---- 50=>x"5900", 51=>x"5b00", 52=>x"5d00", 53=>x"6000", 54=>x"6300", 55=>x"6900", 56=>x"6400",
---- 57=>x"5a00", 58=>x"5c00", 59=>x"5b00", 60=>x"5d00", 61=>x"6500", 62=>x"6500", 63=>x"6600",
---- 64=>x"6100", 65=>x"5900", 66=>x"5700", 67=>x"5b00", 68=>x"5c00", 69=>x"6500", 70=>x"9700",
---- 71=>x"6200", 72=>x"6100", 73=>x"5b00", 74=>x"5700", 75=>x"5d00", 76=>x"5f00", 77=>x"6400",
---- 78=>x"6600", 79=>x"6200", 80=>x"6600", 81=>x"a300", 82=>x"5700", 83=>x"5d00", 84=>x"5e00",
---- 85=>x"6100", 86=>x"6700", 87=>x"6700", 88=>x"6100", 89=>x"5a00", 90=>x"5b00", 91=>x"5f00",
---- 92=>x"6100", 93=>x"6200", 94=>x"6400", 95=>x"6600", 96=>x"6300", 97=>x"5800", 98=>x"5600",
---- 99=>x"5d00", 100=>x"6000", 101=>x"6000", 102=>x"6300", 103=>x"6800", 104=>x"5c00", 105=>x"5800",
---- 106=>x"5200", 107=>x"5600", 108=>x"5d00", 109=>x"6000", 110=>x"6500", 111=>x"6700", 112=>x"5f00",
---- 113=>x"5700", 114=>x"5500", 115=>x"5700", 116=>x"5f00", 117=>x"6200", 118=>x"6400", 119=>x"6700",
---- 120=>x"6100", 121=>x"5a00", 122=>x"5600", 123=>x"5a00", 124=>x"6100", 125=>x"6200", 126=>x"6200",
---- 127=>x"6800", 128=>x"6100", 129=>x"5a00", 130=>x"5700", 131=>x"5e00", 132=>x"5f00", 133=>x"6000",
---- 134=>x"6400", 135=>x"6400", 136=>x"5f00", 137=>x"5800", 138=>x"5a00", 139=>x"5d00", 140=>x"5f00",
---- 141=>x"6400", 142=>x"6200", 143=>x"6700", 144=>x"6000", 145=>x"5600", 146=>x"5600", 147=>x"5a00",
---- 148=>x"6100", 149=>x"6100", 150=>x"6500", 151=>x"6600", 152=>x"5b00", 153=>x"5300", 154=>x"5300",
---- 155=>x"5700", 156=>x"5f00", 157=>x"5f00", 158=>x"6400", 159=>x"6500", 160=>x"5d00", 161=>x"5400",
---- 162=>x"5100", 163=>x"5b00", 164=>x"5e00", 165=>x"6000", 166=>x"6800", 167=>x"6800", 168=>x"5d00",
---- 169=>x"5400", 170=>x"5300", 171=>x"5900", 172=>x"5c00", 173=>x"6200", 174=>x"6700", 175=>x"6700",
---- 176=>x"5d00", 177=>x"5300", 178=>x"5300", 179=>x"5b00", 180=>x"5e00", 181=>x"6200", 182=>x"6400",
---- 183=>x"6500", 184=>x"5e00", 185=>x"5400", 186=>x"5100", 187=>x"5b00", 188=>x"5d00", 189=>x"5f00",
---- 190=>x"6200", 191=>x"6600", 192=>x"6100", 193=>x"5800", 194=>x"5300", 195=>x"5900", 196=>x"5e00",
---- 197=>x"6000", 198=>x"6200", 199=>x"6500", 200=>x"5c00", 201=>x"5600", 202=>x"5500", 203=>x"5900",
---- 204=>x"5c00", 205=>x"6000", 206=>x"6100", 207=>x"6300", 208=>x"5e00", 209=>x"5200", 210=>x"ae00",
---- 211=>x"5700", 212=>x"5e00", 213=>x"5c00", 214=>x"6200", 215=>x"6500", 216=>x"5c00", 217=>x"5100",
---- 218=>x"5500", 219=>x"5800", 220=>x"5d00", 221=>x"5e00", 222=>x"6300", 223=>x"6200", 224=>x"5900",
---- 225=>x"4f00", 226=>x"5000", 227=>x"5600", 228=>x"5600", 229=>x"5b00", 230=>x"6000", 231=>x"6000",
---- 232=>x"5900", 233=>x"4c00", 234=>x"4e00", 235=>x"5300", 236=>x"5a00", 237=>x"5f00", 238=>x"9c00",
---- 239=>x"6000", 240=>x"a600", 241=>x"5100", 242=>x"4e00", 243=>x"5300", 244=>x"5f00", 245=>x"5b00",
---- 246=>x"5e00", 247=>x"6100", 248=>x"5900", 249=>x"5200", 250=>x"4d00", 251=>x"5000", 252=>x"5700",
---- 253=>x"5600", 254=>x"5a00", 255=>x"5c00", 256=>x"5a00", 257=>x"4c00", 258=>x"4c00", 259=>x"5100",
---- 260=>x"5300", 261=>x"5600", 262=>x"5b00", 263=>x"5e00", 264=>x"5700", 265=>x"4b00", 266=>x"4900",
---- 267=>x"5100", 268=>x"5200", 269=>x"5700", 270=>x"5b00", 271=>x"5d00", 272=>x"5900", 273=>x"4e00",
---- 274=>x"4700", 275=>x"5000", 276=>x"5200", 277=>x"5a00", 278=>x"5e00", 279=>x"5d00", 280=>x"5500",
---- 281=>x"4b00", 282=>x"4700", 283=>x"5000", 284=>x"5700", 285=>x"5800", 286=>x"5900", 287=>x"5d00",
---- 288=>x"5300", 289=>x"4b00", 290=>x"4800", 291=>x"5000", 292=>x"5600", 293=>x"5800", 294=>x"5b00",
---- 295=>x"5f00", 296=>x"5300", 297=>x"4b00", 298=>x"4800", 299=>x"5000", 300=>x"5600", 301=>x"5a00",
---- 302=>x"5e00", 303=>x"6000", 304=>x"5400", 305=>x"4900", 306=>x"4b00", 307=>x"5100", 308=>x"5400",
---- 309=>x"5800", 310=>x"5c00", 311=>x"6000", 312=>x"5700", 313=>x"4a00", 314=>x"4e00", 315=>x"5100",
---- 316=>x"5800", 317=>x"5600", 318=>x"5c00", 319=>x"6200", 320=>x"5600", 321=>x"4d00", 322=>x"4700",
---- 323=>x"5000", 324=>x"5500", 325=>x"5900", 326=>x"5f00", 327=>x"6100", 328=>x"5400", 329=>x"4d00",
---- 330=>x"4a00", 331=>x"5000", 332=>x"5800", 333=>x"5a00", 334=>x"5e00", 335=>x"5f00", 336=>x"5900",
---- 337=>x"4c00", 338=>x"4a00", 339=>x"5000", 340=>x"5600", 341=>x"5a00", 342=>x"6100", 343=>x"5f00",
---- 344=>x"5b00", 345=>x"5000", 346=>x"4f00", 347=>x"5300", 348=>x"5800", 349=>x"5a00", 350=>x"5c00",
---- 351=>x"5c00", 352=>x"5900", 353=>x"4f00", 354=>x"4a00", 355=>x"5000", 356=>x"5500", 357=>x"5b00",
---- 358=>x"5c00", 359=>x"5e00", 360=>x"5800", 361=>x"4b00", 362=>x"4900", 363=>x"5200", 364=>x"5800",
---- 365=>x"5b00", 366=>x"5d00", 367=>x"6200", 368=>x"5a00", 369=>x"4c00", 370=>x"4b00", 371=>x"5300",
---- 372=>x"5800", 373=>x"5a00", 374=>x"6000", 375=>x"6100", 376=>x"a500", 377=>x"4d00", 378=>x"4e00",
---- 379=>x"5200", 380=>x"5800", 381=>x"5f00", 382=>x"6200", 383=>x"6100", 384=>x"5c00", 385=>x"4900",
---- 386=>x"4e00", 387=>x"5300", 388=>x"5900", 389=>x"5b00", 390=>x"6200", 391=>x"5d00", 392=>x"5a00",
---- 393=>x"4d00", 394=>x"4c00", 395=>x"4d00", 396=>x"5600", 397=>x"5c00", 398=>x"6000", 399=>x"6100",
---- 400=>x"5900", 401=>x"4c00", 402=>x"4b00", 403=>x"4d00", 404=>x"5600", 405=>x"5900", 406=>x"5e00",
---- 407=>x"6100", 408=>x"5e00", 409=>x"4e00", 410=>x"b700", 411=>x"4f00", 412=>x"5600", 413=>x"5800",
---- 414=>x"5e00", 415=>x"5f00", 416=>x"5e00", 417=>x"4e00", 418=>x"4900", 419=>x"5000", 420=>x"5500",
---- 421=>x"5a00", 422=>x"5e00", 423=>x"5e00", 424=>x"5900", 425=>x"5000", 426=>x"4c00", 427=>x"4e00",
---- 428=>x"5500", 429=>x"5b00", 430=>x"5e00", 431=>x"5f00", 432=>x"5e00", 433=>x"4f00", 434=>x"4b00",
---- 435=>x"5100", 436=>x"5500", 437=>x"5a00", 438=>x"5c00", 439=>x"5b00", 440=>x"a400", 441=>x"4e00",
---- 442=>x"4a00", 443=>x"5200", 444=>x"5500", 445=>x"5400", 446=>x"5a00", 447=>x"5d00", 448=>x"5900",
---- 449=>x"4c00", 450=>x"4a00", 451=>x"5100", 452=>x"5600", 453=>x"5600", 454=>x"5c00", 455=>x"6000",
---- 456=>x"5c00", 457=>x"5000", 458=>x"4b00", 459=>x"5000", 460=>x"5400", 461=>x"5a00", 462=>x"5d00",
---- 463=>x"5f00", 464=>x"5c00", 465=>x"4900", 466=>x"4700", 467=>x"4f00", 468=>x"5000", 469=>x"5600",
---- 470=>x"5800", 471=>x"5800", 472=>x"5600", 473=>x"4600", 474=>x"4700", 475=>x"4f00", 476=>x"5300",
---- 477=>x"5500", 478=>x"5800", 479=>x"5800", 480=>x"5300", 481=>x"4800", 482=>x"4600", 483=>x"4b00",
---- 484=>x"4f00", 485=>x"5300", 486=>x"5900", 487=>x"5c00", 488=>x"5600", 489=>x"4700", 490=>x"4500",
---- 491=>x"4a00", 492=>x"4d00", 493=>x"5200", 494=>x"5b00", 495=>x"5f00", 496=>x"5500", 497=>x"4d00",
---- 498=>x"4900", 499=>x"4c00", 500=>x"4900", 501=>x"5300", 502=>x"5800", 503=>x"5f00", 504=>x"5300",
---- 505=>x"4a00", 506=>x"4b00", 507=>x"4d00", 508=>x"4f00", 509=>x"5500", 510=>x"5b00", 511=>x"5e00",
---- 512=>x"5700", 513=>x"4900", 514=>x"4b00", 515=>x"4d00", 516=>x"5000", 517=>x"5700", 518=>x"5b00",
---- 519=>x"5c00", 520=>x"5900", 521=>x"5000", 522=>x"4c00", 523=>x"5000", 524=>x"5200", 525=>x"5700",
---- 526=>x"5b00", 527=>x"a100", 528=>x"5900", 529=>x"4f00", 530=>x"4c00", 531=>x"5100", 532=>x"5400",
---- 533=>x"5c00", 534=>x"6000", 535=>x"5f00", 536=>x"5800", 537=>x"4d00", 538=>x"4e00", 539=>x"5300",
---- 540=>x"5500", 541=>x"5700", 542=>x"5d00", 543=>x"5f00", 544=>x"5b00", 545=>x"4b00", 546=>x"4d00",
---- 547=>x"5000", 548=>x"5600", 549=>x"5400", 550=>x"5d00", 551=>x"5f00", 552=>x"a700", 553=>x"4d00",
---- 554=>x"4e00", 555=>x"5100", 556=>x"5500", 557=>x"5a00", 558=>x"5d00", 559=>x"5f00", 560=>x"5900",
---- 561=>x"4c00", 562=>x"4c00", 563=>x"4f00", 564=>x"5600", 565=>x"5d00", 566=>x"5d00", 567=>x"5e00",
---- 568=>x"5800", 569=>x"4e00", 570=>x"4d00", 571=>x"5000", 572=>x"5900", 573=>x"5b00", 574=>x"5d00",
---- 575=>x"6000", 576=>x"5b00", 577=>x"4d00", 578=>x"4e00", 579=>x"5200", 580=>x"5c00", 581=>x"6200",
---- 582=>x"5a00", 583=>x"5d00", 584=>x"5b00", 585=>x"4d00", 586=>x"4b00", 587=>x"4d00", 588=>x"5400",
---- 589=>x"5800", 590=>x"a500", 591=>x"5d00", 592=>x"5900", 593=>x"4e00", 594=>x"4c00", 595=>x"4f00",
---- 596=>x"5400", 597=>x"5a00", 598=>x"5d00", 599=>x"5e00", 600=>x"5900", 601=>x"4b00", 602=>x"4900",
---- 603=>x"5000", 604=>x"5400", 605=>x"5900", 606=>x"5b00", 607=>x"6000", 608=>x"5a00", 609=>x"4c00",
---- 610=>x"4b00", 611=>x"5100", 612=>x"5500", 613=>x"5b00", 614=>x"5e00", 615=>x"6000", 616=>x"5a00",
---- 617=>x"4f00", 618=>x"4d00", 619=>x"5100", 620=>x"5800", 621=>x"a500", 622=>x"5f00", 623=>x"5e00",
---- 624=>x"5900", 625=>x"5100", 626=>x"4d00", 627=>x"5200", 628=>x"5a00", 629=>x"5d00", 630=>x"6000",
---- 631=>x"5f00", 632=>x"5900", 633=>x"5000", 634=>x"4c00", 635=>x"5000", 636=>x"5500", 637=>x"5e00",
---- 638=>x"6000", 639=>x"5f00", 640=>x"5b00", 641=>x"4f00", 642=>x"4f00", 643=>x"4f00", 644=>x"5500",
---- 645=>x"5c00", 646=>x"5e00", 647=>x"6100", 648=>x"5b00", 649=>x"4b00", 650=>x"4d00", 651=>x"5000",
---- 652=>x"5500", 653=>x"5c00", 654=>x"5e00", 655=>x"6100", 656=>x"5e00", 657=>x"5000", 658=>x"4d00",
---- 659=>x"5300", 660=>x"5700", 661=>x"5d00", 662=>x"5e00", 663=>x"6100", 664=>x"5d00", 665=>x"4f00",
---- 666=>x"4c00", 667=>x"5300", 668=>x"5900", 669=>x"5b00", 670=>x"5c00", 671=>x"6200", 672=>x"6200",
---- 673=>x"4c00", 674=>x"4b00", 675=>x"5000", 676=>x"5600", 677=>x"5900", 678=>x"5c00", 679=>x"5f00",
---- 680=>x"5a00", 681=>x"4d00", 682=>x"4b00", 683=>x"4d00", 684=>x"5300", 685=>x"5a00", 686=>x"5f00",
---- 687=>x"6000", 688=>x"5a00", 689=>x"4f00", 690=>x"4700", 691=>x"5000", 692=>x"5400", 693=>x"5800",
---- 694=>x"a300", 695=>x"6200", 696=>x"5a00", 697=>x"4f00", 698=>x"4600", 699=>x"4c00", 700=>x"5600",
---- 701=>x"5900", 702=>x"5b00", 703=>x"6100", 704=>x"5900", 705=>x"4900", 706=>x"4700", 707=>x"4e00",
---- 708=>x"5300", 709=>x"5600", 710=>x"5c00", 711=>x"5f00", 712=>x"5b00", 713=>x"4a00", 714=>x"4800",
---- 715=>x"4d00", 716=>x"5100", 717=>x"5600", 718=>x"5e00", 719=>x"5e00", 720=>x"5b00", 721=>x"4e00",
---- 722=>x"4700", 723=>x"4c00", 724=>x"5300", 725=>x"5500", 726=>x"6000", 727=>x"5e00", 728=>x"5800",
---- 729=>x"4b00", 730=>x"4700", 731=>x"4f00", 732=>x"5300", 733=>x"5600", 734=>x"5e00", 735=>x"5f00",
---- 736=>x"5700", 737=>x"4d00", 738=>x"4800", 739=>x"5100", 740=>x"5300", 741=>x"5900", 742=>x"5d00",
---- 743=>x"6100", 744=>x"5a00", 745=>x"4b00", 746=>x"4900", 747=>x"5100", 748=>x"5100", 749=>x"5a00",
---- 750=>x"5e00", 751=>x"6000", 752=>x"5900", 753=>x"4e00", 754=>x"4d00", 755=>x"4e00", 756=>x"5100",
---- 757=>x"5800", 758=>x"5e00", 759=>x"5d00", 760=>x"5c00", 761=>x"4f00", 762=>x"4700", 763=>x"4d00",
---- 764=>x"5400", 765=>x"5b00", 766=>x"5c00", 767=>x"6000", 768=>x"5d00", 769=>x"4d00", 770=>x"4900",
---- 771=>x"4e00", 772=>x"5300", 773=>x"5500", 774=>x"5c00", 775=>x"5e00", 776=>x"5c00", 777=>x"4d00",
---- 778=>x"4900", 779=>x"4c00", 780=>x"5200", 781=>x"ac00", 782=>x"5b00", 783=>x"5e00", 784=>x"5c00",
---- 785=>x"4e00", 786=>x"4700", 787=>x"5000", 788=>x"aa00", 789=>x"5800", 790=>x"5d00", 791=>x"5e00",
---- 792=>x"a100", 793=>x"4e00", 794=>x"4800", 795=>x"4e00", 796=>x"a900", 797=>x"a600", 798=>x"5d00",
---- 799=>x"5e00", 800=>x"5c00", 801=>x"4a00", 802=>x"4500", 803=>x"4b00", 804=>x"5300", 805=>x"5900",
---- 806=>x"5b00", 807=>x"5b00", 808=>x"5b00", 809=>x"4b00", 810=>x"4400", 811=>x"4c00", 812=>x"5300",
---- 813=>x"5700", 814=>x"5b00", 815=>x"5b00", 816=>x"5900", 817=>x"4d00", 818=>x"4900", 819=>x"4d00",
---- 820=>x"5400", 821=>x"5400", 822=>x"5a00", 823=>x"5d00", 824=>x"5a00", 825=>x"4900", 826=>x"4800",
---- 827=>x"4d00", 828=>x"5200", 829=>x"5300", 830=>x"5800", 831=>x"5d00", 832=>x"5b00", 833=>x"4c00",
---- 834=>x"4600", 835=>x"4b00", 836=>x"5000", 837=>x"5500", 838=>x"5700", 839=>x"5b00", 840=>x"5900",
---- 841=>x"4b00", 842=>x"4400", 843=>x"4900", 844=>x"5000", 845=>x"5400", 846=>x"5900", 847=>x"5a00",
---- 848=>x"6000", 849=>x"4a00", 850=>x"4300", 851=>x"4a00", 852=>x"5100", 853=>x"5200", 854=>x"5800",
---- 855=>x"5900", 856=>x"5d00", 857=>x"4900", 858=>x"4300", 859=>x"4e00", 860=>x"4f00", 861=>x"5200",
---- 862=>x"5a00", 863=>x"5c00", 864=>x"5c00", 865=>x"4a00", 866=>x"4600", 867=>x"4b00", 868=>x"5100",
---- 869=>x"5400", 870=>x"5c00", 871=>x"5a00", 872=>x"5e00", 873=>x"4c00", 874=>x"4900", 875=>x"4900",
---- 876=>x"5200", 877=>x"5800", 878=>x"5e00", 879=>x"5c00", 880=>x"5f00", 881=>x"4d00", 882=>x"4800",
---- 883=>x"4c00", 884=>x"5000", 885=>x"5400", 886=>x"5d00", 887=>x"5f00", 888=>x"6000", 889=>x"4c00",
---- 890=>x"4500", 891=>x"4d00", 892=>x"5100", 893=>x"5400", 894=>x"5e00", 895=>x"5c00", 896=>x"6200",
---- 897=>x"4d00", 898=>x"4600", 899=>x"4d00", 900=>x"4f00", 901=>x"5400", 902=>x"5b00", 903=>x"5e00",
---- 904=>x"6300", 905=>x"5100", 906=>x"4900", 907=>x"4d00", 908=>x"4f00", 909=>x"5300", 910=>x"5b00",
---- 911=>x"5b00", 912=>x"6300", 913=>x"5000", 914=>x"4700", 915=>x"4c00", 916=>x"5100", 917=>x"5700",
---- 918=>x"5d00", 919=>x"5e00", 920=>x"6400", 921=>x"5300", 922=>x"4a00", 923=>x"5300", 924=>x"5300",
---- 925=>x"5700", 926=>x"5e00", 927=>x"6100", 928=>x"6200", 929=>x"5200", 930=>x"4f00", 931=>x"5400",
---- 932=>x"5800", 933=>x"5a00", 934=>x"5f00", 935=>x"5e00", 936=>x"6200", 937=>x"4e00", 938=>x"4c00",
---- 939=>x"4e00", 940=>x"5900", 941=>x"5c00", 942=>x"5e00", 943=>x"6000", 944=>x"5f00", 945=>x"4d00",
---- 946=>x"4b00", 947=>x"4e00", 948=>x"5800", 949=>x"5b00", 950=>x"5f00", 951=>x"5f00", 952=>x"5e00",
---- 953=>x"5100", 954=>x"4d00", 955=>x"4f00", 956=>x"5500", 957=>x"5700", 958=>x"5e00", 959=>x"5f00",
---- 960=>x"6200", 961=>x"5100", 962=>x"4a00", 963=>x"4e00", 964=>x"5500", 965=>x"5600", 966=>x"5c00",
---- 967=>x"6000", 968=>x"6100", 969=>x"5000", 970=>x"4a00", 971=>x"4d00", 972=>x"5200", 973=>x"5900",
---- 974=>x"5d00", 975=>x"6000", 976=>x"5f00", 977=>x"5100", 978=>x"4900", 979=>x"5100", 980=>x"5400",
---- 981=>x"5700", 982=>x"5c00", 983=>x"5e00", 984=>x"6100", 985=>x"5200", 986=>x"4a00", 987=>x"5000",
---- 988=>x"5600", 989=>x"5600", 990=>x"5b00", 991=>x"5d00", 992=>x"5e00", 993=>x"4f00", 994=>x"4a00",
---- 995=>x"4f00", 996=>x"5500", 997=>x"5300", 998=>x"5e00", 999=>x"6000", 1000=>x"5f00", 1001=>x"4e00",
---- 1002=>x"4c00", 1003=>x"5000", 1004=>x"5500", 1005=>x"5800", 1006=>x"5b00", 1007=>x"6000", 1008=>x"5e00",
---- 1009=>x"4e00", 1010=>x"5100", 1011=>x"5300", 1012=>x"5500", 1013=>x"5900", 1014=>x"5e00", 1015=>x"6100",
---- 1016=>x"6400", 1017=>x"5000", 1018=>x"4a00", 1019=>x"5100", 1020=>x"5700", 1021=>x"5900", 1022=>x"5e00",
---- 1023=>x"6000", 1024=>x"6000", 1025=>x"4e00", 1026=>x"4a00", 1027=>x"4f00", 1028=>x"5300", 1029=>x"5300",
---- 1030=>x"5c00", 1031=>x"6100", 1032=>x"6300", 1033=>x"5100", 1034=>x"4c00", 1035=>x"4b00", 1036=>x"5200",
---- 1037=>x"5500", 1038=>x"5a00", 1039=>x"5e00", 1040=>x"6100", 1041=>x"5400", 1042=>x"4800", 1043=>x"4b00",
---- 1044=>x"5300", 1045=>x"5500", 1046=>x"5900", 1047=>x"5900", 1048=>x"6200", 1049=>x"4a00", 1050=>x"4700",
---- 1051=>x"4900", 1052=>x"5100", 1053=>x"5600", 1054=>x"5900", 1055=>x"a500", 1056=>x"6200", 1057=>x"4d00",
---- 1058=>x"4900", 1059=>x"4a00", 1060=>x"5300", 1061=>x"5800", 1062=>x"5d00", 1063=>x"5f00", 1064=>x"6100",
---- 1065=>x"4c00", 1066=>x"4900", 1067=>x"5000", 1068=>x"5600", 1069=>x"5a00", 1070=>x"6000", 1071=>x"6100",
---- 1072=>x"6500", 1073=>x"4f00", 1074=>x"4900", 1075=>x"5000", 1076=>x"5500", 1077=>x"5b00", 1078=>x"6200",
---- 1079=>x"6200", 1080=>x"6500", 1081=>x"5300", 1082=>x"4e00", 1083=>x"5300", 1084=>x"5600", 1085=>x"5c00",
---- 1086=>x"6200", 1087=>x"6100", 1088=>x"6900", 1089=>x"5300", 1090=>x"5000", 1091=>x"5400", 1092=>x"5a00",
---- 1093=>x"5e00", 1094=>x"6700", 1095=>x"6600", 1096=>x"6600", 1097=>x"5600", 1098=>x"5400", 1099=>x"5600",
---- 1100=>x"5a00", 1101=>x"5e00", 1102=>x"6300", 1103=>x"6600", 1104=>x"6600", 1105=>x"5700", 1106=>x"5200",
---- 1107=>x"5600", 1108=>x"5d00", 1109=>x"6000", 1110=>x"6600", 1111=>x"6900", 1112=>x"6a00", 1113=>x"aa00",
---- 1114=>x"5000", 1115=>x"5700", 1116=>x"5c00", 1117=>x"6300", 1118=>x"6600", 1119=>x"6900", 1120=>x"6c00",
---- 1121=>x"5500", 1122=>x"4f00", 1123=>x"5600", 1124=>x"5b00", 1125=>x"6100", 1126=>x"6500", 1127=>x"9600",
---- 1128=>x"6900", 1129=>x"5200", 1130=>x"4c00", 1131=>x"ac00", 1132=>x"5c00", 1133=>x"5e00", 1134=>x"6300",
---- 1135=>x"6700", 1136=>x"6800", 1137=>x"5300", 1138=>x"5000", 1139=>x"5500", 1140=>x"5c00", 1141=>x"5d00",
---- 1142=>x"6300", 1143=>x"6900", 1144=>x"6700", 1145=>x"5600", 1146=>x"4d00", 1147=>x"5500", 1148=>x"5900",
---- 1149=>x"5f00", 1150=>x"6400", 1151=>x"6800", 1152=>x"6900", 1153=>x"5700", 1154=>x"4f00", 1155=>x"5300",
---- 1156=>x"5a00", 1157=>x"5e00", 1158=>x"6300", 1159=>x"6800", 1160=>x"6700", 1161=>x"5600", 1162=>x"4e00",
---- 1163=>x"5200", 1164=>x"5b00", 1165=>x"5c00", 1166=>x"6200", 1167=>x"6300", 1168=>x"6900", 1169=>x"5200",
---- 1170=>x"4d00", 1171=>x"5300", 1172=>x"5900", 1173=>x"5a00", 1174=>x"6100", 1175=>x"6300", 1176=>x"6600",
---- 1177=>x"5100", 1178=>x"4e00", 1179=>x"5000", 1180=>x"5400", 1181=>x"5a00", 1182=>x"6300", 1183=>x"7500",
---- 1184=>x"9800", 1185=>x"5600", 1186=>x"4c00", 1187=>x"5300", 1188=>x"5a00", 1189=>x"5d00", 1190=>x"6600",
---- 1191=>x"7200", 1192=>x"6800", 1193=>x"5500", 1194=>x"4c00", 1195=>x"5500", 1196=>x"5900", 1197=>x"5f00",
---- 1198=>x"6400", 1199=>x"6800", 1200=>x"6900", 1201=>x"5300", 1202=>x"4d00", 1203=>x"5200", 1204=>x"5600",
---- 1205=>x"5b00", 1206=>x"6200", 1207=>x"6800", 1208=>x"6800", 1209=>x"5100", 1210=>x"4c00", 1211=>x"5400",
---- 1212=>x"5b00", 1213=>x"6100", 1214=>x"6000", 1215=>x"6300", 1216=>x"9700", 1217=>x"5200", 1218=>x"4800",
---- 1219=>x"4e00", 1220=>x"5d00", 1221=>x"7e00", 1222=>x"6b00", 1223=>x"6100", 1224=>x"6900", 1225=>x"4f00",
---- 1226=>x"4a00", 1227=>x"4900", 1228=>x"6100", 1229=>x"8800", 1230=>x"6200", 1231=>x"5c00", 1232=>x"6500",
---- 1233=>x"4d00", 1234=>x"4800", 1235=>x"4800", 1236=>x"5800", 1237=>x"8b00", 1238=>x"7300", 1239=>x"6000",
---- 1240=>x"6500", 1241=>x"4f00", 1242=>x"4800", 1243=>x"4a00", 1244=>x"b200", 1245=>x"7200", 1246=>x"9500",
---- 1247=>x"8600", 1248=>x"6400", 1249=>x"4f00", 1250=>x"4a00", 1251=>x"4a00", 1252=>x"4f00", 1253=>x"5b00",
---- 1254=>x"6e00", 1255=>x"7800", 1256=>x"6700", 1257=>x"5100", 1258=>x"4900", 1259=>x"4d00", 1260=>x"5200",
---- 1261=>x"5800", 1262=>x"5c00", 1263=>x"6f00", 1264=>x"6b00", 1265=>x"4f00", 1266=>x"4400", 1267=>x"4800",
---- 1268=>x"5500", 1269=>x"6b00", 1270=>x"8000", 1271=>x"7d00", 1272=>x"6800", 1273=>x"4e00", 1274=>x"4700",
---- 1275=>x"5800", 1276=>x"7800", 1277=>x"8c00", 1278=>x"7d00", 1279=>x"6700", 1280=>x"6d00", 1281=>x"5a00",
---- 1282=>x"6600", 1283=>x"7800", 1284=>x"7800", 1285=>x"6a00", 1286=>x"5f00", 1287=>x"6300", 1288=>x"6f00",
---- 1289=>x"6500", 1290=>x"5700", 1291=>x"5100", 1292=>x"5200", 1293=>x"5700", 1294=>x"5f00", 1295=>x"6500",
---- 1296=>x"7200", 1297=>x"5700", 1298=>x"4600", 1299=>x"4b00", 1300=>x"5500", 1301=>x"5b00", 1302=>x"5e00",
---- 1303=>x"6500", 1304=>x"6d00", 1305=>x"5300", 1306=>x"4900", 1307=>x"5000", 1308=>x"5600", 1309=>x"5b00",
---- 1310=>x"6100", 1311=>x"6400", 1312=>x"6d00", 1313=>x"5500", 1314=>x"4800", 1315=>x"4e00", 1316=>x"5600",
---- 1317=>x"5c00", 1318=>x"6100", 1319=>x"6400", 1320=>x"6c00", 1321=>x"5500", 1322=>x"4a00", 1323=>x"4e00",
---- 1324=>x"5500", 1325=>x"5a00", 1326=>x"5f00", 1327=>x"6000", 1328=>x"6d00", 1329=>x"5500", 1330=>x"4b00",
---- 1331=>x"5000", 1332=>x"5600", 1333=>x"5a00", 1334=>x"5d00", 1335=>x"6200", 1336=>x"6f00", 1337=>x"5500",
---- 1338=>x"4a00", 1339=>x"4e00", 1340=>x"5600", 1341=>x"5d00", 1342=>x"5e00", 1343=>x"6300", 1344=>x"6e00",
---- 1345=>x"5600", 1346=>x"4a00", 1347=>x"4d00", 1348=>x"5200", 1349=>x"5900", 1350=>x"5f00", 1351=>x"5e00",
---- 1352=>x"6d00", 1353=>x"5700", 1354=>x"4700", 1355=>x"4a00", 1356=>x"af00", 1357=>x"5800", 1358=>x"5d00",
---- 1359=>x"9b00", 1360=>x"6d00", 1361=>x"5500", 1362=>x"4600", 1363=>x"4b00", 1364=>x"ac00", 1365=>x"5500",
---- 1366=>x"5800", 1367=>x"7c00", 1368=>x"7000", 1369=>x"5300", 1370=>x"4500", 1371=>x"4c00", 1372=>x"5300",
---- 1373=>x"5400", 1374=>x"7200", 1375=>x"9100", 1376=>x"7200", 1377=>x"5300", 1378=>x"4500", 1379=>x"4b00",
---- 1380=>x"4e00", 1381=>x"6400", 1382=>x"9000", 1383=>x"7100", 1384=>x"6d00", 1385=>x"5300", 1386=>x"4800",
---- 1387=>x"4900", 1388=>x"5100", 1389=>x"8500", 1390=>x"7e00", 1391=>x"5900", 1392=>x"6c00", 1393=>x"5200",
---- 1394=>x"4500", 1395=>x"4900", 1396=>x"7000", 1397=>x"8800", 1398=>x"5e00", 1399=>x"5a00", 1400=>x"6d00",
---- 1401=>x"5200", 1402=>x"3f00", 1403=>x"6b00", 1404=>x"9300", 1405=>x"6900", 1406=>x"5500", 1407=>x"5900",
---- 1408=>x"6e00", 1409=>x"5000", 1410=>x"5b00", 1411=>x"9500", 1412=>x"7600", 1413=>x"5200", 1414=>x"5300",
---- 1415=>x"5e00", 1416=>x"6800", 1417=>x"6600", 1418=>x"9800", 1419=>x"7f00", 1420=>x"4d00", 1421=>x"5000",
---- 1422=>x"5700", 1423=>x"7300", 1424=>x"7800", 1425=>x"9800", 1426=>x"8500", 1427=>x"4e00", 1428=>x"4c00",
---- 1429=>x"5100", 1430=>x"5d00", 1431=>x"8900", 1432=>x"9000", 1433=>x"7c00", 1434=>x"4c00", 1435=>x"4400",
---- 1436=>x"4c00", 1437=>x"5100", 1438=>x"6d00", 1439=>x"9600", 1440=>x"7b00", 1441=>x"5300", 1442=>x"3e00",
---- 1443=>x"4600", 1444=>x"4b00", 1445=>x"5c00", 1446=>x"9100", 1447=>x"8900", 1448=>x"6900", 1449=>x"4d00",
---- 1450=>x"4400", 1451=>x"4800", 1452=>x"5000", 1453=>x"8100", 1454=>x"9900", 1455=>x"6900", 1456=>x"6900",
---- 1457=>x"4f00", 1458=>x"4300", 1459=>x"4200", 1460=>x"5d00", 1461=>x"9900", 1462=>x"7700", 1463=>x"5f00",
---- 1464=>x"6a00", 1465=>x"b000", 1466=>x"4100", 1467=>x"4300", 1468=>x"6600", 1469=>x"9800", 1470=>x"6400",
---- 1471=>x"6200", 1472=>x"6e00", 1473=>x"4f00", 1474=>x"4000", 1475=>x"4200", 1476=>x"6800", 1477=>x"9400",
---- 1478=>x"6200", 1479=>x"6000", 1480=>x"6d00", 1481=>x"5100", 1482=>x"4100", 1483=>x"4300", 1484=>x"5e00",
---- 1485=>x"8900", 1486=>x"6d00", 1487=>x"6100", 1488=>x"6e00", 1489=>x"5800", 1490=>x"4500", 1491=>x"4400",
---- 1492=>x"5300", 1493=>x"7600", 1494=>x"7600", 1495=>x"6b00", 1496=>x"6c00", 1497=>x"5500", 1498=>x"4300",
---- 1499=>x"4400", 1500=>x"5300", 1501=>x"6700", 1502=>x"6c00", 1503=>x"6600", 1504=>x"6c00", 1505=>x"5200",
---- 1506=>x"4100", 1507=>x"4900", 1508=>x"5400", 1509=>x"6500", 1510=>x"6600", 1511=>x"6600", 1512=>x"6f00",
---- 1513=>x"5200", 1514=>x"4300", 1515=>x"4800", 1516=>x"5300", 1517=>x"6200", 1518=>x"6600", 1519=>x"5c00",
---- 1520=>x"6c00", 1521=>x"4f00", 1522=>x"4200", 1523=>x"4600", 1524=>x"5200", 1525=>x"5f00", 1526=>x"7600",
---- 1527=>x"4800", 1528=>x"6c00", 1529=>x"4d00", 1530=>x"3e00", 1531=>x"4200", 1532=>x"4700", 1533=>x"6a00",
---- 1534=>x"6200", 1535=>x"3500", 1536=>x"6a00", 1537=>x"4d00", 1538=>x"3900", 1539=>x"3b00", 1540=>x"6100",
---- 1541=>x"8200", 1542=>x"5200", 1543=>x"5600", 1544=>x"6600", 1545=>x"4500", 1546=>x"3800", 1547=>x"6900",
---- 1548=>x"b800", 1549=>x"8b00", 1550=>x"5f00", 1551=>x"9000", 1552=>x"5f00", 1553=>x"4800", 1554=>x"7900",
---- 1555=>x"cf00", 1556=>x"9a00", 1557=>x"4500", 1558=>x"6000", 1559=>x"9100", 1560=>x"6100", 1561=>x"8800",
---- 1562=>x"d700", 1563=>x"9900", 1564=>x"5300", 1565=>x"4000", 1566=>x"6300", 1567=>x"8400", 1568=>x"9c00",
---- 1569=>x"d400", 1570=>x"9100", 1571=>x"3e00", 1572=>x"5600", 1573=>x"3c00", 1574=>x"5800", 1575=>x"5c00",
---- 1576=>x"c400", 1577=>x"7a00", 1578=>x"3700", 1579=>x"5100", 1580=>x"4100", 1581=>x"3400", 1582=>x"8700",
---- 1583=>x"4700", 1584=>x"7a00", 1585=>x"4000", 1586=>x"4100", 1587=>x"4f00", 1588=>x"3900", 1589=>x"7100",
---- 1590=>x"9700", 1591=>x"3000", 1592=>x"6300", 1593=>x"4c00", 1594=>x"4100", 1595=>x"5700", 1596=>x"6600",
---- 1597=>x"9700", 1598=>x"5a00", 1599=>x"2400", 1600=>x"6c00", 1601=>x"4c00", 1602=>x"5400", 1603=>x"7100",
---- 1604=>x"a800", 1605=>x"7100", 1606=>x"2a00", 1607=>x"2800", 1608=>x"6700", 1609=>x"5600", 1610=>x"7500",
---- 1611=>x"8200", 1612=>x"bd00", 1613=>x"3f00", 1614=>x"2900", 1615=>x"2a00", 1616=>x"7200", 1617=>x"7c00",
---- 1618=>x"8600", 1619=>x"7d00", 1620=>x"9200", 1621=>x"2900", 1622=>x"2b00", 1623=>x"2a00", 1624=>x"8900",
---- 1625=>x"ae00", 1626=>x"8000", 1627=>x"7300", 1628=>x"5d00", 1629=>x"2700", 1630=>x"2c00", 1631=>x"2d00",
---- 1632=>x"4400", 1633=>x"c200", 1634=>x"5e00", 1635=>x"6100", 1636=>x"5700", 1637=>x"3800", 1638=>x"2e00",
---- 1639=>x"2800", 1640=>x"de00", 1641=>x"a700", 1642=>x"5b00", 1643=>x"5700", 1644=>x"4200", 1645=>x"3c00",
---- 1646=>x"3800", 1647=>x"2e00", 1648=>x"de00", 1649=>x"9000", 1650=>x"8200", 1651=>x"9200", 1652=>x"3000",
---- 1653=>x"2500", 1654=>x"2d00", 1655=>x"2f00", 1656=>x"cd00", 1657=>x"7700", 1658=>x"5b00", 1659=>x"9e00",
---- 1660=>x"2b00", 1661=>x"2300", 1662=>x"2900", 1663=>x"2d00", 1664=>x"a800", 1665=>x"7600", 1666=>x"4f00",
---- 1667=>x"4c00", 1668=>x"2500", 1669=>x"2700", 1670=>x"2f00", 1671=>x"2c00", 1672=>x"b300", 1673=>x"7800",
---- 1674=>x"5a00", 1675=>x"3a00", 1676=>x"2a00", 1677=>x"2900", 1678=>x"2b00", 1679=>x"2c00", 1680=>x"c000",
---- 1681=>x"7700", 1682=>x"5600", 1683=>x"5a00", 1684=>x"2700", 1685=>x"2700", 1686=>x"2c00", 1687=>x"2900",
---- 1688=>x"8100", 1689=>x"9200", 1690=>x"6d00", 1691=>x"6500", 1692=>x"1f00", 1693=>x"2600", 1694=>x"3100",
---- 1695=>x"2a00", 1696=>x"6d00", 1697=>x"ab00", 1698=>x"a200", 1699=>x"3700", 1700=>x"2700", 1701=>x"2d00",
---- 1702=>x"2f00", 1703=>x"2900", 1704=>x"6d00", 1705=>x"7100", 1706=>x"7700", 1707=>x"4100", 1708=>x"2200",
---- 1709=>x"3100", 1710=>x"2e00", 1711=>x"2900", 1712=>x"7800", 1713=>x"8e00", 1714=>x"9200", 1715=>x"3d00",
---- 1716=>x"2d00", 1717=>x"3300", 1718=>x"2f00", 1719=>x"2c00", 1720=>x"9800", 1721=>x"9100", 1722=>x"6700",
---- 1723=>x"2b00", 1724=>x"3500", 1725=>x"3100", 1726=>x"2600", 1727=>x"3200", 1728=>x"9e00", 1729=>x"8c00",
---- 1730=>x"5c00", 1731=>x"2c00", 1732=>x"3500", 1733=>x"2d00", 1734=>x"2b00", 1735=>x"4000", 1736=>x"9500",
---- 1737=>x"7d00", 1738=>x"3300", 1739=>x"2a00", 1740=>x"3400", 1741=>x"2f00", 1742=>x"3800", 1743=>x"3b00",
---- 1744=>x"8d00", 1745=>x"7600", 1746=>x"2a00", 1747=>x"2d00", 1748=>x"3800", 1749=>x"3c00", 1750=>x"3d00",
---- 1751=>x"2a00", 1752=>x"8400", 1753=>x"7000", 1754=>x"3500", 1755=>x"3800", 1756=>x"4300", 1757=>x"3500",
---- 1758=>x"3000", 1759=>x"2800", 1760=>x"7e00", 1761=>x"6900", 1762=>x"4300", 1763=>x"3e00", 1764=>x"4000",
---- 1765=>x"2d00", 1766=>x"2b00", 1767=>x"2b00", 1768=>x"8000", 1769=>x"7f00", 1770=>x"5100", 1771=>x"3100",
---- 1772=>x"3500", 1773=>x"2d00", 1774=>x"2d00", 1775=>x"2e00", 1776=>x"8a00", 1777=>x"8a00", 1778=>x"4c00",
---- 1779=>x"3f00", 1780=>x"2c00", 1781=>x"2b00", 1782=>x"2e00", 1783=>x"2e00", 1784=>x"9400", 1785=>x"6f00",
---- 1786=>x"4400", 1787=>x"3d00", 1788=>x"2d00", 1789=>x"3100", 1790=>x"2b00", 1791=>x"3400", 1792=>x"9100",
---- 1793=>x"6900", 1794=>x"3d00", 1795=>x"2f00", 1796=>x"2e00", 1797=>x"3900", 1798=>x"3100", 1799=>x"2e00",
---- 1800=>x"9800", 1801=>x"6d00", 1802=>x"4000", 1803=>x"3500", 1804=>x"2e00", 1805=>x"3800", 1806=>x"3000",
---- 1807=>x"2b00", 1808=>x"9c00", 1809=>x"7e00", 1810=>x"4600", 1811=>x"3700", 1812=>x"3200", 1813=>x"3200",
---- 1814=>x"2f00", 1815=>x"2b00", 1816=>x"9f00", 1817=>x"8600", 1818=>x"4000", 1819=>x"4a00", 1820=>x"3b00",
---- 1821=>x"3100", 1822=>x"2a00", 1823=>x"2900", 1824=>x"a400", 1825=>x"8700", 1826=>x"4300", 1827=>x"5800",
---- 1828=>x"4000", 1829=>x"2e00", 1830=>x"2600", 1831=>x"2900", 1832=>x"9b00", 1833=>x"9100", 1834=>x"4500",
---- 1835=>x"5800", 1836=>x"4000", 1837=>x"3000", 1838=>x"2c00", 1839=>x"2e00", 1840=>x"8d00", 1841=>x"8c00",
---- 1842=>x"4500", 1843=>x"5100", 1844=>x"3d00", 1845=>x"3600", 1846=>x"2b00", 1847=>x"2a00", 1848=>x"8100",
---- 1849=>x"7f00", 1850=>x"5000", 1851=>x"5600", 1852=>x"4400", 1853=>x"3200", 1854=>x"d800", 1855=>x"2d00",
---- 1856=>x"7f00", 1857=>x"7300", 1858=>x"5400", 1859=>x"5200", 1860=>x"5200", 1861=>x"2b00", 1862=>x"2600",
---- 1863=>x"2d00", 1864=>x"8100", 1865=>x"7200", 1866=>x"5800", 1867=>x"5000", 1868=>x"5a00", 1869=>x"2d00",
---- 1870=>x"2800", 1871=>x"3000", 1872=>x"6e00", 1873=>x"7100", 1874=>x"6300", 1875=>x"5400", 1876=>x"5700",
---- 1877=>x"2800", 1878=>x"2600", 1879=>x"3500", 1880=>x"5100", 1881=>x"7000", 1882=>x"6700", 1883=>x"5500",
---- 1884=>x"5400", 1885=>x"2600", 1886=>x"2e00", 1887=>x"3800", 1888=>x"5000", 1889=>x"7500", 1890=>x"6100",
---- 1891=>x"4400", 1892=>x"4200", 1893=>x"2800", 1894=>x"3300", 1895=>x"3100", 1896=>x"5700", 1897=>x"7d00",
---- 1898=>x"6c00", 1899=>x"3900", 1900=>x"3800", 1901=>x"2c00", 1902=>x"3200", 1903=>x"2e00", 1904=>x"5f00",
---- 1905=>x"8100", 1906=>x"7200", 1907=>x"3f00", 1908=>x"3200", 1909=>x"2b00", 1910=>x"3500", 1911=>x"3100",
---- 1912=>x"6700", 1913=>x"7d00", 1914=>x"6a00", 1915=>x"4c00", 1916=>x"2700", 1917=>x"2a00", 1918=>x"2f00",
---- 1919=>x"3500", 1920=>x"6700", 1921=>x"7a00", 1922=>x"6300", 1923=>x"4e00", 1924=>x"3000", 1925=>x"2c00",
---- 1926=>x"3100", 1927=>x"2e00", 1928=>x"6a00", 1929=>x"8500", 1930=>x"6000", 1931=>x"4400", 1932=>x"2b00",
---- 1933=>x"3300", 1934=>x"2f00", 1935=>x"2d00", 1936=>x"6d00", 1937=>x"7a00", 1938=>x"5b00", 1939=>x"3800",
---- 1940=>x"2700", 1941=>x"3500", 1942=>x"2f00", 1943=>x"3300", 1944=>x"6400", 1945=>x"7a00", 1946=>x"6400",
---- 1947=>x"3200", 1948=>x"2a00", 1949=>x"3100", 1950=>x"2a00", 1951=>x"3600", 1952=>x"5600", 1953=>x"7300",
---- 1954=>x"5c00", 1955=>x"2d00", 1956=>x"2600", 1957=>x"2e00", 1958=>x"2c00", 1959=>x"3500", 1960=>x"5400",
---- 1961=>x"6400", 1962=>x"5100", 1963=>x"2900", 1964=>x"2c00", 1965=>x"2c00", 1966=>x"3200", 1967=>x"3500",
---- 1968=>x"4900", 1969=>x"5100", 1970=>x"3d00", 1971=>x"2b00", 1972=>x"3100", 1973=>x"2900", 1974=>x"2a00",
---- 1975=>x"3000", 1976=>x"4500", 1977=>x"4900", 1978=>x"3400", 1979=>x"d500", 1980=>x"3000", 1981=>x"2b00",
---- 1982=>x"3600", 1983=>x"3200", 1984=>x"4600", 1985=>x"4700", 1986=>x"3900", 1987=>x"3200", 1988=>x"3000",
---- 1989=>x"2f00", 1990=>x"3b00", 1991=>x"3600", 1992=>x"4100", 1993=>x"4100", 1994=>x"4300", 1995=>x"3d00",
---- 1996=>x"3000", 1997=>x"2e00", 1998=>x"2f00", 1999=>x"3000", 2000=>x"3400", 2001=>x"3b00", 2002=>x"3a00",
---- 2003=>x"3600", 2004=>x"2d00", 2005=>x"3300", 2006=>x"3600", 2007=>x"2d00", 2008=>x"4700", 2009=>x"3a00",
---- 2010=>x"3300", 2011=>x"3200", 2012=>x"3a00", 2013=>x"2e00", 2014=>x"3300", 2015=>x"2d00", 2016=>x"5c00",
---- 2017=>x"3a00", 2018=>x"2e00", 2019=>x"3100", 2020=>x"3e00", 2021=>x"2f00", 2022=>x"3800", 2023=>x"2f00",
---- 2024=>x"5500", 2025=>x"3300", 2026=>x"3200", 2027=>x"2e00", 2028=>x"3100", 2029=>x"2b00", 2030=>x"3700",
---- 2031=>x"3300", 2032=>x"4700", 2033=>x"3600", 2034=>x"3c00", 2035=>x"2b00", 2036=>x"2800", 2037=>x"2e00",
---- 2038=>x"3e00", 2039=>x"2e00", 2040=>x"4600", 2041=>x"3900", 2042=>x"3800", 2043=>x"2800", 2044=>x"2600",
---- 2045=>x"3300", 2046=>x"4400", 2047=>x"2700"),
---- 5  => (0=>x"6d00", 1=>x"6a00", 2=>x"6900", 3=>x"6d00", 4=>x"6c00", 5=>x"6a00", 6=>x"6d00", 7=>x"6c00",
---- 8=>x"6e00", 9=>x"6a00", 10=>x"6900", 11=>x"6e00", 12=>x"6c00", 13=>x"6b00", 14=>x"6d00",
---- 15=>x"6b00", 16=>x"6d00", 17=>x"6a00", 18=>x"6800", 19=>x"6c00", 20=>x"6b00", 21=>x"6a00",
---- 22=>x"6d00", 23=>x"6b00", 24=>x"6700", 25=>x"6800", 26=>x"6700", 27=>x"6800", 28=>x"6700",
---- 29=>x"6800", 30=>x"6900", 31=>x"6800", 32=>x"9500", 33=>x"6900", 34=>x"6500", 35=>x"6a00",
---- 36=>x"6900", 37=>x"6800", 38=>x"6800", 39=>x"6700", 40=>x"9b00", 41=>x"6600", 42=>x"6700",
---- 43=>x"6700", 44=>x"6800", 45=>x"6b00", 46=>x"6700", 47=>x"6600", 48=>x"6600", 49=>x"6900",
---- 50=>x"6a00", 51=>x"6b00", 52=>x"6c00", 53=>x"6900", 54=>x"6600", 55=>x"6700", 56=>x"6900",
---- 57=>x"6e00", 58=>x"6b00", 59=>x"6b00", 60=>x"6b00", 61=>x"6b00", 62=>x"6600", 63=>x"6800",
---- 64=>x"6a00", 65=>x"6a00", 66=>x"6900", 67=>x"6a00", 68=>x"6700", 69=>x"9700", 70=>x"6700",
---- 71=>x"6a00", 72=>x"6600", 73=>x"6700", 74=>x"6a00", 75=>x"6b00", 76=>x"6900", 77=>x"6a00",
---- 78=>x"6900", 79=>x"6a00", 80=>x"6b00", 81=>x"6c00", 82=>x"6b00", 83=>x"6c00", 84=>x"6800",
---- 85=>x"6800", 86=>x"6600", 87=>x"6500", 88=>x"7000", 89=>x"6700", 90=>x"6700", 91=>x"6700",
---- 92=>x"6700", 93=>x"9500", 94=>x"6500", 95=>x"6600", 96=>x"6a00", 97=>x"6800", 98=>x"6900",
---- 99=>x"6600", 100=>x"6400", 101=>x"6a00", 102=>x"6700", 103=>x"6800", 104=>x"6900", 105=>x"6900",
---- 106=>x"6900", 107=>x"6900", 108=>x"6900", 109=>x"6a00", 110=>x"6600", 111=>x"6600", 112=>x"6700",
---- 113=>x"6800", 114=>x"6800", 115=>x"6b00", 116=>x"6a00", 117=>x"6900", 118=>x"6800", 119=>x"6700",
---- 120=>x"6b00", 121=>x"6b00", 122=>x"6c00", 123=>x"6700", 124=>x"6900", 125=>x"6a00", 126=>x"6600",
---- 127=>x"6700", 128=>x"6900", 129=>x"6b00", 130=>x"6c00", 131=>x"6c00", 132=>x"6b00", 133=>x"6a00",
---- 134=>x"6400", 135=>x"6600", 136=>x"6800", 137=>x"6900", 138=>x"6800", 139=>x"6a00", 140=>x"6900",
---- 141=>x"6700", 142=>x"6700", 143=>x"6700", 144=>x"6800", 145=>x"6700", 146=>x"6600", 147=>x"6500",
---- 148=>x"6700", 149=>x"6700", 150=>x"6700", 151=>x"6400", 152=>x"6600", 153=>x"6900", 154=>x"6500",
---- 155=>x"6500", 156=>x"6600", 157=>x"6800", 158=>x"6600", 159=>x"6600", 160=>x"6700", 161=>x"6700",
---- 162=>x"6400", 163=>x"6700", 164=>x"6600", 165=>x"6500", 166=>x"6500", 167=>x"6700", 168=>x"6700",
---- 169=>x"9a00", 170=>x"6600", 171=>x"6700", 172=>x"6600", 173=>x"6a00", 174=>x"6400", 175=>x"9800",
---- 176=>x"6700", 177=>x"6600", 178=>x"6900", 179=>x"6700", 180=>x"6700", 181=>x"6800", 182=>x"6a00",
---- 183=>x"6600", 184=>x"6800", 185=>x"6900", 186=>x"6900", 187=>x"6b00", 188=>x"6700", 189=>x"6600",
---- 190=>x"6900", 191=>x"6700", 192=>x"6700", 193=>x"6900", 194=>x"6900", 195=>x"6c00", 196=>x"6700",
---- 197=>x"6600", 198=>x"6800", 199=>x"6600", 200=>x"6700", 201=>x"6700", 202=>x"6600", 203=>x"6700",
---- 204=>x"6600", 205=>x"6400", 206=>x"6700", 207=>x"6900", 208=>x"6800", 209=>x"6900", 210=>x"6700",
---- 211=>x"6800", 212=>x"6600", 213=>x"6a00", 214=>x"6700", 215=>x"6600", 216=>x"6500", 217=>x"6900",
---- 218=>x"6500", 219=>x"6500", 220=>x"6800", 221=>x"6900", 222=>x"6600", 223=>x"6700", 224=>x"6300",
---- 225=>x"6400", 226=>x"6800", 227=>x"6300", 228=>x"6600", 229=>x"6600", 230=>x"6700", 231=>x"6500",
---- 232=>x"5f00", 233=>x"6100", 234=>x"6300", 235=>x"6600", 236=>x"6500", 237=>x"6300", 238=>x"9b00",
---- 239=>x"6200", 240=>x"6500", 241=>x"6500", 242=>x"6400", 243=>x"9d00", 244=>x"6300", 245=>x"6500",
---- 246=>x"6100", 247=>x"6400", 248=>x"6100", 249=>x"6400", 250=>x"6100", 251=>x"5f00", 252=>x"6300",
---- 253=>x"6200", 254=>x"6200", 255=>x"6500", 256=>x"5f00", 257=>x"5e00", 258=>x"5d00", 259=>x"6200",
---- 260=>x"6400", 261=>x"6300", 262=>x"6300", 263=>x"6300", 264=>x"5e00", 265=>x"5f00", 266=>x"5f00",
---- 267=>x"6200", 268=>x"6100", 269=>x"6300", 270=>x"6400", 271=>x"6500", 272=>x"5f00", 273=>x"6100",
---- 274=>x"6200", 275=>x"6100", 276=>x"6200", 277=>x"6500", 278=>x"6300", 279=>x"6300", 280=>x"6400",
---- 281=>x"6700", 282=>x"6600", 283=>x"6900", 284=>x"6300", 285=>x"6500", 286=>x"6500", 287=>x"6300",
---- 288=>x"6400", 289=>x"6500", 290=>x"6000", 291=>x"6700", 292=>x"6600", 293=>x"6400", 294=>x"6100",
---- 295=>x"9d00", 296=>x"6100", 297=>x"6200", 298=>x"6100", 299=>x"6600", 300=>x"6400", 301=>x"6600",
---- 302=>x"9c00", 303=>x"6300", 304=>x"6500", 305=>x"6200", 306=>x"6200", 307=>x"6400", 308=>x"6200",
---- 309=>x"6400", 310=>x"6300", 311=>x"6500", 312=>x"6900", 313=>x"6200", 314=>x"6300", 315=>x"6400",
---- 316=>x"9b00", 317=>x"6100", 318=>x"6500", 319=>x"6200", 320=>x"6100", 321=>x"6000", 322=>x"6000",
---- 323=>x"6100", 324=>x"6600", 325=>x"6400", 326=>x"6200", 327=>x"6400", 328=>x"5f00", 329=>x"6500",
---- 330=>x"6900", 331=>x"6000", 332=>x"6400", 333=>x"6500", 334=>x"6300", 335=>x"6300", 336=>x"6100",
---- 337=>x"6300", 338=>x"6300", 339=>x"6300", 340=>x"6300", 341=>x"6000", 342=>x"6800", 343=>x"6700",
---- 344=>x"6000", 345=>x"6300", 346=>x"6300", 347=>x"6300", 348=>x"6200", 349=>x"6400", 350=>x"6a00",
---- 351=>x"6700", 352=>x"5f00", 353=>x"5e00", 354=>x"6200", 355=>x"6600", 356=>x"6600", 357=>x"6600",
---- 358=>x"6900", 359=>x"6500", 360=>x"5f00", 361=>x"5e00", 362=>x"6500", 363=>x"6700", 364=>x"6500",
---- 365=>x"6500", 366=>x"6900", 367=>x"6600", 368=>x"6100", 369=>x"5f00", 370=>x"6200", 371=>x"6300",
---- 372=>x"6200", 373=>x"6300", 374=>x"6500", 375=>x"9c00", 376=>x"6700", 377=>x"6200", 378=>x"6100",
---- 379=>x"6100", 380=>x"6300", 381=>x"6200", 382=>x"6600", 383=>x"9e00", 384=>x"6400", 385=>x"6600",
---- 386=>x"6100", 387=>x"6300", 388=>x"6400", 389=>x"6400", 390=>x"6300", 391=>x"6600", 392=>x"6300",
---- 393=>x"6300", 394=>x"6300", 395=>x"6500", 396=>x"6200", 397=>x"6100", 398=>x"6200", 399=>x"6200",
---- 400=>x"6000", 401=>x"6600", 402=>x"6300", 403=>x"6400", 404=>x"6200", 405=>x"6500", 406=>x"6100",
---- 407=>x"6400", 408=>x"6200", 409=>x"6200", 410=>x"6200", 411=>x"6100", 412=>x"6200", 413=>x"6600",
---- 414=>x"6300", 415=>x"6400", 416=>x"6100", 417=>x"6000", 418=>x"6000", 419=>x"6600", 420=>x"6700",
---- 421=>x"6500", 422=>x"6300", 423=>x"6300", 424=>x"5f00", 425=>x"6000", 426=>x"6100", 427=>x"6100",
---- 428=>x"6900", 429=>x"6600", 430=>x"6300", 431=>x"6200", 432=>x"6000", 433=>x"6200", 434=>x"6400",
---- 435=>x"6200", 436=>x"6500", 437=>x"6400", 438=>x"6600", 439=>x"6400", 440=>x"5f00", 441=>x"6300",
---- 442=>x"6300", 443=>x"6200", 444=>x"6500", 445=>x"6400", 446=>x"6500", 447=>x"6600", 448=>x"5e00",
---- 449=>x"6100", 450=>x"5d00", 451=>x"6200", 452=>x"6400", 453=>x"6600", 454=>x"6a00", 455=>x"6500",
---- 456=>x"5c00", 457=>x"5d00", 458=>x"6100", 459=>x"6300", 460=>x"6500", 461=>x"6200", 462=>x"6600",
---- 463=>x"6300", 464=>x"5c00", 465=>x"5f00", 466=>x"5f00", 467=>x"5f00", 468=>x"6100", 469=>x"6000",
---- 470=>x"5f00", 471=>x"6000", 472=>x"5e00", 473=>x"5d00", 474=>x"5f00", 475=>x"6000", 476=>x"5f00",
---- 477=>x"6100", 478=>x"6000", 479=>x"5e00", 480=>x"5d00", 481=>x"6100", 482=>x"6200", 483=>x"6200",
---- 484=>x"6100", 485=>x"6200", 486=>x"6200", 487=>x"5f00", 488=>x"5b00", 489=>x"5e00", 490=>x"6200",
---- 491=>x"6200", 492=>x"6200", 493=>x"6500", 494=>x"6300", 495=>x"6300", 496=>x"5e00", 497=>x"6200",
---- 498=>x"6400", 499=>x"6300", 500=>x"6100", 501=>x"6500", 502=>x"6400", 503=>x"6300", 504=>x"6200",
---- 505=>x"6500", 506=>x"6400", 507=>x"6300", 508=>x"6300", 509=>x"6600", 510=>x"6600", 511=>x"6300",
---- 512=>x"6100", 513=>x"6100", 514=>x"6200", 515=>x"6300", 516=>x"6300", 517=>x"6600", 518=>x"6600",
---- 519=>x"6300", 520=>x"6100", 521=>x"6400", 522=>x"6300", 523=>x"6500", 524=>x"6400", 525=>x"6500",
---- 526=>x"6500", 527=>x"6500", 528=>x"6300", 529=>x"6500", 530=>x"6300", 531=>x"6700", 532=>x"6600",
---- 533=>x"6400", 534=>x"6800", 535=>x"6a00", 536=>x"6200", 537=>x"6200", 538=>x"6300", 539=>x"6700",
---- 540=>x"6600", 541=>x"6700", 542=>x"6900", 543=>x"6a00", 544=>x"6500", 545=>x"6600", 546=>x"6200",
---- 547=>x"6400", 548=>x"6500", 549=>x"6600", 550=>x"6500", 551=>x"6600", 552=>x"6300", 553=>x"6500",
---- 554=>x"6400", 555=>x"6600", 556=>x"6500", 557=>x"6800", 558=>x"6100", 559=>x"6500", 560=>x"6200",
---- 561=>x"6200", 562=>x"6100", 563=>x"6600", 564=>x"6600", 565=>x"6500", 566=>x"6500", 567=>x"6600",
---- 568=>x"6400", 569=>x"6300", 570=>x"6100", 571=>x"6200", 572=>x"6600", 573=>x"6400", 574=>x"6500",
---- 575=>x"6500", 576=>x"6100", 577=>x"6400", 578=>x"6300", 579=>x"6400", 580=>x"6300", 581=>x"6400",
---- 582=>x"6300", 583=>x"6400", 584=>x"5e00", 585=>x"6300", 586=>x"6400", 587=>x"6500", 588=>x"6400",
---- 589=>x"6100", 590=>x"6300", 591=>x"6200", 592=>x"5d00", 593=>x"5f00", 594=>x"6200", 595=>x"6700",
---- 596=>x"6500", 597=>x"6300", 598=>x"6200", 599=>x"6100", 600=>x"6000", 601=>x"6300", 602=>x"6000",
---- 603=>x"6200", 604=>x"6100", 605=>x"6300", 606=>x"6200", 607=>x"6400", 608=>x"5f00", 609=>x"6300",
---- 610=>x"6300", 611=>x"6300", 612=>x"6100", 613=>x"6300", 614=>x"6500", 615=>x"6100", 616=>x"5f00",
---- 617=>x"6400", 618=>x"6400", 619=>x"6400", 620=>x"6400", 621=>x"9f00", 622=>x"6400", 623=>x"6300",
---- 624=>x"5f00", 625=>x"6300", 626=>x"6700", 627=>x"9a00", 628=>x"6400", 629=>x"6000", 630=>x"6200",
---- 631=>x"6400", 632=>x"9d00", 633=>x"6600", 634=>x"6300", 635=>x"6100", 636=>x"6300", 637=>x"6200",
---- 638=>x"6300", 639=>x"6300", 640=>x"6200", 641=>x"6600", 642=>x"6300", 643=>x"6200", 644=>x"6200",
---- 645=>x"6400", 646=>x"6200", 647=>x"6200", 648=>x"6000", 649=>x"6300", 650=>x"6300", 651=>x"6300",
---- 652=>x"6300", 653=>x"5f00", 654=>x"5f00", 655=>x"6200", 656=>x"6200", 657=>x"6200", 658=>x"6200",
---- 659=>x"6200", 660=>x"6200", 661=>x"6000", 662=>x"6200", 663=>x"6200", 664=>x"6300", 665=>x"6100",
---- 666=>x"6300", 667=>x"6000", 668=>x"6300", 669=>x"6200", 670=>x"6400", 671=>x"6200", 672=>x"5f00",
---- 673=>x"6300", 674=>x"6000", 675=>x"5f00", 676=>x"6200", 677=>x"6000", 678=>x"6000", 679=>x"6100",
---- 680=>x"5c00", 681=>x"6100", 682=>x"6300", 683=>x"6100", 684=>x"6000", 685=>x"5d00", 686=>x"6100",
---- 687=>x"6300", 688=>x"6400", 689=>x"6000", 690=>x"6200", 691=>x"6100", 692=>x"5e00", 693=>x"5d00",
---- 694=>x"6200", 695=>x"6000", 696=>x"6300", 697=>x"6000", 698=>x"6100", 699=>x"6100", 700=>x"6200",
---- 701=>x"6300", 702=>x"6100", 703=>x"6100", 704=>x"6100", 705=>x"6400", 706=>x"6000", 707=>x"6200",
---- 708=>x"6500", 709=>x"6200", 710=>x"6100", 711=>x"6500", 712=>x"5d00", 713=>x"5f00", 714=>x"6000",
---- 715=>x"6400", 716=>x"6600", 717=>x"6400", 718=>x"6000", 719=>x"6700", 720=>x"6200", 721=>x"6000",
---- 722=>x"6200", 723=>x"6300", 724=>x"6600", 725=>x"6100", 726=>x"6100", 727=>x"6600", 728=>x"5e00",
---- 729=>x"6300", 730=>x"6300", 731=>x"6100", 732=>x"6100", 733=>x"6200", 734=>x"6300", 735=>x"6600",
---- 736=>x"6000", 737=>x"6000", 738=>x"6200", 739=>x"6200", 740=>x"6100", 741=>x"6200", 742=>x"6500",
---- 743=>x"6400", 744=>x"5f00", 745=>x"6000", 746=>x"6300", 747=>x"6200", 748=>x"6400", 749=>x"6200",
---- 750=>x"6300", 751=>x"6500", 752=>x"5e00", 753=>x"6100", 754=>x"6500", 755=>x"6200", 756=>x"6200",
---- 757=>x"6200", 758=>x"6200", 759=>x"6500", 760=>x"6000", 761=>x"5f00", 762=>x"6000", 763=>x"5f00",
---- 764=>x"6100", 765=>x"6200", 766=>x"6400", 767=>x"6500", 768=>x"5e00", 769=>x"5e00", 770=>x"5f00",
---- 771=>x"6200", 772=>x"6200", 773=>x"5f00", 774=>x"6300", 775=>x"6300", 776=>x"6000", 777=>x"6000",
---- 778=>x"5f00", 779=>x"6400", 780=>x"6200", 781=>x"6300", 782=>x"6200", 783=>x"9d00", 784=>x"5f00",
---- 785=>x"6000", 786=>x"5f00", 787=>x"6100", 788=>x"6500", 789=>x"6400", 790=>x"6500", 791=>x"6500",
---- 792=>x"5e00", 793=>x"6000", 794=>x"5f00", 795=>x"6000", 796=>x"6300", 797=>x"6100", 798=>x"6300",
---- 799=>x"6300", 800=>x"5d00", 801=>x"6000", 802=>x"6000", 803=>x"5f00", 804=>x"6000", 805=>x"5f00",
---- 806=>x"6400", 807=>x"6600", 808=>x"5e00", 809=>x"5e00", 810=>x"a100", 811=>x"6000", 812=>x"6000",
---- 813=>x"6100", 814=>x"5f00", 815=>x"6000", 816=>x"5e00", 817=>x"5e00", 818=>x"6200", 819=>x"6300",
---- 820=>x"6100", 821=>x"6300", 822=>x"6000", 823=>x"5f00", 824=>x"5b00", 825=>x"6100", 826=>x"6000",
---- 827=>x"6100", 828=>x"6200", 829=>x"6200", 830=>x"6000", 831=>x"6300", 832=>x"5c00", 833=>x"6200",
---- 834=>x"6100", 835=>x"5f00", 836=>x"6000", 837=>x"5f00", 838=>x"6000", 839=>x"6300", 840=>x"5e00",
---- 841=>x"5f00", 842=>x"5d00", 843=>x"5f00", 844=>x"6100", 845=>x"6000", 846=>x"6100", 847=>x"6200",
---- 848=>x"5d00", 849=>x"6000", 850=>x"6000", 851=>x"6100", 852=>x"5f00", 853=>x"6000", 854=>x"5f00",
---- 855=>x"5d00", 856=>x"5c00", 857=>x"6200", 858=>x"6400", 859=>x"6400", 860=>x"6200", 861=>x"9c00",
---- 862=>x"6400", 863=>x"6100", 864=>x"5e00", 865=>x"6000", 866=>x"6100", 867=>x"6200", 868=>x"6300",
---- 869=>x"6300", 870=>x"6400", 871=>x"6200", 872=>x"6100", 873=>x"6200", 874=>x"6200", 875=>x"6300",
---- 876=>x"6400", 877=>x"9a00", 878=>x"6200", 879=>x"6400", 880=>x"5d00", 881=>x"6100", 882=>x"6300",
---- 883=>x"6400", 884=>x"6200", 885=>x"6700", 886=>x"6400", 887=>x"6300", 888=>x"5f00", 889=>x"6000",
---- 890=>x"9d00", 891=>x"6300", 892=>x"6400", 893=>x"6400", 894=>x"6700", 895=>x"6500", 896=>x"5e00",
---- 897=>x"6300", 898=>x"6300", 899=>x"6300", 900=>x"6200", 901=>x"6500", 902=>x"6500", 903=>x"6500",
---- 904=>x"5f00", 905=>x"6200", 906=>x"6700", 907=>x"6500", 908=>x"6700", 909=>x"6900", 910=>x"6700",
---- 911=>x"6700", 912=>x"6100", 913=>x"6400", 914=>x"6600", 915=>x"6600", 916=>x"6800", 917=>x"6900",
---- 918=>x"6800", 919=>x"6800", 920=>x"6600", 921=>x"6600", 922=>x"6500", 923=>x"6600", 924=>x"6900",
---- 925=>x"6900", 926=>x"6600", 927=>x"6400", 928=>x"6100", 929=>x"6300", 930=>x"6400", 931=>x"6500",
---- 932=>x"6500", 933=>x"6400", 934=>x"6500", 935=>x"6700", 936=>x"6100", 937=>x"6300", 938=>x"6400",
---- 939=>x"6500", 940=>x"6500", 941=>x"6600", 942=>x"6800", 943=>x"6900", 944=>x"6200", 945=>x"6500",
---- 946=>x"6500", 947=>x"6600", 948=>x"6600", 949=>x"6600", 950=>x"6900", 951=>x"6900", 952=>x"9d00",
---- 953=>x"6200", 954=>x"6600", 955=>x"6500", 956=>x"6800", 957=>x"6700", 958=>x"6900", 959=>x"6a00",
---- 960=>x"6400", 961=>x"6400", 962=>x"6800", 963=>x"6400", 964=>x"6500", 965=>x"6800", 966=>x"6800",
---- 967=>x"6800", 968=>x"6400", 969=>x"6500", 970=>x"6400", 971=>x"6400", 972=>x"9800", 973=>x"6900",
---- 974=>x"6700", 975=>x"6600", 976=>x"6300", 977=>x"6400", 978=>x"6700", 979=>x"6800", 980=>x"6600",
---- 981=>x"6600", 982=>x"6400", 983=>x"6500", 984=>x"6100", 985=>x"6500", 986=>x"6700", 987=>x"6700",
---- 988=>x"6700", 989=>x"6600", 990=>x"6400", 991=>x"6600", 992=>x"6000", 993=>x"6400", 994=>x"6600",
---- 995=>x"6700", 996=>x"6600", 997=>x"6600", 998=>x"9600", 999=>x"6800", 1000=>x"5f00", 1001=>x"9c00",
---- 1002=>x"6a00", 1003=>x"6700", 1004=>x"6600", 1005=>x"6400", 1006=>x"6400", 1007=>x"6300", 1008=>x"6200",
---- 1009=>x"6500", 1010=>x"9600", 1011=>x"6600", 1012=>x"6600", 1013=>x"6500", 1014=>x"6400", 1015=>x"6300",
---- 1016=>x"6400", 1017=>x"6a00", 1018=>x"6700", 1019=>x"6300", 1020=>x"6600", 1021=>x"6400", 1022=>x"6700",
---- 1023=>x"6400", 1024=>x"6200", 1025=>x"9c00", 1026=>x"6500", 1027=>x"6500", 1028=>x"6600", 1029=>x"6300",
---- 1030=>x"6200", 1031=>x"6400", 1032=>x"6200", 1033=>x"6600", 1034=>x"6500", 1035=>x"6800", 1036=>x"6500",
---- 1037=>x"6500", 1038=>x"6400", 1039=>x"6400", 1040=>x"6000", 1041=>x"6100", 1042=>x"6800", 1043=>x"6600",
---- 1044=>x"6300", 1045=>x"6300", 1046=>x"6200", 1047=>x"6200", 1048=>x"5e00", 1049=>x"5e00", 1050=>x"6200",
---- 1051=>x"6400", 1052=>x"6000", 1053=>x"5e00", 1054=>x"6200", 1055=>x"5e00", 1056=>x"6100", 1057=>x"6200",
---- 1058=>x"9f00", 1059=>x"6100", 1060=>x"6100", 1061=>x"6300", 1062=>x"6200", 1063=>x"6000", 1064=>x"6100",
---- 1065=>x"6300", 1066=>x"6400", 1067=>x"6000", 1068=>x"6100", 1069=>x"6200", 1070=>x"6400", 1071=>x"6500",
---- 1072=>x"6500", 1073=>x"6500", 1074=>x"6500", 1075=>x"6600", 1076=>x"6700", 1077=>x"6600", 1078=>x"6700",
---- 1079=>x"6200", 1080=>x"6700", 1081=>x"6a00", 1082=>x"6600", 1083=>x"6600", 1084=>x"6a00", 1085=>x"6600",
---- 1086=>x"6800", 1087=>x"6a00", 1088=>x"6600", 1089=>x"9400", 1090=>x"6b00", 1091=>x"6800", 1092=>x"6900",
---- 1093=>x"6600", 1094=>x"6900", 1095=>x"6300", 1096=>x"6b00", 1097=>x"6e00", 1098=>x"6a00", 1099=>x"6d00",
---- 1100=>x"9200", 1101=>x"7900", 1102=>x"4b00", 1103=>x"3100", 1104=>x"6d00", 1105=>x"6f00", 1106=>x"6f00",
---- 1107=>x"6c00", 1108=>x"7600", 1109=>x"8900", 1110=>x"2900", 1111=>x"2600", 1112=>x"6e00", 1113=>x"6f00",
---- 1114=>x"6f00", 1115=>x"9300", 1116=>x"7600", 1117=>x"8900", 1118=>x"3000", 1119=>x"3000", 1120=>x"6b00",
---- 1121=>x"7000", 1122=>x"7000", 1123=>x"6c00", 1124=>x"6b00", 1125=>x"8a00", 1126=>x"6d00", 1127=>x"7000",
---- 1128=>x"6b00", 1129=>x"6d00", 1130=>x"6b00", 1131=>x"6b00", 1132=>x"6600", 1133=>x"8000", 1134=>x"9f00",
---- 1135=>x"9200", 1136=>x"6a00", 1137=>x"6e00", 1138=>x"6c00", 1139=>x"6c00", 1140=>x"6b00", 1141=>x"6e00",
---- 1142=>x"8a00", 1143=>x"9e00", 1144=>x"6c00", 1145=>x"6f00", 1146=>x"6d00", 1147=>x"6e00", 1148=>x"6c00",
---- 1149=>x"7400", 1150=>x"7700", 1151=>x"8900", 1152=>x"6b00", 1153=>x"6f00", 1154=>x"6d00", 1155=>x"6e00",
---- 1156=>x"6e00", 1157=>x"7500", 1158=>x"7500", 1159=>x"6500", 1160=>x"6800", 1161=>x"6900", 1162=>x"6d00",
---- 1163=>x"7500", 1164=>x"7e00", 1165=>x"8a00", 1166=>x"8600", 1167=>x"8b00", 1168=>x"6800", 1169=>x"7900",
---- 1170=>x"9200", 1171=>x"9800", 1172=>x"9b00", 1173=>x"9700", 1174=>x"9200", 1175=>x"9c00", 1176=>x"8400",
---- 1177=>x"8600", 1178=>x"8400", 1179=>x"7b00", 1180=>x"8300", 1181=>x"7d00", 1182=>x"7e00", 1183=>x"7600",
---- 1184=>x"7100", 1185=>x"6e00", 1186=>x"6d00", 1187=>x"7300", 1188=>x"8300", 1189=>x"7800", 1190=>x"6b00",
---- 1191=>x"6200", 1192=>x"6800", 1193=>x"6d00", 1194=>x"7000", 1195=>x"7500", 1196=>x"8200", 1197=>x"6d00",
---- 1198=>x"5500", 1199=>x"4c00", 1200=>x"6b00", 1201=>x"6c00", 1202=>x"7000", 1203=>x"7200", 1204=>x"7900",
---- 1205=>x"5b00", 1206=>x"4300", 1207=>x"6e00", 1208=>x"6800", 1209=>x"9400", 1210=>x"6e00", 1211=>x"6f00",
---- 1212=>x"6e00", 1213=>x"5900", 1214=>x"7c00", 1215=>x"9700", 1216=>x"6700", 1217=>x"6700", 1218=>x"6c00",
---- 1219=>x"7f00", 1220=>x"8d00", 1221=>x"9100", 1222=>x"8300", 1223=>x"5d00", 1224=>x"6600", 1225=>x"7d00",
---- 1226=>x"9d00", 1227=>x"9c00", 1228=>x"9500", 1229=>x"7200", 1230=>x"2e00", 1231=>x"2e00", 1232=>x"9000",
---- 1233=>x"a100", 1234=>x"8500", 1235=>x"7800", 1236=>x"8300", 1237=>x"5500", 1238=>x"2c00", 1239=>x"3c00",
---- 1240=>x"8900", 1241=>x"7000", 1242=>x"6800", 1243=>x"7c00", 1244=>x"7d00", 1245=>x"5800", 1246=>x"3800",
---- 1247=>x"5500", 1248=>x"8c00", 1249=>x"7500", 1250=>x"7700", 1251=>x"7d00", 1252=>x"8200", 1253=>x"6500",
---- 1254=>x"3400", 1255=>x"4300", 1256=>x"7a00", 1257=>x"7000", 1258=>x"8100", 1259=>x"8600", 1260=>x"8100",
---- 1261=>x"5400", 1262=>x"3a00", 1263=>x"5200", 1264=>x"6f00", 1265=>x"6800", 1266=>x"6f00", 1267=>x"7800",
---- 1268=>x"6900", 1269=>x"4000", 1270=>x"4a00", 1271=>x"5e00", 1272=>x"6800", 1273=>x"6d00", 1274=>x"7400",
---- 1275=>x"7500", 1276=>x"5f00", 1277=>x"4900", 1278=>x"4200", 1279=>x"5300", 1280=>x"6800", 1281=>x"7100",
---- 1282=>x"7900", 1283=>x"7600", 1284=>x"5a00", 1285=>x"4600", 1286=>x"3b00", 1287=>x"aa00", 1288=>x"6500",
---- 1289=>x"6d00", 1290=>x"7a00", 1291=>x"7600", 1292=>x"5700", 1293=>x"4a00", 1294=>x"3f00", 1295=>x"5b00",
---- 1296=>x"6800", 1297=>x"6d00", 1298=>x"7100", 1299=>x"6500", 1300=>x"4a00", 1301=>x"5700", 1302=>x"4a00",
---- 1303=>x"5c00", 1304=>x"6900", 1305=>x"6d00", 1306=>x"7500", 1307=>x"6600", 1308=>x"5400", 1309=>x"5e00",
---- 1310=>x"4800", 1311=>x"5d00", 1312=>x"6900", 1313=>x"7700", 1314=>x"7900", 1315=>x"6600", 1316=>x"5600",
---- 1317=>x"4000", 1318=>x"4300", 1319=>x"5e00", 1320=>x"6b00", 1321=>x"7600", 1322=>x"7400", 1323=>x"7000",
---- 1324=>x"4500", 1325=>x"2500", 1326=>x"3700", 1327=>x"5c00", 1328=>x"6700", 1329=>x"6b00", 1330=>x"7b00",
---- 1331=>x"9300", 1332=>x"5500", 1333=>x"2400", 1334=>x"3400", 1335=>x"5600", 1336=>x"6800", 1337=>x"7600",
---- 1338=>x"9500", 1339=>x"8e00", 1340=>x"5400", 1341=>x"2f00", 1342=>x"3a00", 1343=>x"5a00", 1344=>x"6b00",
---- 1345=>x"9300", 1346=>x"8b00", 1347=>x"6d00", 1348=>x"5300", 1349=>x"3900", 1350=>x"3f00", 1351=>x"4e00",
---- 1352=>x"8b00", 1353=>x"8a00", 1354=>x"6e00", 1355=>x"7700", 1356=>x"4c00", 1357=>x"3d00", 1358=>x"4300",
---- 1359=>x"4c00", 1360=>x"8e00", 1361=>x"6b00", 1362=>x"7600", 1363=>x"7800", 1364=>x"4300", 1365=>x"3b00",
---- 1366=>x"4a00", 1367=>x"6800", 1368=>x"6d00", 1369=>x"6600", 1370=>x"7f00", 1371=>x"7500", 1372=>x"3d00",
---- 1373=>x"b700", 1374=>x"5d00", 1375=>x"6400", 1376=>x"6200", 1377=>x"6800", 1378=>x"7b00", 1379=>x"6700",
---- 1380=>x"4100", 1381=>x"5100", 1382=>x"3600", 1383=>x"5800", 1384=>x"6000", 1385=>x"6600", 1386=>x"8000",
---- 1387=>x"6900", 1388=>x"3f00", 1389=>x"3400", 1390=>x"2900", 1391=>x"6800", 1392=>x"6200", 1393=>x"7400",
---- 1394=>x"9000", 1395=>x"6500", 1396=>x"cb00", 1397=>x"2800", 1398=>x"3f00", 1399=>x"4f00", 1400=>x"7100",
---- 1401=>x"9300", 1402=>x"9600", 1403=>x"5d00", 1404=>x"3600", 1405=>x"3600", 1406=>x"5800", 1407=>x"3400",
---- 1408=>x"7600", 1409=>x"9700", 1410=>x"8300", 1411=>x"5700", 1412=>x"3200", 1413=>x"4a00", 1414=>x"4500",
---- 1415=>x"3300", 1416=>x"9200", 1417=>x"7f00", 1418=>x"7500", 1419=>x"5700", 1420=>x"3e00", 1421=>x"4500",
---- 1422=>x"3d00", 1423=>x"3800", 1424=>x"8700", 1425=>x"6e00", 1426=>x"7100", 1427=>x"5d00", 1428=>x"4300",
---- 1429=>x"3a00", 1430=>x"5700", 1431=>x"4c00", 1432=>x"7400", 1433=>x"6700", 1434=>x"6900", 1435=>x"5200",
---- 1436=>x"4600", 1437=>x"3f00", 1438=>x"7c00", 1439=>x"5900", 1440=>x"6600", 1441=>x"6e00", 1442=>x"6400",
---- 1443=>x"3c00", 1444=>x"4000", 1445=>x"5700", 1446=>x"8800", 1447=>x"4700", 1448=>x"6300", 1449=>x"7600",
---- 1450=>x"6300", 1451=>x"3a00", 1452=>x"2e00", 1453=>x"6600", 1454=>x"8a00", 1455=>x"3300", 1456=>x"6a00",
---- 1457=>x"7600", 1458=>x"4d00", 1459=>x"3500", 1460=>x"3600", 1461=>x"7a00", 1462=>x"8700", 1463=>x"2a00",
---- 1464=>x"7100", 1465=>x"5f00", 1466=>x"3500", 1467=>x"3200", 1468=>x"4000", 1469=>x"7c00", 1470=>x"7500",
---- 1471=>x"2c00", 1472=>x"6200", 1473=>x"4d00", 1474=>x"4000", 1475=>x"3300", 1476=>x"4300", 1477=>x"7800",
---- 1478=>x"5100", 1479=>x"3000", 1480=>x"5d00", 1481=>x"5700", 1482=>x"4200", 1483=>x"4700", 1484=>x"4a00",
---- 1485=>x"5b00", 1486=>x"3c00", 1487=>x"3400", 1488=>x"5b00", 1489=>x"4b00", 1490=>x"4300", 1491=>x"5d00",
---- 1492=>x"5b00", 1493=>x"5200", 1494=>x"3900", 1495=>x"3200", 1496=>x"5d00", 1497=>x"4600", 1498=>x"4b00",
---- 1499=>x"5900", 1500=>x"5e00", 1501=>x"5400", 1502=>x"3800", 1503=>x"3400", 1504=>x"5600", 1505=>x"3c00",
---- 1506=>x"4b00", 1507=>x"3900", 1508=>x"6200", 1509=>x"5900", 1510=>x"3200", 1511=>x"3c00", 1512=>x"4100",
---- 1513=>x"3c00", 1514=>x"4100", 1515=>x"3200", 1516=>x"7400", 1517=>x"5700", 1518=>x"2d00", 1519=>x"3d00",
---- 1520=>x"3000", 1521=>x"3900", 1522=>x"3300", 1523=>x"3500", 1524=>x"7500", 1525=>x"5d00", 1526=>x"3000",
---- 1527=>x"3900", 1528=>x"3000", 1529=>x"3100", 1530=>x"3900", 1531=>x"4500", 1532=>x"6400", 1533=>x"5600",
---- 1534=>x"3500", 1535=>x"3800", 1536=>x"3e00", 1537=>x"2800", 1538=>x"3f00", 1539=>x"5f00", 1540=>x"4f00",
---- 1541=>x"4600", 1542=>x"3e00", 1543=>x"3900", 1544=>x"4100", 1545=>x"2500", 1546=>x"3500", 1547=>x"5300",
---- 1548=>x"4c00", 1549=>x"3a00", 1550=>x"4000", 1551=>x"3c00", 1552=>x"3700", 1553=>x"2600", 1554=>x"2b00",
---- 1555=>x"4d00", 1556=>x"5600", 1557=>x"3500", 1558=>x"3a00", 1559=>x"4300", 1560=>x"3600", 1561=>x"3400",
---- 1562=>x"2800", 1563=>x"4700", 1564=>x"5900", 1565=>x"4200", 1566=>x"3e00", 1567=>x"4000", 1568=>x"2900",
---- 1569=>x"2b00", 1570=>x"2600", 1571=>x"4400", 1572=>x"6000", 1573=>x"4800", 1574=>x"3a00", 1575=>x"3f00",
---- 1576=>x"2400", 1577=>x"2a00", 1578=>x"2400", 1579=>x"3d00", 1580=>x"6000", 1581=>x"4c00", 1582=>x"3b00",
---- 1583=>x"3b00", 1584=>x"2600", 1585=>x"2a00", 1586=>x"2400", 1587=>x"3000", 1588=>x"5600", 1589=>x"4f00",
---- 1590=>x"2c00", 1591=>x"3700", 1592=>x"2900", 1593=>x"2b00", 1594=>x"2700", 1595=>x"2900", 1596=>x"3a00",
---- 1597=>x"5400", 1598=>x"3f00", 1599=>x"4400", 1600=>x"2800", 1601=>x"2700", 1602=>x"2600", 1603=>x"2d00",
---- 1604=>x"2b00", 1605=>x"4000", 1606=>x"6100", 1607=>x"6600", 1608=>x"2a00", 1609=>x"2b00", 1610=>x"2b00",
---- 1611=>x"2c00", 1612=>x"2a00", 1613=>x"3100", 1614=>x"5c00", 1615=>x"7400", 1616=>x"2a00", 1617=>x"2a00",
---- 1618=>x"2a00", 1619=>x"2500", 1620=>x"4200", 1621=>x"6500", 1622=>x"6400", 1623=>x"6700", 1624=>x"2a00",
---- 1625=>x"2400", 1626=>x"2600", 1627=>x"de00", 1628=>x"d100", 1629=>x"6500", 1630=>x"8100", 1631=>x"8100",
---- 1632=>x"2a00", 1633=>x"2500", 1634=>x"2b00", 1635=>x"2600", 1636=>x"2700", 1637=>x"3a00", 1638=>x"4800",
---- 1639=>x"4e00", 1640=>x"2f00", 1641=>x"2f00", 1642=>x"2b00", 1643=>x"2b00", 1644=>x"3600", 1645=>x"4b00",
---- 1646=>x"3700", 1647=>x"1e00", 1648=>x"3900", 1649=>x"3c00", 1650=>x"3900", 1651=>x"3a00", 1652=>x"4300",
---- 1653=>x"4b00", 1654=>x"4100", 1655=>x"2a00", 1656=>x"3200", 1657=>x"ca00", 1658=>x"3100", 1659=>x"3500",
---- 1660=>x"4400", 1661=>x"4300", 1662=>x"4400", 1663=>x"3500", 1664=>x"2a00", 1665=>x"3100", 1666=>x"2c00",
---- 1667=>x"2d00", 1668=>x"4700", 1669=>x"3700", 1670=>x"3a00", 1671=>x"3e00", 1672=>x"2700", 1673=>x"3100",
---- 1674=>x"2a00", 1675=>x"3f00", 1676=>x"5000", 1677=>x"2d00", 1678=>x"3700", 1679=>x"3600", 1680=>x"2b00",
---- 1681=>x"3300", 1682=>x"2a00", 1683=>x"5700", 1684=>x"4300", 1685=>x"2c00", 1686=>x"3000", 1687=>x"3600",
---- 1688=>x"2d00", 1689=>x"2e00", 1690=>x"3b00", 1691=>x"5300", 1692=>x"3200", 1693=>x"2900", 1694=>x"3000",
---- 1695=>x"3500", 1696=>x"3200", 1697=>x"3600", 1698=>x"4400", 1699=>x"3800", 1700=>x"2c00", 1701=>x"2d00",
---- 1702=>x"3100", 1703=>x"3200", 1704=>x"2f00", 1705=>x"3b00", 1706=>x"3a00", 1707=>x"3500", 1708=>x"2e00",
---- 1709=>x"2e00", 1710=>x"3000", 1711=>x"3100", 1712=>x"3500", 1713=>x"3b00", 1714=>x"3200", 1715=>x"3500",
---- 1716=>x"3300", 1717=>x"d100", 1718=>x"3000", 1719=>x"3200", 1720=>x"4000", 1721=>x"3400", 1722=>x"2e00",
---- 1723=>x"3400", 1724=>x"2c00", 1725=>x"2900", 1726=>x"3100", 1727=>x"3400", 1728=>x"3b00", 1729=>x"cf00",
---- 1730=>x"2c00", 1731=>x"3200", 1732=>x"2d00", 1733=>x"2900", 1734=>x"3500", 1735=>x"2d00", 1736=>x"3000",
---- 1737=>x"2c00", 1738=>x"2a00", 1739=>x"2d00", 1740=>x"2a00", 1741=>x"2c00", 1742=>x"3300", 1743=>x"2500",
---- 1744=>x"2d00", 1745=>x"2c00", 1746=>x"2a00", 1747=>x"2e00", 1748=>x"2d00", 1749=>x"3100", 1750=>x"2900",
---- 1751=>x"2500", 1752=>x"2c00", 1753=>x"3000", 1754=>x"2d00", 1755=>x"2d00", 1756=>x"2d00", 1757=>x"2f00",
---- 1758=>x"2800", 1759=>x"2800", 1760=>x"3000", 1761=>x"2e00", 1762=>x"2c00", 1763=>x"2f00", 1764=>x"2e00",
---- 1765=>x"2d00", 1766=>x"3600", 1767=>x"4200", 1768=>x"2e00", 1769=>x"2c00", 1770=>x"3200", 1771=>x"3100",
---- 1772=>x"2e00", 1773=>x"3b00", 1774=>x"5d00", 1775=>x"4400", 1776=>x"2b00", 1777=>x"2b00", 1778=>x"3200",
---- 1779=>x"3600", 1780=>x"2c00", 1781=>x"3d00", 1782=>x"4c00", 1783=>x"2c00", 1784=>x"2f00", 1785=>x"2e00",
---- 1786=>x"3300", 1787=>x"3100", 1788=>x"2b00", 1789=>x"3100", 1790=>x"2f00", 1791=>x"3300", 1792=>x"2e00",
---- 1793=>x"2c00", 1794=>x"3100", 1795=>x"3100", 1796=>x"2f00", 1797=>x"3200", 1798=>x"2f00", 1799=>x"c200",
---- 1800=>x"2b00", 1801=>x"2a00", 1802=>x"3400", 1803=>x"2f00", 1804=>x"2c00", 1805=>x"3100", 1806=>x"4400",
---- 1807=>x"4400", 1808=>x"2600", 1809=>x"2d00", 1810=>x"3700", 1811=>x"2800", 1812=>x"3c00", 1813=>x"5400",
---- 1814=>x"4800", 1815=>x"3b00", 1816=>x"2700", 1817=>x"2d00", 1818=>x"3600", 1819=>x"4900", 1820=>x"5b00",
---- 1821=>x"4c00", 1822=>x"3200", 1823=>x"2e00", 1824=>x"2c00", 1825=>x"4600", 1826=>x"5400", 1827=>x"5000",
---- 1828=>x"3c00", 1829=>x"2b00", 1830=>x"2d00", 1831=>x"2c00", 1832=>x"3300", 1833=>x"4000", 1834=>x"3b00",
---- 1835=>x"3100", 1836=>x"3200", 1837=>x"3100", 1838=>x"2f00", 1839=>x"3200", 1840=>x"2d00", 1841=>x"2f00",
---- 1842=>x"2e00", 1843=>x"3300", 1844=>x"3000", 1845=>x"2c00", 1846=>x"2e00", 1847=>x"3700", 1848=>x"3000",
---- 1849=>x"3600", 1850=>x"3600", 1851=>x"3200", 1852=>x"3100", 1853=>x"2d00", 1854=>x"2d00", 1855=>x"3100",
---- 1856=>x"3a00", 1857=>x"3900", 1858=>x"2e00", 1859=>x"2d00", 1860=>x"3100", 1861=>x"2f00", 1862=>x"2f00",
---- 1863=>x"3a00", 1864=>x"3d00", 1865=>x"2d00", 1866=>x"2c00", 1867=>x"2d00", 1868=>x"3000", 1869=>x"2f00",
---- 1870=>x"2e00", 1871=>x"bc00", 1872=>x"2f00", 1873=>x"2a00", 1874=>x"2e00", 1875=>x"2b00", 1876=>x"2c00",
---- 1877=>x"2d00", 1878=>x"3e00", 1879=>x"4600", 1880=>x"2900", 1881=>x"2e00", 1882=>x"2c00", 1883=>x"2700",
---- 1884=>x"2b00", 1885=>x"4300", 1886=>x"4800", 1887=>x"3800", 1888=>x"2700", 1889=>x"2c00", 1890=>x"2b00",
---- 1891=>x"2b00", 1892=>x"3900", 1893=>x"4700", 1894=>x"3500", 1895=>x"3500", 1896=>x"2b00", 1897=>x"2f00",
---- 1898=>x"3600", 1899=>x"3b00", 1900=>x"3200", 1901=>x"2e00", 1902=>x"3100", 1903=>x"3900", 1904=>x"3100",
---- 1905=>x"4100", 1906=>x"4700", 1907=>x"3200", 1908=>x"2c00", 1909=>x"2d00", 1910=>x"2f00", 1911=>x"3a00",
---- 1912=>x"3b00", 1913=>x"3b00", 1914=>x"3500", 1915=>x"2e00", 1916=>x"3200", 1917=>x"2d00", 1918=>x"3100",
---- 1919=>x"3000", 1920=>x"2e00", 1921=>x"2f00", 1922=>x"3100", 1923=>x"2e00", 1924=>x"2e00", 1925=>x"2e00",
---- 1926=>x"3200", 1927=>x"3700", 1928=>x"3000", 1929=>x"2f00", 1930=>x"3100", 1931=>x"2d00", 1932=>x"3000",
---- 1933=>x"2e00", 1934=>x"3100", 1935=>x"3a00", 1936=>x"2f00", 1937=>x"2f00", 1938=>x"2d00", 1939=>x"3200",
---- 1940=>x"3800", 1941=>x"2d00", 1942=>x"3000", 1943=>x"3700", 1944=>x"3300", 1945=>x"3800", 1946=>x"2f00",
---- 1947=>x"3800", 1948=>x"3a00", 1949=>x"2f00", 1950=>x"3300", 1951=>x"3b00", 1952=>x"3300", 1953=>x"3a00",
---- 1954=>x"3000", 1955=>x"3b00", 1956=>x"3c00", 1957=>x"d300", 1958=>x"2f00", 1959=>x"3500", 1960=>x"3500",
---- 1961=>x"3600", 1962=>x"2800", 1963=>x"3f00", 1964=>x"3f00", 1965=>x"2f00", 1966=>x"3000", 1967=>x"2f00",
---- 1968=>x"3300", 1969=>x"3500", 1970=>x"3300", 1971=>x"3e00", 1972=>x"3f00", 1973=>x"3100", 1974=>x"3400",
---- 1975=>x"3000", 1976=>x"2e00", 1977=>x"3100", 1978=>x"3400", 1979=>x"4000", 1980=>x"3a00", 1981=>x"3600",
---- 1982=>x"3700", 1983=>x"3600", 1984=>x"2a00", 1985=>x"2d00", 1986=>x"3800", 1987=>x"4300", 1988=>x"4000",
---- 1989=>x"3c00", 1990=>x"3900", 1991=>x"3500", 1992=>x"2e00", 1993=>x"3300", 1994=>x"3600", 1995=>x"3f00",
---- 1996=>x"c800", 1997=>x"3900", 1998=>x"3900", 1999=>x"3c00", 2000=>x"2f00", 2001=>x"3400", 2002=>x"3900",
---- 2003=>x"3f00", 2004=>x"3500", 2005=>x"3600", 2006=>x"3a00", 2007=>x"4200", 2008=>x"2e00", 2009=>x"3400",
---- 2010=>x"3800", 2011=>x"3c00", 2012=>x"3600", 2013=>x"3900", 2014=>x"3d00", 2015=>x"4300", 2016=>x"3500",
---- 2017=>x"3e00", 2018=>x"3d00", 2019=>x"3700", 2020=>x"3800", 2021=>x"3b00", 2022=>x"4000", 2023=>x"4200",
---- 2024=>x"3800", 2025=>x"3600", 2026=>x"3c00", 2027=>x"3900", 2028=>x"3d00", 2029=>x"3f00", 2030=>x"5000",
---- 2031=>x"4c00", 2032=>x"3900", 2033=>x"3d00", 2034=>x"3c00", 2035=>x"3e00", 2036=>x"3d00", 2037=>x"4300",
---- 2038=>x"4b00", 2039=>x"4d00", 2040=>x"3800", 2041=>x"3700", 2042=>x"3c00", 2043=>x"4700", 2044=>x"4000",
---- 2045=>x"4200", 2046=>x"4300", 2047=>x"4100"),
---- 6  => (0=>x"6d00", 1=>x"6d00", 2=>x"6800", 3=>x"6a00", 4=>x"9200", 5=>x"7000", 6=>x"7100", 7=>x"7800",
---- 8=>x"6f00", 9=>x"6d00", 10=>x"6900", 11=>x"6a00", 12=>x"6e00", 13=>x"7200", 14=>x"7100",
---- 15=>x"7800", 16=>x"6c00", 17=>x"6c00", 18=>x"6900", 19=>x"6800", 20=>x"6d00", 21=>x"7200",
---- 22=>x"7200", 23=>x"7700", 24=>x"6a00", 25=>x"6a00", 26=>x"6800", 27=>x"6b00", 28=>x"6b00",
---- 29=>x"6e00", 30=>x"7400", 31=>x"7500", 32=>x"6700", 33=>x"6a00", 34=>x"6800", 35=>x"6b00",
---- 36=>x"6e00", 37=>x"6e00", 38=>x"7000", 39=>x"7400", 40=>x"6800", 41=>x"6600", 42=>x"6700",
---- 43=>x"6c00", 44=>x"6e00", 45=>x"6d00", 46=>x"7200", 47=>x"7400", 48=>x"6700", 49=>x"6700",
---- 50=>x"6500", 51=>x"6700", 52=>x"7000", 53=>x"8f00", 54=>x"7100", 55=>x"7400", 56=>x"6900",
---- 57=>x"6500", 58=>x"6600", 59=>x"6800", 60=>x"6e00", 61=>x"6e00", 62=>x"7000", 63=>x"7400",
---- 64=>x"6700", 65=>x"6800", 66=>x"6500", 67=>x"6700", 68=>x"6b00", 69=>x"6f00", 70=>x"7000",
---- 71=>x"7400", 72=>x"6500", 73=>x"6700", 74=>x"6600", 75=>x"6900", 76=>x"9200", 77=>x"7100",
---- 78=>x"7300", 79=>x"7500", 80=>x"6900", 81=>x"6800", 82=>x"6600", 83=>x"6500", 84=>x"6e00",
---- 85=>x"7100", 86=>x"7300", 87=>x"7100", 88=>x"6600", 89=>x"6700", 90=>x"6700", 91=>x"6900",
---- 92=>x"6d00", 93=>x"6f00", 94=>x"6f00", 95=>x"7300", 96=>x"6600", 97=>x"6600", 98=>x"6800",
---- 99=>x"6b00", 100=>x"6b00", 101=>x"6e00", 102=>x"6f00", 103=>x"6f00", 104=>x"6800", 105=>x"6600",
---- 106=>x"6700", 107=>x"6c00", 108=>x"6e00", 109=>x"6d00", 110=>x"6f00", 111=>x"7200", 112=>x"6700",
---- 113=>x"6500", 114=>x"6800", 115=>x"6b00", 116=>x"6b00", 117=>x"6c00", 118=>x"7100", 119=>x"7300",
---- 120=>x"6900", 121=>x"6600", 122=>x"6600", 123=>x"6b00", 124=>x"6c00", 125=>x"6b00", 126=>x"6e00",
---- 127=>x"7300", 128=>x"6700", 129=>x"6500", 130=>x"6800", 131=>x"6a00", 132=>x"6b00", 133=>x"6e00",
---- 134=>x"7100", 135=>x"7100", 136=>x"6400", 137=>x"6500", 138=>x"6600", 139=>x"6800", 140=>x"6b00",
---- 141=>x"6f00", 142=>x"6f00", 143=>x"7200", 144=>x"6600", 145=>x"6800", 146=>x"6800", 147=>x"6900",
---- 148=>x"6b00", 149=>x"6e00", 150=>x"7200", 151=>x"7000", 152=>x"6600", 153=>x"6900", 154=>x"6500",
---- 155=>x"6800", 156=>x"6b00", 157=>x"6e00", 158=>x"7000", 159=>x"7300", 160=>x"6600", 161=>x"6600",
---- 162=>x"6600", 163=>x"6700", 164=>x"6900", 165=>x"6f00", 166=>x"7200", 167=>x"7400", 168=>x"6500",
---- 169=>x"6500", 170=>x"6700", 171=>x"6700", 172=>x"6900", 173=>x"6d00", 174=>x"6f00", 175=>x"7100",
---- 176=>x"6700", 177=>x"6500", 178=>x"6700", 179=>x"6800", 180=>x"6d00", 181=>x"6c00", 182=>x"6f00",
---- 183=>x"7400", 184=>x"6600", 185=>x"6600", 186=>x"6800", 187=>x"6900", 188=>x"7000", 189=>x"6c00",
---- 190=>x"7200", 191=>x"7500", 192=>x"6500", 193=>x"6500", 194=>x"6700", 195=>x"6a00", 196=>x"6f00",
---- 197=>x"7000", 198=>x"7000", 199=>x"6f00", 200=>x"6700", 201=>x"6500", 202=>x"6700", 203=>x"6a00",
---- 204=>x"6e00", 205=>x"7200", 206=>x"7100", 207=>x"7100", 208=>x"6900", 209=>x"6900", 210=>x"6a00",
---- 211=>x"6d00", 212=>x"6c00", 213=>x"6f00", 214=>x"7100", 215=>x"7400", 216=>x"6a00", 217=>x"6700",
---- 218=>x"6800", 219=>x"6b00", 220=>x"6d00", 221=>x"7100", 222=>x"7700", 223=>x"7300", 224=>x"6800",
---- 225=>x"6800", 226=>x"6900", 227=>x"6800", 228=>x"6c00", 229=>x"6f00", 230=>x"7700", 231=>x"7300",
---- 232=>x"6200", 233=>x"6a00", 234=>x"6c00", 235=>x"9600", 236=>x"6a00", 237=>x"6e00", 238=>x"7100",
---- 239=>x"7100", 240=>x"6500", 241=>x"6800", 242=>x"6800", 243=>x"6a00", 244=>x"6b00", 245=>x"6e00",
---- 246=>x"7000", 247=>x"7100", 248=>x"9800", 249=>x"6400", 250=>x"6700", 251=>x"6900", 252=>x"6b00",
---- 253=>x"6e00", 254=>x"6e00", 255=>x"7200", 256=>x"6400", 257=>x"6600", 258=>x"6900", 259=>x"6800",
---- 260=>x"6900", 261=>x"6d00", 262=>x"6c00", 263=>x"6f00", 264=>x"6400", 265=>x"6600", 266=>x"6800",
---- 267=>x"6700", 268=>x"6700", 269=>x"6a00", 270=>x"6600", 271=>x"6d00", 272=>x"6500", 273=>x"6600",
---- 274=>x"6300", 275=>x"6400", 276=>x"6900", 277=>x"6a00", 278=>x"6c00", 279=>x"6f00", 280=>x"6500",
---- 281=>x"6500", 282=>x"6700", 283=>x"6800", 284=>x"6b00", 285=>x"6c00", 286=>x"6c00", 287=>x"6f00",
---- 288=>x"6400", 289=>x"6500", 290=>x"6100", 291=>x"6400", 292=>x"6800", 293=>x"6b00", 294=>x"6d00",
---- 295=>x"6d00", 296=>x"6300", 297=>x"6300", 298=>x"6300", 299=>x"6700", 300=>x"6900", 301=>x"6a00",
---- 302=>x"6d00", 303=>x"6d00", 304=>x"6400", 305=>x"6400", 306=>x"6600", 307=>x"6600", 308=>x"6800",
---- 309=>x"6800", 310=>x"6c00", 311=>x"6e00", 312=>x"6500", 313=>x"6500", 314=>x"6500", 315=>x"6800",
---- 316=>x"6700", 317=>x"6a00", 318=>x"6e00", 319=>x"7000", 320=>x"6700", 321=>x"6600", 322=>x"9b00",
---- 323=>x"6700", 324=>x"6a00", 325=>x"6c00", 326=>x"6d00", 327=>x"6e00", 328=>x"6400", 329=>x"6500",
---- 330=>x"6600", 331=>x"6800", 332=>x"6900", 333=>x"6b00", 334=>x"6e00", 335=>x"6e00", 336=>x"6300",
---- 337=>x"6500", 338=>x"6500", 339=>x"6700", 340=>x"6600", 341=>x"6900", 342=>x"7000", 343=>x"7000",
---- 344=>x"6600", 345=>x"6400", 346=>x"6400", 347=>x"6600", 348=>x"6700", 349=>x"6a00", 350=>x"6b00",
---- 351=>x"6e00", 352=>x"6600", 353=>x"6300", 354=>x"6500", 355=>x"6600", 356=>x"6900", 357=>x"6d00",
---- 358=>x"9200", 359=>x"6c00", 360=>x"6400", 361=>x"6400", 362=>x"6300", 363=>x"6500", 364=>x"6b00",
---- 365=>x"6e00", 366=>x"6c00", 367=>x"6c00", 368=>x"6200", 369=>x"6200", 370=>x"6600", 371=>x"6700",
---- 372=>x"6a00", 373=>x"6600", 374=>x"6b00", 375=>x"6e00", 376=>x"6600", 377=>x"6300", 378=>x"6300",
---- 379=>x"6a00", 380=>x"6900", 381=>x"6700", 382=>x"6b00", 383=>x"6e00", 384=>x"6500", 385=>x"6500",
---- 386=>x"6400", 387=>x"6800", 388=>x"6500", 389=>x"6700", 390=>x"6b00", 391=>x"6f00", 392=>x"6300",
---- 393=>x"6300", 394=>x"6700", 395=>x"6800", 396=>x"9800", 397=>x"6a00", 398=>x"6900", 399=>x"6d00",
---- 400=>x"6300", 401=>x"6600", 402=>x"6800", 403=>x"6600", 404=>x"6700", 405=>x"6a00", 406=>x"6e00",
---- 407=>x"6d00", 408=>x"6500", 409=>x"6800", 410=>x"6400", 411=>x"6600", 412=>x"6600", 413=>x"6a00",
---- 414=>x"6d00", 415=>x"6f00", 416=>x"6400", 417=>x"6600", 418=>x"6200", 419=>x"6500", 420=>x"6700",
---- 421=>x"6900", 422=>x"6d00", 423=>x"6e00", 424=>x"6200", 425=>x"6100", 426=>x"6600", 427=>x"6300",
---- 428=>x"6700", 429=>x"6a00", 430=>x"6b00", 431=>x"6e00", 432=>x"6200", 433=>x"6300", 434=>x"6500",
---- 435=>x"6500", 436=>x"6700", 437=>x"6800", 438=>x"6a00", 439=>x"6e00", 440=>x"9b00", 441=>x"6400",
---- 442=>x"6500", 443=>x"6400", 444=>x"6b00", 445=>x"6c00", 446=>x"6d00", 447=>x"6d00", 448=>x"6600",
---- 449=>x"6400", 450=>x"6700", 451=>x"6b00", 452=>x"6d00", 453=>x"6a00", 454=>x"6e00", 455=>x"6f00",
---- 456=>x"6000", 457=>x"6500", 458=>x"6800", 459=>x"6d00", 460=>x"6c00", 461=>x"6b00", 462=>x"6b00",
---- 463=>x"6c00", 464=>x"6300", 465=>x"6300", 466=>x"6300", 467=>x"6700", 468=>x"6400", 469=>x"6900",
---- 470=>x"6b00", 471=>x"6e00", 472=>x"6100", 473=>x"6100", 474=>x"6300", 475=>x"6a00", 476=>x"6700",
---- 477=>x"6800", 478=>x"6900", 479=>x"6a00", 480=>x"6300", 481=>x"6300", 482=>x"6400", 483=>x"6600",
---- 484=>x"6800", 485=>x"9700", 486=>x"6b00", 487=>x"6b00", 488=>x"6300", 489=>x"6400", 490=>x"6300",
---- 491=>x"6600", 492=>x"6800", 493=>x"6800", 494=>x"6900", 495=>x"6900", 496=>x"6300", 497=>x"6500",
---- 498=>x"6300", 499=>x"6500", 500=>x"6800", 501=>x"6800", 502=>x"6a00", 503=>x"6a00", 504=>x"6500",
---- 505=>x"6400", 506=>x"6400", 507=>x"6700", 508=>x"6500", 509=>x"6900", 510=>x"6d00", 511=>x"6f00",
---- 512=>x"6500", 513=>x"6400", 514=>x"6800", 515=>x"6900", 516=>x"6a00", 517=>x"6900", 518=>x"6d00",
---- 519=>x"6d00", 520=>x"6400", 521=>x"6400", 522=>x"6600", 523=>x"6c00", 524=>x"6900", 525=>x"6a00",
---- 526=>x"6d00", 527=>x"6c00", 528=>x"6700", 529=>x"6500", 530=>x"6600", 531=>x"6900", 532=>x"6c00",
---- 533=>x"6c00", 534=>x"6e00", 535=>x"6e00", 536=>x"6600", 537=>x"6300", 538=>x"6300", 539=>x"6600",
---- 540=>x"6d00", 541=>x"6f00", 542=>x"6d00", 543=>x"6e00", 544=>x"6700", 545=>x"6200", 546=>x"6000",
---- 547=>x"6600", 548=>x"9300", 549=>x"6900", 550=>x"6c00", 551=>x"6e00", 552=>x"6700", 553=>x"6200",
---- 554=>x"6300", 555=>x"6600", 556=>x"6500", 557=>x"6a00", 558=>x"6c00", 559=>x"6c00", 560=>x"6500",
---- 561=>x"6400", 562=>x"6300", 563=>x"6400", 564=>x"6600", 565=>x"6a00", 566=>x"6a00", 567=>x"6c00",
---- 568=>x"6100", 569=>x"6500", 570=>x"6400", 571=>x"6400", 572=>x"6600", 573=>x"6b00", 574=>x"6c00",
---- 575=>x"6c00", 576=>x"6000", 577=>x"6200", 578=>x"6500", 579=>x"6600", 580=>x"6600", 581=>x"6800",
---- 582=>x"6900", 583=>x"6900", 584=>x"6000", 585=>x"6300", 586=>x"6300", 587=>x"6200", 588=>x"6500",
---- 589=>x"6500", 590=>x"6700", 591=>x"6a00", 592=>x"6200", 593=>x"6200", 594=>x"6300", 595=>x"6300",
---- 596=>x"6300", 597=>x"6500", 598=>x"6a00", 599=>x"6900", 600=>x"6300", 601=>x"6000", 602=>x"6200",
---- 603=>x"6500", 604=>x"6400", 605=>x"6600", 606=>x"6d00", 607=>x"6900", 608=>x"6100", 609=>x"6400",
---- 610=>x"6100", 611=>x"6300", 612=>x"6600", 613=>x"6700", 614=>x"6700", 615=>x"6800", 616=>x"6100",
---- 617=>x"6300", 618=>x"6200", 619=>x"6200", 620=>x"6500", 621=>x"6800", 622=>x"6600", 623=>x"6a00",
---- 624=>x"6200", 625=>x"6200", 626=>x"6200", 627=>x"6400", 628=>x"6300", 629=>x"6600", 630=>x"6500",
---- 631=>x"6700", 632=>x"6200", 633=>x"6200", 634=>x"6200", 635=>x"6600", 636=>x"6300", 637=>x"6500",
---- 638=>x"6800", 639=>x"6600", 640=>x"6400", 641=>x"6100", 642=>x"6100", 643=>x"6300", 644=>x"6500",
---- 645=>x"6500", 646=>x"6700", 647=>x"6600", 648=>x"6200", 649=>x"6200", 650=>x"6100", 651=>x"6300",
---- 652=>x"6600", 653=>x"9b00", 654=>x"6400", 655=>x"6200", 656=>x"6200", 657=>x"6200", 658=>x"6800",
---- 659=>x"6600", 660=>x"6400", 661=>x"6400", 662=>x"6400", 663=>x"6200", 664=>x"6100", 665=>x"6000",
---- 666=>x"6300", 667=>x"6200", 668=>x"6200", 669=>x"6100", 670=>x"6400", 671=>x"6500", 672=>x"6200",
---- 673=>x"9e00", 674=>x"6200", 675=>x"6100", 676=>x"6200", 677=>x"6200", 678=>x"6500", 679=>x"6200",
---- 680=>x"6300", 681=>x"6200", 682=>x"6400", 683=>x"6200", 684=>x"6000", 685=>x"6200", 686=>x"6200",
---- 687=>x"5e00", 688=>x"6000", 689=>x"6100", 690=>x"6200", 691=>x"6200", 692=>x"6600", 693=>x"6400",
---- 694=>x"6400", 695=>x"6000", 696=>x"9d00", 697=>x"6300", 698=>x"6000", 699=>x"9d00", 700=>x"6200",
---- 701=>x"6300", 702=>x"5f00", 703=>x"5f00", 704=>x"6300", 705=>x"6400", 706=>x"6200", 707=>x"6300",
---- 708=>x"6500", 709=>x"6200", 710=>x"6100", 711=>x"5f00", 712=>x"6300", 713=>x"6400", 714=>x"6400",
---- 715=>x"6100", 716=>x"6400", 717=>x"6300", 718=>x"6300", 719=>x"5e00", 720=>x"6200", 721=>x"5f00",
---- 722=>x"6200", 723=>x"6200", 724=>x"6400", 725=>x"6400", 726=>x"6100", 727=>x"5f00", 728=>x"6200",
---- 729=>x"6300", 730=>x"6400", 731=>x"6300", 732=>x"6400", 733=>x"6500", 734=>x"6600", 735=>x"6100",
---- 736=>x"6400", 737=>x"6100", 738=>x"6400", 739=>x"6400", 740=>x"6500", 741=>x"6200", 742=>x"6200",
---- 743=>x"6000", 744=>x"6500", 745=>x"6100", 746=>x"6500", 747=>x"6400", 748=>x"6300", 749=>x"6100",
---- 750=>x"6200", 751=>x"6000", 752=>x"6500", 753=>x"5d00", 754=>x"6100", 755=>x"6500", 756=>x"6300",
---- 757=>x"6100", 758=>x"5f00", 759=>x"a200", 760=>x"6500", 761=>x"6100", 762=>x"6000", 763=>x"6400",
---- 764=>x"6400", 765=>x"6000", 766=>x"6000", 767=>x"6200", 768=>x"6300", 769=>x"6100", 770=>x"6300",
---- 771=>x"6200", 772=>x"6700", 773=>x"6400", 774=>x"6400", 775=>x"6300", 776=>x"6200", 777=>x"6300",
---- 778=>x"6300", 779=>x"6100", 780=>x"6100", 781=>x"6200", 782=>x"6400", 783=>x"6500", 784=>x"6500",
---- 785=>x"6300", 786=>x"6200", 787=>x"6200", 788=>x"6100", 789=>x"6000", 790=>x"6000", 791=>x"6500",
---- 792=>x"6000", 793=>x"6000", 794=>x"6000", 795=>x"6400", 796=>x"6200", 797=>x"6100", 798=>x"9a00",
---- 799=>x"6600", 800=>x"5f00", 801=>x"5d00", 802=>x"5f00", 803=>x"6100", 804=>x"6000", 805=>x"5f00",
---- 806=>x"6600", 807=>x"6800", 808=>x"6100", 809=>x"6400", 810=>x"6000", 811=>x"6200", 812=>x"6200",
---- 813=>x"6100", 814=>x"6600", 815=>x"6800", 816=>x"6000", 817=>x"6300", 818=>x"5f00", 819=>x"6100",
---- 820=>x"6300", 821=>x"6000", 822=>x"6700", 823=>x"6800", 824=>x"9b00", 825=>x"6200", 826=>x"a100",
---- 827=>x"6000", 828=>x"6300", 829=>x"6500", 830=>x"6800", 831=>x"6900", 832=>x"6100", 833=>x"6300",
---- 834=>x"6500", 835=>x"6500", 836=>x"6400", 837=>x"6600", 838=>x"6800", 839=>x"6700", 840=>x"6200",
---- 841=>x"6000", 842=>x"6400", 843=>x"6200", 844=>x"6100", 845=>x"6700", 846=>x"6b00", 847=>x"6800",
---- 848=>x"6000", 849=>x"6300", 850=>x"6200", 851=>x"6300", 852=>x"6400", 853=>x"6400", 854=>x"6700",
---- 855=>x"6c00", 856=>x"6000", 857=>x"6100", 858=>x"6100", 859=>x"6100", 860=>x"6600", 861=>x"6400",
---- 862=>x"6900", 863=>x"6700", 864=>x"6300", 865=>x"6300", 866=>x"6000", 867=>x"6000", 868=>x"6300",
---- 869=>x"6400", 870=>x"6900", 871=>x"6800", 872=>x"6300", 873=>x"6300", 874=>x"6300", 875=>x"6300",
---- 876=>x"6200", 877=>x"6700", 878=>x"6900", 879=>x"6a00", 880=>x"6200", 881=>x"6200", 882=>x"6300",
---- 883=>x"6500", 884=>x"6400", 885=>x"6900", 886=>x"6b00", 887=>x"6a00", 888=>x"6100", 889=>x"6300",
---- 890=>x"6300", 891=>x"6500", 892=>x"6800", 893=>x"6700", 894=>x"6800", 895=>x"6e00", 896=>x"6500",
---- 897=>x"6600", 898=>x"6500", 899=>x"6500", 900=>x"6600", 901=>x"6800", 902=>x"6400", 903=>x"9b00",
---- 904=>x"6400", 905=>x"6400", 906=>x"6300", 907=>x"6400", 908=>x"6300", 909=>x"6400", 910=>x"6300",
---- 911=>x"7700", 912=>x"6500", 913=>x"6100", 914=>x"6300", 915=>x"6300", 916=>x"6300", 917=>x"6300",
---- 918=>x"6d00", 919=>x"9600", 920=>x"6400", 921=>x"6300", 922=>x"6300", 923=>x"6400", 924=>x"6800",
---- 925=>x"6700", 926=>x"7200", 927=>x"7700", 928=>x"6300", 929=>x"6800", 930=>x"6500", 931=>x"6700",
---- 932=>x"6800", 933=>x"6800", 934=>x"6d00", 935=>x"7800", 936=>x"6600", 937=>x"6700", 938=>x"6600",
---- 939=>x"6600", 940=>x"6500", 941=>x"6700", 942=>x"6a00", 943=>x"7f00", 944=>x"6500", 945=>x"6700",
---- 946=>x"6600", 947=>x"6600", 948=>x"6800", 949=>x"6b00", 950=>x"6b00", 951=>x"7200", 952=>x"6800",
---- 953=>x"6500", 954=>x"6400", 955=>x"6700", 956=>x"6a00", 957=>x"6b00", 958=>x"6c00", 959=>x"7000",
---- 960=>x"6700", 961=>x"6600", 962=>x"6700", 963=>x"6900", 964=>x"6800", 965=>x"6b00", 966=>x"6d00",
---- 967=>x"6e00", 968=>x"6500", 969=>x"6800", 970=>x"6800", 971=>x"6400", 972=>x"6800", 973=>x"6b00",
---- 974=>x"6f00", 975=>x"7000", 976=>x"6400", 977=>x"9a00", 978=>x"6400", 979=>x"6700", 980=>x"6900",
---- 981=>x"6b00", 982=>x"6f00", 983=>x"7200", 984=>x"6800", 985=>x"6200", 986=>x"6600", 987=>x"6700",
---- 988=>x"6900", 989=>x"6900", 990=>x"6d00", 991=>x"7100", 992=>x"6700", 993=>x"6700", 994=>x"6700",
---- 995=>x"6500", 996=>x"6600", 997=>x"6800", 998=>x"6b00", 999=>x"7400", 1000=>x"6500", 1001=>x"6600",
---- 1002=>x"6600", 1003=>x"6400", 1004=>x"6700", 1005=>x"6b00", 1006=>x"6d00", 1007=>x"7100", 1008=>x"5f00",
---- 1009=>x"6300", 1010=>x"6500", 1011=>x"6600", 1012=>x"6700", 1013=>x"6800", 1014=>x"6a00", 1015=>x"6b00",
---- 1016=>x"6100", 1017=>x"6500", 1018=>x"6400", 1019=>x"6500", 1020=>x"6500", 1021=>x"6500", 1022=>x"6b00",
---- 1023=>x"6c00", 1024=>x"6400", 1025=>x"6500", 1026=>x"9f00", 1027=>x"6300", 1028=>x"6700", 1029=>x"6600",
---- 1030=>x"6800", 1031=>x"6900", 1032=>x"6200", 1033=>x"6000", 1034=>x"6300", 1035=>x"6100", 1036=>x"6000",
---- 1037=>x"6200", 1038=>x"6500", 1039=>x"8100", 1040=>x"6200", 1041=>x"6200", 1042=>x"6000", 1043=>x"5d00",
---- 1044=>x"5b00", 1045=>x"5c00", 1046=>x"7d00", 1047=>x"a000", 1048=>x"6200", 1049=>x"5f00", 1050=>x"5b00",
---- 1051=>x"5700", 1052=>x"5000", 1053=>x"7700", 1054=>x"c000", 1055=>x"ba00", 1056=>x"5f00", 1057=>x"5b00",
---- 1058=>x"5900", 1059=>x"5900", 1060=>x"4f00", 1061=>x"8f00", 1062=>x"ca00", 1063=>x"c000", 1064=>x"5f00",
---- 1065=>x"5d00", 1066=>x"5a00", 1067=>x"5b00", 1068=>x"4c00", 1069=>x"6b00", 1070=>x"b700", 1071=>x"ba00",
---- 1072=>x"6300", 1073=>x"6300", 1074=>x"6300", 1075=>x"5700", 1076=>x"3200", 1077=>x"5100", 1078=>x"ad00",
---- 1079=>x"6800", 1080=>x"7500", 1081=>x"6500", 1082=>x"4700", 1083=>x"4000", 1084=>x"2c00", 1085=>x"2c00",
---- 1086=>x"9100", 1087=>x"7a00", 1088=>x"6000", 1089=>x"3800", 1090=>x"3d00", 1091=>x"3900", 1092=>x"3d00",
---- 1093=>x"5600", 1094=>x"9500", 1095=>x"a000", 1096=>x"2a00", 1097=>x"2d00", 1098=>x"5800", 1099=>x"7800",
---- 1100=>x"8400", 1101=>x"9a00", 1102=>x"ac00", 1103=>x"bb00", 1104=>x"3600", 1105=>x"4f00", 1106=>x"8100",
---- 1107=>x"9e00", 1108=>x"9600", 1109=>x"9800", 1110=>x"9500", 1111=>x"a500", 1112=>x"6600", 1113=>x"8500",
---- 1114=>x"a200", 1115=>x"9b00", 1116=>x"8300", 1117=>x"8700", 1118=>x"7d00", 1119=>x"9700", 1120=>x"8a00",
---- 1121=>x"8300", 1122=>x"8600", 1123=>x"9800", 1124=>x"8600", 1125=>x"6800", 1126=>x"5100", 1127=>x"5700",
---- 1128=>x"a200", 1129=>x"a300", 1130=>x"9900", 1131=>x"8600", 1132=>x"5f00", 1133=>x"4500", 1134=>x"4100",
---- 1135=>x"4100", 1136=>x"a500", 1137=>x"8b00", 1138=>x"7900", 1139=>x"6c00", 1140=>x"4700", 1141=>x"3900",
---- 1142=>x"4500", 1143=>x"6300", 1144=>x"7600", 1145=>x"9700", 1146=>x"6b00", 1147=>x"5000", 1148=>x"4300",
---- 1149=>x"4f00", 1150=>x"6400", 1151=>x"5c00", 1152=>x"7600", 1153=>x"8b00", 1154=>x"7200", 1155=>x"7100",
---- 1156=>x"9100", 1157=>x"9100", 1158=>x"7200", 1159=>x"4200", 1160=>x"9e00", 1161=>x"ad00", 1162=>x"9a00",
---- 1163=>x"8a00", 1164=>x"7f00", 1165=>x"6a00", 1166=>x"4c00", 1167=>x"3d00", 1168=>x"9900", 1169=>x"7700",
---- 1170=>x"4600", 1171=>x"3b00", 1172=>x"4800", 1173=>x"4d00", 1174=>x"3700", 1175=>x"3b00", 1176=>x"5d00",
---- 1177=>x"3d00", 1178=>x"3400", 1179=>x"4c00", 1180=>x"aa00", 1181=>x"3f00", 1182=>x"3a00", 1183=>x"3e00",
---- 1184=>x"5e00", 1185=>x"5900", 1186=>x"5400", 1187=>x"5a00", 1188=>x"4e00", 1189=>x"3e00", 1190=>x"3f00",
---- 1191=>x"3400", 1192=>x"4c00", 1193=>x"5700", 1194=>x"6900", 1195=>x"5200", 1196=>x"5700", 1197=>x"5300",
---- 1198=>x"3800", 1199=>x"3900", 1200=>x"6f00", 1201=>x"7c00", 1202=>x"a300", 1203=>x"4b00", 1204=>x"7500",
---- 1205=>x"5b00", 1206=>x"4100", 1207=>x"5e00", 1208=>x"8800", 1209=>x"5c00", 1210=>x"4200", 1211=>x"6700",
---- 1212=>x"6a00", 1213=>x"4400", 1214=>x"6100", 1215=>x"7a00", 1216=>x"3b00", 1217=>x"4300", 1218=>x"7100",
---- 1219=>x"8000", 1220=>x"4b00", 1221=>x"5f00", 1222=>x"7e00", 1223=>x"3e00", 1224=>x"3800", 1225=>x"6a00",
---- 1226=>x"9c00", 1227=>x"7200", 1228=>x"5900", 1229=>x"7600", 1230=>x"4200", 1231=>x"2f00", 1232=>x"6200",
---- 1233=>x"8700", 1234=>x"7700", 1235=>x"5e00", 1236=>x"6f00", 1237=>x"3c00", 1238=>x"3a00", 1239=>x"3600",
---- 1240=>x"8800", 1241=>x"7200", 1242=>x"4d00", 1243=>x"5f00", 1244=>x"5100", 1245=>x"5e00", 1246=>x"4500",
---- 1247=>x"c500", 1248=>x"8a00", 1249=>x"5e00", 1250=>x"5200", 1251=>x"5c00", 1252=>x"5900", 1253=>x"4a00",
---- 1254=>x"4000", 1255=>x"5d00", 1256=>x"5b00", 1257=>x"4e00", 1258=>x"6600", 1259=>x"6500", 1260=>x"5800",
---- 1261=>x"4100", 1262=>x"5e00", 1263=>x"5600", 1264=>x"4e00", 1265=>x"4900", 1266=>x"7e00", 1267=>x"6100",
---- 1268=>x"4400", 1269=>x"5700", 1270=>x"4e00", 1271=>x"3b00", 1272=>x"5300", 1273=>x"6b00", 1274=>x"7a00",
---- 1275=>x"4e00", 1276=>x"5500", 1277=>x"4a00", 1278=>x"4a00", 1279=>x"3300", 1280=>x"6400", 1281=>x"7000",
---- 1282=>x"6b00", 1283=>x"5200", 1284=>x"4a00", 1285=>x"3700", 1286=>x"3b00", 1287=>x"5000", 1288=>x"5d00",
---- 1289=>x"7000", 1290=>x"7900", 1291=>x"5600", 1292=>x"4800", 1293=>x"2900", 1294=>x"3200", 1295=>x"8a00",
---- 1296=>x"5700", 1297=>x"8700", 1298=>x"7800", 1299=>x"5200", 1300=>x"3d00", 1301=>x"1e00", 1302=>x"4c00",
---- 1303=>x"9200", 1304=>x"5000", 1305=>x"5f00", 1306=>x"5c00", 1307=>x"4900", 1308=>x"2b00", 1309=>x"3100",
---- 1310=>x"8100", 1311=>x"7a00", 1312=>x"4c00", 1313=>x"4a00", 1314=>x"4800", 1315=>x"2900", 1316=>x"2b00",
---- 1317=>x"7000", 1318=>x"7e00", 1319=>x"4e00", 1320=>x"5200", 1321=>x"4600", 1322=>x"3900", 1323=>x"2500",
---- 1324=>x"5d00", 1325=>x"7b00", 1326=>x"4600", 1327=>x"3200", 1328=>x"4700", 1329=>x"4500", 1330=>x"3500",
---- 1331=>x"5300", 1332=>x"8900", 1333=>x"4e00", 1334=>x"2c00", 1335=>x"3100", 1336=>x"4700", 1337=>x"4c00",
---- 1338=>x"6000", 1339=>x"8600", 1340=>x"5c00", 1341=>x"3900", 1342=>x"3100", 1343=>x"3300", 1344=>x"4800",
---- 1345=>x"7500", 1346=>x"7c00", 1347=>x"5a00", 1348=>x"3800", 1349=>x"3300", 1350=>x"2f00", 1351=>x"3000",
---- 1352=>x"7100", 1353=>x"8600", 1354=>x"3e00", 1355=>x"2a00", 1356=>x"4900", 1357=>x"3a00", 1358=>x"3800",
---- 1359=>x"3200", 1360=>x"7e00", 1361=>x"6c00", 1362=>x"2800", 1363=>x"2f00", 1364=>x"4500", 1365=>x"4c00",
---- 1366=>x"4500", 1367=>x"3a00", 1368=>x"7700", 1369=>x"5600", 1370=>x"2e00", 1371=>x"3900", 1372=>x"3400",
---- 1373=>x"4e00", 1374=>x"4500", 1375=>x"b800", 1376=>x"6d00", 1377=>x"3d00", 1378=>x"3500", 1379=>x"3500",
---- 1380=>x"4400", 1381=>x"4300", 1382=>x"3a00", 1383=>x"4d00", 1384=>x"7a00", 1385=>x"4400", 1386=>x"3700",
---- 1387=>x"3c00", 1388=>x"4100", 1389=>x"4100", 1390=>x"3700", 1391=>x"4600", 1392=>x"5d00", 1393=>x"4d00",
---- 1394=>x"3600", 1395=>x"3d00", 1396=>x"4000", 1397=>x"4200", 1398=>x"3900", 1399=>x"3400", 1400=>x"3100",
---- 1401=>x"4100", 1402=>x"3f00", 1403=>x"3f00", 1404=>x"4200", 1405=>x"4d00", 1406=>x"3b00", 1407=>x"3500",
---- 1408=>x"2700", 1409=>x"ca00", 1410=>x"4600", 1411=>x"b800", 1412=>x"4400", 1413=>x"4500", 1414=>x"3c00",
---- 1415=>x"4900", 1416=>x"2f00", 1417=>x"3600", 1418=>x"3400", 1419=>x"3100", 1420=>x"4600", 1421=>x"4500",
---- 1422=>x"3b00", 1423=>x"5700", 1424=>x"3a00", 1425=>x"2a00", 1426=>x"2d00", 1427=>x"2700", 1428=>x"4900",
---- 1429=>x"5100", 1430=>x"3400", 1431=>x"5a00", 1432=>x"2d00", 1433=>x"2800", 1434=>x"2d00", 1435=>x"2d00",
---- 1436=>x"5d00", 1437=>x"4f00", 1438=>x"3600", 1439=>x"5400", 1440=>x"2e00", 1441=>x"3100", 1442=>x"2b00",
---- 1443=>x"3600", 1444=>x"6400", 1445=>x"4400", 1446=>x"5100", 1447=>x"4900", 1448=>x"2900", 1449=>x"3400",
---- 1450=>x"2c00", 1451=>x"4900", 1452=>x"6700", 1453=>x"3300", 1454=>x"5100", 1455=>x"5500", 1456=>x"3000",
---- 1457=>x"3000", 1458=>x"2400", 1459=>x"5c00", 1460=>x"5b00", 1461=>x"3100", 1462=>x"3600", 1463=>x"5700",
---- 1464=>x"2f00", 1465=>x"2c00", 1466=>x"2f00", 1467=>x"5e00", 1468=>x"4600", 1469=>x"3500", 1470=>x"2a00",
---- 1471=>x"3b00", 1472=>x"3100", 1473=>x"2400", 1474=>x"3600", 1475=>x"5a00", 1476=>x"3f00", 1477=>x"3e00",
---- 1478=>x"3700", 1479=>x"2600", 1480=>x"2e00", 1481=>x"2600", 1482=>x"3a00", 1483=>x"5c00", 1484=>x"3700",
---- 1485=>x"3f00", 1486=>x"3d00", 1487=>x"3300", 1488=>x"2900", 1489=>x"2600", 1490=>x"4300", 1491=>x"5c00",
---- 1492=>x"2e00", 1493=>x"3300", 1494=>x"4100", 1495=>x"2d00", 1496=>x"d600", 1497=>x"2500", 1498=>x"4a00",
---- 1499=>x"5d00", 1500=>x"3000", 1501=>x"2e00", 1502=>x"3d00", 1503=>x"3c00", 1504=>x"3200", 1505=>x"2500",
---- 1506=>x"4600", 1507=>x"5a00", 1508=>x"2e00", 1509=>x"3300", 1510=>x"3900", 1511=>x"4500", 1512=>x"3600",
---- 1513=>x"2c00", 1514=>x"4200", 1515=>x"5500", 1516=>x"3000", 1517=>x"3700", 1518=>x"3600", 1519=>x"3a00",
---- 1520=>x"3f00", 1521=>x"2f00", 1522=>x"3e00", 1523=>x"4c00", 1524=>x"3000", 1525=>x"3200", 1526=>x"3200",
---- 1527=>x"2b00", 1528=>x"4400", 1529=>x"3c00", 1530=>x"4300", 1531=>x"4700", 1532=>x"3300", 1533=>x"2d00",
---- 1534=>x"3500", 1535=>x"2400", 1536=>x"3f00", 1537=>x"3e00", 1538=>x"4700", 1539=>x"3f00", 1540=>x"3300",
---- 1541=>x"2a00", 1542=>x"3900", 1543=>x"2600", 1544=>x"3800", 1545=>x"4300", 1546=>x"3b00", 1547=>x"3300",
---- 1548=>x"3400", 1549=>x"2d00", 1550=>x"3300", 1551=>x"2900", 1552=>x"3800", 1553=>x"4600", 1554=>x"3500",
---- 1555=>x"3100", 1556=>x"3000", 1557=>x"2e00", 1558=>x"3000", 1559=>x"2800", 1560=>x"4700", 1561=>x"3d00",
---- 1562=>x"3200", 1563=>x"4200", 1564=>x"3300", 1565=>x"2b00", 1566=>x"3100", 1567=>x"2d00", 1568=>x"4b00",
---- 1569=>x"3800", 1570=>x"3400", 1571=>x"5100", 1572=>x"4100", 1573=>x"2f00", 1574=>x"3600", 1575=>x"2f00",
---- 1576=>x"3f00", 1577=>x"3600", 1578=>x"3600", 1579=>x"4e00", 1580=>x"5d00", 1581=>x"c700", 1582=>x"3800",
---- 1583=>x"3200", 1584=>x"3e00", 1585=>x"3300", 1586=>x"3400", 1587=>x"4d00", 1588=>x"7000", 1589=>x"4600",
---- 1590=>x"3d00", 1591=>x"3f00", 1592=>x"3400", 1593=>x"2800", 1594=>x"3100", 1595=>x"4200", 1596=>x"6c00",
---- 1597=>x"5400", 1598=>x"4400", 1599=>x"4100", 1600=>x"2900", 1601=>x"2100", 1602=>x"3100", 1603=>x"3b00",
---- 1604=>x"6a00", 1605=>x"6400", 1606=>x"4d00", 1607=>x"4800", 1608=>x"2500", 1609=>x"2100", 1610=>x"2900",
---- 1611=>x"3200", 1612=>x"7000", 1613=>x"7000", 1614=>x"4500", 1615=>x"5b00", 1616=>x"2900", 1617=>x"1c00",
---- 1618=>x"2100", 1619=>x"4b00", 1620=>x"8c00", 1621=>x"6200", 1622=>x"4400", 1623=>x"6600", 1624=>x"7100",
---- 1625=>x"5b00", 1626=>x"6700", 1627=>x"8800", 1628=>x"6d00", 1629=>x"4300", 1630=>x"4800", 1631=>x"4a00",
---- 1632=>x"6400", 1633=>x"7500", 1634=>x"7c00", 1635=>x"6000", 1636=>x"4200", 1637=>x"5200", 1638=>x"4300",
---- 1639=>x"3b00", 1640=>x"3100", 1641=>x"4c00", 1642=>x"4100", 1643=>x"3d00", 1644=>x"3c00", 1645=>x"c700",
---- 1646=>x"3a00", 1647=>x"4900", 1648=>x"3d00", 1649=>x"5800", 1650=>x"4400", 1651=>x"3a00", 1652=>x"3b00",
---- 1653=>x"3900", 1654=>x"c300", 1655=>x"3900", 1656=>x"3300", 1657=>x"3c00", 1658=>x"3300", 1659=>x"2d00",
---- 1660=>x"4400", 1661=>x"aa00", 1662=>x"4300", 1663=>x"3900", 1664=>x"2c00", 1665=>x"2f00", 1666=>x"2b00",
---- 1667=>x"2900", 1668=>x"5100", 1669=>x"6a00", 1670=>x"4300", 1671=>x"3b00", 1672=>x"3500", 1673=>x"2d00",
---- 1674=>x"2a00", 1675=>x"3000", 1676=>x"6100", 1677=>x"6a00", 1678=>x"3600", 1679=>x"4800", 1680=>x"3800",
---- 1681=>x"3100", 1682=>x"2a00", 1683=>x"3400", 1684=>x"6c00", 1685=>x"6b00", 1686=>x"2d00", 1687=>x"4000",
---- 1688=>x"3200", 1689=>x"3100", 1690=>x"2f00", 1691=>x"3500", 1692=>x"7100", 1693=>x"7300", 1694=>x"3000",
---- 1695=>x"3600", 1696=>x"2a00", 1697=>x"2d00", 1698=>x"2e00", 1699=>x"3700", 1700=>x"7400", 1701=>x"7000",
---- 1702=>x"2d00", 1703=>x"3700", 1704=>x"2d00", 1705=>x"2d00", 1706=>x"2a00", 1707=>x"3f00", 1708=>x"8500",
---- 1709=>x"6c00", 1710=>x"2200", 1711=>x"3300", 1712=>x"3300", 1713=>x"3100", 1714=>x"2b00", 1715=>x"5300",
---- 1716=>x"9400", 1717=>x"6600", 1718=>x"2600", 1719=>x"2500", 1720=>x"3000", 1721=>x"d300", 1722=>x"2e00",
---- 1723=>x"6e00", 1724=>x"9500", 1725=>x"5b00", 1726=>x"2700", 1727=>x"dd00", 1728=>x"2600", 1729=>x"2600",
---- 1730=>x"3d00", 1731=>x"7f00", 1732=>x"8800", 1733=>x"5400", 1734=>x"2a00", 1735=>x"2c00", 1736=>x"2200",
---- 1737=>x"2800", 1738=>x"7300", 1739=>x"8900", 1740=>x"7f00", 1741=>x"5800", 1742=>x"2b00", 1743=>x"2900",
---- 1744=>x"2800", 1745=>x"5a00", 1746=>x"8500", 1747=>x"6100", 1748=>x"7000", 1749=>x"3f00", 1750=>x"2800",
---- 1751=>x"2900", 1752=>x"6000", 1753=>x"7800", 1754=>x"4100", 1755=>x"4b00", 1756=>x"6a00", 1757=>x"3c00",
---- 1758=>x"3100", 1759=>x"2a00", 1760=>x"5900", 1761=>x"3a00", 1762=>x"2400", 1763=>x"6400", 1764=>x"6600",
---- 1765=>x"4b00", 1766=>x"3600", 1767=>x"2d00", 1768=>x"2d00", 1769=>x"2a00", 1770=>x"3300", 1771=>x"5a00",
---- 1772=>x"5600", 1773=>x"5700", 1774=>x"3600", 1775=>x"3000", 1776=>x"2f00", 1777=>x"3400", 1778=>x"3200",
---- 1779=>x"5000", 1780=>x"5600", 1781=>x"5500", 1782=>x"3800", 1783=>x"2e00", 1784=>x"3b00", 1785=>x"3400",
---- 1786=>x"2c00", 1787=>x"4c00", 1788=>x"5300", 1789=>x"4300", 1790=>x"3900", 1791=>x"3100", 1792=>x"3900",
---- 1793=>x"2d00", 1794=>x"3300", 1795=>x"4600", 1796=>x"4700", 1797=>x"3b00", 1798=>x"3100", 1799=>x"3500",
---- 1800=>x"3200", 1801=>x"3000", 1802=>x"3100", 1803=>x"3f00", 1804=>x"4300", 1805=>x"3d00", 1806=>x"3d00",
---- 1807=>x"3d00", 1808=>x"2f00", 1809=>x"2d00", 1810=>x"2e00", 1811=>x"3f00", 1812=>x"3c00", 1813=>x"3800",
---- 1814=>x"4000", 1815=>x"3700", 1816=>x"2a00", 1817=>x"2c00", 1818=>x"3a00", 1819=>x"4200", 1820=>x"3e00",
---- 1821=>x"3b00", 1822=>x"3100", 1823=>x"2d00", 1824=>x"2b00", 1825=>x"2c00", 1826=>x"4100", 1827=>x"3d00",
---- 1828=>x"4200", 1829=>x"3500", 1830=>x"3200", 1831=>x"3800", 1832=>x"2d00", 1833=>x"3300", 1834=>x"3d00",
---- 1835=>x"3d00", 1836=>x"4900", 1837=>x"3a00", 1838=>x"3300", 1839=>x"3d00", 1840=>x"2c00", 1841=>x"3d00",
---- 1842=>x"3900", 1843=>x"4000", 1844=>x"3b00", 1845=>x"3600", 1846=>x"3700", 1847=>x"4d00", 1848=>x"3600",
---- 1849=>x"4300", 1850=>x"3700", 1851=>x"4500", 1852=>x"3400", 1853=>x"3200", 1854=>x"3c00", 1855=>x"5100",
---- 1856=>x"4400", 1857=>x"3500", 1858=>x"3a00", 1859=>x"4100", 1860=>x"3200", 1861=>x"3200", 1862=>x"3c00",
---- 1863=>x"3f00", 1864=>x"3f00", 1865=>x"2d00", 1866=>x"3e00", 1867=>x"3d00", 1868=>x"3000", 1869=>x"cb00",
---- 1870=>x"4000", 1871=>x"4100", 1872=>x"3300", 1873=>x"d200", 1874=>x"4100", 1875=>x"3d00", 1876=>x"2e00",
---- 1877=>x"2f00", 1878=>x"3d00", 1879=>x"4300", 1880=>x"2e00", 1881=>x"2c00", 1882=>x"4700", 1883=>x"3d00",
---- 1884=>x"2e00", 1885=>x"3100", 1886=>x"3f00", 1887=>x"3e00", 1888=>x"3600", 1889=>x"2d00", 1890=>x"3f00",
---- 1891=>x"3800", 1892=>x"2a00", 1893=>x"3600", 1894=>x"4900", 1895=>x"3b00", 1896=>x"3300", 1897=>x"2c00",
---- 1898=>x"3400", 1899=>x"3e00", 1900=>x"2e00", 1901=>x"3700", 1902=>x"4500", 1903=>x"3d00", 1904=>x"3300",
---- 1905=>x"3100", 1906=>x"3100", 1907=>x"3d00", 1908=>x"3500", 1909=>x"3f00", 1910=>x"3e00", 1911=>x"3800",
---- 1912=>x"3200", 1913=>x"3100", 1914=>x"3200", 1915=>x"3300", 1916=>x"3800", 1917=>x"4600", 1918=>x"3400",
---- 1919=>x"3b00", 1920=>x"3a00", 1921=>x"3100", 1922=>x"3200", 1923=>x"2b00", 1924=>x"3200", 1925=>x"3400",
---- 1926=>x"2f00", 1927=>x"4000", 1928=>x"3c00", 1929=>x"3000", 1930=>x"3300", 1931=>x"3300", 1932=>x"2d00",
---- 1933=>x"2800", 1934=>x"3400", 1935=>x"3f00", 1936=>x"3a00", 1937=>x"2d00", 1938=>x"3100", 1939=>x"3000",
---- 1940=>x"2d00", 1941=>x"3700", 1942=>x"4500", 1943=>x"4500", 1944=>x"3c00", 1945=>x"3000", 1946=>x"2b00",
---- 1947=>x"2c00", 1948=>x"2e00", 1949=>x"3900", 1950=>x"5100", 1951=>x"4e00", 1952=>x"4800", 1953=>x"4000",
---- 1954=>x"2b00", 1955=>x"2d00", 1956=>x"2e00", 1957=>x"3900", 1958=>x"4c00", 1959=>x"5100", 1960=>x"4800",
---- 1961=>x"3e00", 1962=>x"d400", 1963=>x"3400", 1964=>x"2e00", 1965=>x"3e00", 1966=>x"4800", 1967=>x"4d00",
---- 1968=>x"4f00", 1969=>x"3e00", 1970=>x"2800", 1971=>x"3300", 1972=>x"3000", 1973=>x"3c00", 1974=>x"3c00",
---- 1975=>x"5000", 1976=>x"5400", 1977=>x"4800", 1978=>x"2900", 1979=>x"3500", 1980=>x"3000", 1981=>x"3b00",
---- 1982=>x"3f00", 1983=>x"5b00", 1984=>x"4700", 1985=>x"5900", 1986=>x"2a00", 1987=>x"2f00", 1988=>x"2f00",
---- 1989=>x"3700", 1990=>x"4e00", 1991=>x"5f00", 1992=>x"3500", 1993=>x"5800", 1994=>x"3900", 1995=>x"2c00",
---- 1996=>x"2c00", 1997=>x"2e00", 1998=>x"4e00", 1999=>x"5c00", 2000=>x"d000", 2001=>x"4d00", 2002=>x"5300",
---- 2003=>x"2900", 2004=>x"2e00", 2005=>x"2b00", 2006=>x"6000", 2007=>x"6800", 2008=>x"3400", 2009=>x"3700",
---- 2010=>x"5c00", 2011=>x"2f00", 2012=>x"2700", 2013=>x"3000", 2014=>x"7600", 2015=>x"6c00", 2016=>x"3f00",
---- 2017=>x"2800", 2018=>x"5400", 2019=>x"4800", 2020=>x"2800", 2021=>x"3300", 2022=>x"8000", 2023=>x"5b00",
---- 2024=>x"4a00", 2025=>x"3400", 2026=>x"3b00", 2027=>x"4e00", 2028=>x"3300", 2029=>x"3e00", 2030=>x"7c00",
---- 2031=>x"4d00", 2032=>x"4f00", 2033=>x"3900", 2034=>x"3000", 2035=>x"4300", 2036=>x"4100", 2037=>x"5e00",
---- 2038=>x"7f00", 2039=>x"3400", 2040=>x"4c00", 2041=>x"4400", 2042=>x"3200", 2043=>x"4c00", 2044=>x"5600",
---- 2045=>x"7e00", 2046=>x"6d00", 2047=>x"2e00"),
---- 7  => (0=>x"7400", 1=>x"8500", 2=>x"7c00", 3=>x"7900", 4=>x"7d00", 5=>x"8000", 6=>x"7a00", 7=>x"8300",
---- 8=>x"7500", 9=>x"7a00", 10=>x"7a00", 11=>x"7900", 12=>x"7f00", 13=>x"8000", 14=>x"7b00",
---- 15=>x"8300", 16=>x"7500", 17=>x"7900", 18=>x"7b00", 19=>x"7a00", 20=>x"7e00", 21=>x"8000",
---- 22=>x"7b00", 23=>x"8100", 24=>x"8900", 25=>x"7900", 26=>x"7d00", 27=>x"7c00", 28=>x"7d00",
---- 29=>x"7b00", 30=>x"7c00", 31=>x"7c00", 32=>x"7700", 33=>x"7a00", 34=>x"7a00", 35=>x"7c00",
---- 36=>x"7d00", 37=>x"7d00", 38=>x"7b00", 39=>x"7c00", 40=>x"7400", 41=>x"7900", 42=>x"7b00",
---- 43=>x"7c00", 44=>x"7b00", 45=>x"7c00", 46=>x"7d00", 47=>x"8000", 48=>x"7700", 49=>x"7500",
---- 50=>x"7a00", 51=>x"7a00", 52=>x"7a00", 53=>x"7d00", 54=>x"7f00", 55=>x"7d00", 56=>x"7600",
---- 57=>x"7600", 58=>x"7a00", 59=>x"7800", 60=>x"7d00", 61=>x"7c00", 62=>x"7d00", 63=>x"8000",
---- 64=>x"7300", 65=>x"7800", 66=>x"7a00", 67=>x"7d00", 68=>x"7c00", 69=>x"7e00", 70=>x"7f00",
---- 71=>x"8000", 72=>x"7700", 73=>x"7700", 74=>x"7800", 75=>x"7a00", 76=>x"7b00", 77=>x"7d00",
---- 78=>x"7a00", 79=>x"7f00", 80=>x"7700", 81=>x"7800", 82=>x"7800", 83=>x"7700", 84=>x"7c00",
---- 85=>x"7c00", 86=>x"7a00", 87=>x"7d00", 88=>x"7400", 89=>x"7600", 90=>x"7700", 91=>x"7900",
---- 92=>x"7b00", 93=>x"7d00", 94=>x"7d00", 95=>x"7b00", 96=>x"7500", 97=>x"7900", 98=>x"7a00",
---- 99=>x"7800", 100=>x"7800", 101=>x"7800", 102=>x"7f00", 103=>x"7f00", 104=>x"7700", 105=>x"7900",
---- 106=>x"7700", 107=>x"7a00", 108=>x"7a00", 109=>x"7c00", 110=>x"7b00", 111=>x"7d00", 112=>x"7500",
---- 113=>x"7a00", 114=>x"7800", 115=>x"7800", 116=>x"7c00", 117=>x"7d00", 118=>x"7c00", 119=>x"7f00",
---- 120=>x"7400", 121=>x"7600", 122=>x"7a00", 123=>x"7a00", 124=>x"7a00", 125=>x"7c00", 126=>x"7d00",
---- 127=>x"7b00", 128=>x"7500", 129=>x"7700", 130=>x"7a00", 131=>x"7900", 132=>x"7c00", 133=>x"7800",
---- 134=>x"7a00", 135=>x"8200", 136=>x"7400", 137=>x"7500", 138=>x"7800", 139=>x"7a00", 140=>x"7c00",
---- 141=>x"7c00", 142=>x"7b00", 143=>x"7e00", 144=>x"7700", 145=>x"7400", 146=>x"7800", 147=>x"7800",
---- 148=>x"7600", 149=>x"7800", 150=>x"7d00", 151=>x"7b00", 152=>x"7300", 153=>x"7300", 154=>x"7900",
---- 155=>x"7900", 156=>x"7600", 157=>x"7700", 158=>x"7a00", 159=>x"7c00", 160=>x"7400", 161=>x"7700",
---- 162=>x"7700", 163=>x"7900", 164=>x"7900", 165=>x"7a00", 166=>x"7700", 167=>x"7800", 168=>x"7500",
---- 169=>x"7a00", 170=>x"7800", 171=>x"7700", 172=>x"7600", 173=>x"8500", 174=>x"8300", 175=>x"7a00",
---- 176=>x"7500", 177=>x"7800", 178=>x"7800", 179=>x"7800", 180=>x"7700", 181=>x"7a00", 182=>x"7d00",
---- 183=>x"7b00", 184=>x"7500", 185=>x"7800", 186=>x"7800", 187=>x"7900", 188=>x"7a00", 189=>x"7c00",
---- 190=>x"7a00", 191=>x"7b00", 192=>x"7200", 193=>x"7700", 194=>x"7900", 195=>x"7a00", 196=>x"8700",
---- 197=>x"7c00", 198=>x"7c00", 199=>x"7c00", 200=>x"7400", 201=>x"7900", 202=>x"7900", 203=>x"7900",
---- 204=>x"7800", 205=>x"8500", 206=>x"7e00", 207=>x"7c00", 208=>x"7600", 209=>x"7800", 210=>x"7900",
---- 211=>x"7b00", 212=>x"7800", 213=>x"7800", 214=>x"7a00", 215=>x"7c00", 216=>x"7500", 217=>x"7a00",
---- 218=>x"7900", 219=>x"7a00", 220=>x"7c00", 221=>x"7a00", 222=>x"7b00", 223=>x"7e00", 224=>x"7600",
---- 225=>x"7800", 226=>x"7800", 227=>x"7700", 228=>x"7a00", 229=>x"7a00", 230=>x"7e00", 231=>x"7b00",
---- 232=>x"7400", 233=>x"7500", 234=>x"7600", 235=>x"7900", 236=>x"7a00", 237=>x"7900", 238=>x"7b00",
---- 239=>x"7a00", 240=>x"7500", 241=>x"7500", 242=>x"7500", 243=>x"7500", 244=>x"7800", 245=>x"7b00",
---- 246=>x"7900", 247=>x"7900", 248=>x"7500", 249=>x"7500", 250=>x"7500", 251=>x"7500", 252=>x"7700",
---- 253=>x"7a00", 254=>x"7900", 255=>x"7700", 256=>x"7300", 257=>x"7500", 258=>x"7500", 259=>x"7200",
---- 260=>x"7800", 261=>x"7700", 262=>x"7900", 263=>x"7600", 264=>x"7000", 265=>x"7400", 266=>x"7500",
---- 267=>x"7200", 268=>x"7700", 269=>x"7400", 270=>x"7300", 271=>x"7500", 272=>x"7000", 273=>x"7100",
---- 274=>x"7000", 275=>x"8e00", 276=>x"7200", 277=>x"8900", 278=>x"7500", 279=>x"7600", 280=>x"7200",
---- 281=>x"7600", 282=>x"6f00", 283=>x"7100", 284=>x"7400", 285=>x"7500", 286=>x"7600", 287=>x"7700",
---- 288=>x"7100", 289=>x"7200", 290=>x"7200", 291=>x"7400", 292=>x"7300", 293=>x"7500", 294=>x"7300",
---- 295=>x"7600", 296=>x"7100", 297=>x"6f00", 298=>x"7300", 299=>x"8b00", 300=>x"7100", 301=>x"7200",
---- 302=>x"7400", 303=>x"7600", 304=>x"6d00", 305=>x"7100", 306=>x"7200", 307=>x"7600", 308=>x"8d00",
---- 309=>x"7300", 310=>x"7500", 311=>x"7a00", 312=>x"7200", 313=>x"7500", 314=>x"7400", 315=>x"7300",
---- 316=>x"7200", 317=>x"7100", 318=>x"7200", 319=>x"7400", 320=>x"7000", 321=>x"7200", 322=>x"7700",
---- 323=>x"7100", 324=>x"7400", 325=>x"7400", 326=>x"7800", 327=>x"7700", 328=>x"6e00", 329=>x"7000",
---- 330=>x"7200", 331=>x"7200", 332=>x"7100", 333=>x"7400", 334=>x"7500", 335=>x"7900", 336=>x"7100",
---- 337=>x"7500", 338=>x"7100", 339=>x"7300", 340=>x"7500", 341=>x"7500", 342=>x"7600", 343=>x"7600",
---- 344=>x"7000", 345=>x"7200", 346=>x"7200", 347=>x"7200", 348=>x"7400", 349=>x"7500", 350=>x"7500",
---- 351=>x"7600", 352=>x"6d00", 353=>x"7200", 354=>x"7300", 355=>x"7400", 356=>x"7500", 357=>x"7300",
---- 358=>x"7600", 359=>x"7800", 360=>x"6f00", 361=>x"7200", 362=>x"7400", 363=>x"7300", 364=>x"7400",
---- 365=>x"7500", 366=>x"7800", 367=>x"7b00", 368=>x"7000", 369=>x"7000", 370=>x"7400", 371=>x"7600",
---- 372=>x"7400", 373=>x"7600", 374=>x"7800", 375=>x"7800", 376=>x"7400", 377=>x"7200", 378=>x"7300",
---- 379=>x"7400", 380=>x"7400", 381=>x"7600", 382=>x"7700", 383=>x"7600", 384=>x"7000", 385=>x"7000",
---- 386=>x"7700", 387=>x"7800", 388=>x"7300", 389=>x"7400", 390=>x"7500", 391=>x"7500", 392=>x"7000",
---- 393=>x"7300", 394=>x"7900", 395=>x"7500", 396=>x"7400", 397=>x"7200", 398=>x"7600", 399=>x"7800",
---- 400=>x"6d00", 401=>x"7100", 402=>x"7400", 403=>x"7200", 404=>x"7200", 405=>x"7700", 406=>x"7700",
---- 407=>x"7500", 408=>x"7000", 409=>x"7400", 410=>x"7400", 411=>x"7600", 412=>x"7600", 413=>x"7600",
---- 414=>x"7600", 415=>x"7600", 416=>x"6e00", 417=>x"7100", 418=>x"7400", 419=>x"7500", 420=>x"7700",
---- 421=>x"7a00", 422=>x"7800", 423=>x"7300", 424=>x"7100", 425=>x"7000", 426=>x"7100", 427=>x"7500",
---- 428=>x"7600", 429=>x"7400", 430=>x"7500", 431=>x"7200", 432=>x"7300", 433=>x"7300", 434=>x"7600",
---- 435=>x"7300", 436=>x"7000", 437=>x"7300", 438=>x"7200", 439=>x"7100", 440=>x"7100", 441=>x"7200",
---- 442=>x"7000", 443=>x"7300", 444=>x"7500", 445=>x"7400", 446=>x"6e00", 447=>x"6b00", 448=>x"6d00",
---- 449=>x"7200", 450=>x"7300", 451=>x"7200", 452=>x"6f00", 453=>x"6e00", 454=>x"6d00", 455=>x"6700",
---- 456=>x"6e00", 457=>x"7000", 458=>x"7200", 459=>x"8d00", 460=>x"6f00", 461=>x"6f00", 462=>x"6b00",
---- 463=>x"6b00", 464=>x"6d00", 465=>x"7100", 466=>x"6f00", 467=>x"6f00", 468=>x"6c00", 469=>x"6b00",
---- 470=>x"6100", 471=>x"8300", 472=>x"6a00", 473=>x"6d00", 474=>x"6e00", 475=>x"6e00", 476=>x"6b00",
---- 477=>x"6500", 478=>x"6100", 479=>x"a700", 480=>x"6c00", 481=>x"6f00", 482=>x"7000", 483=>x"6c00",
---- 484=>x"6e00", 485=>x"6500", 486=>x"6f00", 487=>x"c700", 488=>x"6d00", 489=>x"7200", 490=>x"7000",
---- 491=>x"6e00", 492=>x"6c00", 493=>x"6200", 494=>x"8000", 495=>x"d100", 496=>x"6c00", 497=>x"7100",
---- 498=>x"7200", 499=>x"7500", 500=>x"6d00", 501=>x"5f00", 502=>x"9e00", 503=>x"dc00", 504=>x"7000",
---- 505=>x"7000", 506=>x"7300", 507=>x"7300", 508=>x"6e00", 509=>x"6500", 510=>x"b000", 511=>x"d600",
---- 512=>x"6e00", 513=>x"7000", 514=>x"7100", 515=>x"6c00", 516=>x"6400", 517=>x"6900", 518=>x"c400",
---- 519=>x"d100", 520=>x"6f00", 521=>x"7100", 522=>x"6f00", 523=>x"6d00", 524=>x"6400", 525=>x"7300",
---- 526=>x"cf00", 527=>x"cf00", 528=>x"7100", 529=>x"7200", 530=>x"7300", 531=>x"6c00", 532=>x"5f00",
---- 533=>x"8700", 534=>x"d800", 535=>x"cc00", 536=>x"7000", 537=>x"7200", 538=>x"7200", 539=>x"6d00",
---- 540=>x"6000", 541=>x"9a00", 542=>x"2400", 543=>x"ca00", 544=>x"6f00", 545=>x"7000", 546=>x"6e00",
---- 547=>x"6800", 548=>x"5b00", 549=>x"ab00", 550=>x"df00", 551=>x"bf00", 552=>x"7000", 553=>x"6d00",
---- 554=>x"6900", 555=>x"6300", 556=>x"5d00", 557=>x"b700", 558=>x"db00", 559=>x"ac00", 560=>x"6900",
---- 561=>x"6c00", 562=>x"6c00", 563=>x"5e00", 564=>x"6a00", 565=>x"cb00", 566=>x"d400", 567=>x"a400",
---- 568=>x"6a00", 569=>x"6900", 570=>x"6700", 571=>x"5800", 572=>x"7900", 573=>x"d800", 574=>x"cb00",
---- 575=>x"ad00", 576=>x"6900", 577=>x"6800", 578=>x"6200", 579=>x"5400", 580=>x"8d00", 581=>x"de00",
---- 582=>x"c900", 583=>x"aa00", 584=>x"6900", 585=>x"6600", 586=>x"6000", 587=>x"5300", 588=>x"a500",
---- 589=>x"de00", 590=>x"c300", 591=>x"af00", 592=>x"6700", 593=>x"6500", 594=>x"5e00", 595=>x"5b00",
---- 596=>x"bb00", 597=>x"dd00", 598=>x"c200", 599=>x"b000", 600=>x"6500", 601=>x"6700", 602=>x"5b00",
---- 603=>x"5e00", 604=>x"c000", 605=>x"db00", 606=>x"bb00", 607=>x"b700", 608=>x"6700", 609=>x"6600",
---- 610=>x"5b00", 611=>x"6200", 612=>x"c800", 613=>x"d500", 614=>x"be00", 615=>x"af00", 616=>x"6600",
---- 617=>x"6500", 618=>x"5b00", 619=>x"6700", 620=>x"2f00", 621=>x"d500", 622=>x"bb00", 623=>x"b200",
---- 624=>x"6600", 625=>x"6400", 626=>x"5a00", 627=>x"6300", 628=>x"cc00", 629=>x"d000", 630=>x"b900",
---- 631=>x"ad00", 632=>x"6500", 633=>x"6500", 634=>x"5900", 635=>x"6600", 636=>x"d200", 637=>x"cc00",
---- 638=>x"ba00", 639=>x"b100", 640=>x"6100", 641=>x"6200", 642=>x"5500", 643=>x"6b00", 644=>x"d100",
---- 645=>x"c300", 646=>x"bb00", 647=>x"ad00", 648=>x"6100", 649=>x"5e00", 650=>x"5200", 651=>x"7300",
---- 652=>x"d700", 653=>x"c500", 654=>x"b200", 655=>x"b100", 656=>x"6000", 657=>x"5c00", 658=>x"5000",
---- 659=>x"8100", 660=>x"db00", 661=>x"ba00", 662=>x"b900", 663=>x"ad00", 664=>x"5e00", 665=>x"5c00",
---- 666=>x"4b00", 667=>x"8c00", 668=>x"d500", 669=>x"c300", 670=>x"b600", 671=>x"bd00", 672=>x"5d00",
---- 673=>x"5a00", 674=>x"4b00", 675=>x"9d00", 676=>x"db00", 677=>x"c100", 678=>x"c500", 679=>x"b400",
---- 680=>x"5d00", 681=>x"5600", 682=>x"4900", 683=>x"9800", 684=>x"da00", 685=>x"cc00", 686=>x"be00",
---- 687=>x"c100", 688=>x"5c00", 689=>x"5500", 690=>x"4800", 691=>x"9b00", 692=>x"e000", 693=>x"c500",
---- 694=>x"c800", 695=>x"bd00", 696=>x"5f00", 697=>x"5700", 698=>x"4600", 699=>x"9500", 700=>x"dc00",
---- 701=>x"3100", 702=>x"c400", 703=>x"c400", 704=>x"5b00", 705=>x"5500", 706=>x"4700", 707=>x"9000",
---- 708=>x"1d00", 709=>x"c700", 710=>x"c400", 711=>x"c700", 712=>x"5900", 713=>x"5800", 714=>x"4800",
---- 715=>x"8c00", 716=>x"db00", 717=>x"ce00", 718=>x"c800", 719=>x"c000", 720=>x"5f00", 721=>x"5b00",
---- 722=>x"4900", 723=>x"7b00", 724=>x"dd00", 725=>x"ce00", 726=>x"c400", 727=>x"c800", 728=>x"6000",
---- 729=>x"5b00", 730=>x"5000", 731=>x"6600", 732=>x"ce00", 733=>x"2e00", 734=>x"c900", 735=>x"c100",
---- 736=>x"5f00", 737=>x"5b00", 738=>x"5000", 739=>x"5200", 740=>x"bb00", 741=>x"d900", 742=>x"c600",
---- 743=>x"ce00", 744=>x"5c00", 745=>x"5a00", 746=>x"5200", 747=>x"4b00", 748=>x"ab00", 749=>x"da00",
---- 750=>x"cf00", 751=>x"c700", 752=>x"5f00", 753=>x"5f00", 754=>x"5900", 755=>x"4900", 756=>x"8a00",
---- 757=>x"e000", 758=>x"c200", 759=>x"d000", 760=>x"6300", 761=>x"5f00", 762=>x"5c00", 763=>x"4900",
---- 764=>x"6c00", 765=>x"d200", 766=>x"d200", 767=>x"c500", 768=>x"6400", 769=>x"6000", 770=>x"5b00",
---- 771=>x"5100", 772=>x"4f00", 773=>x"ba00", 774=>x"d900", 775=>x"ca00", 776=>x"6500", 777=>x"6400",
---- 778=>x"5e00", 779=>x"5600", 780=>x"4900", 781=>x"8d00", 782=>x"dd00", 783=>x"c500", 784=>x"6400",
---- 785=>x"6500", 786=>x"6000", 787=>x"5700", 788=>x"4a00", 789=>x"7300", 790=>x"da00", 791=>x"ce00",
---- 792=>x"6500", 793=>x"6400", 794=>x"6200", 795=>x"5d00", 796=>x"5200", 797=>x"5c00", 798=>x"c300",
---- 799=>x"d300", 800=>x"9300", 801=>x"6700", 802=>x"6500", 803=>x"6100", 804=>x"5b00", 805=>x"5100",
---- 806=>x"8100", 807=>x"dd00", 808=>x"6700", 809=>x"6a00", 810=>x"9800", 811=>x"6500", 812=>x"6000",
---- 813=>x"5500", 814=>x"5a00", 815=>x"bb00", 816=>x"6800", 817=>x"6b00", 818=>x"6700", 819=>x"6500",
---- 820=>x"6400", 821=>x"5f00", 822=>x"5100", 823=>x"7500", 824=>x"6b00", 825=>x"6800", 826=>x"6a00",
---- 827=>x"6900", 828=>x"6600", 829=>x"5f00", 830=>x"5b00", 831=>x"5000", 832=>x"6c00", 833=>x"6a00",
---- 834=>x"6c00", 835=>x"6d00", 836=>x"6a00", 837=>x"6600", 838=>x"5f00", 839=>x"5100", 840=>x"6c00",
---- 841=>x"6f00", 842=>x"7000", 843=>x"6c00", 844=>x"6b00", 845=>x"6900", 846=>x"6200", 847=>x"5c00",
---- 848=>x"6b00", 849=>x"6d00", 850=>x"7200", 851=>x"7100", 852=>x"6c00", 853=>x"6900", 854=>x"6500",
---- 855=>x"5f00", 856=>x"6b00", 857=>x"7200", 858=>x"7100", 859=>x"6e00", 860=>x"6d00", 861=>x"9200",
---- 862=>x"6900", 863=>x"5f00", 864=>x"6c00", 865=>x"7000", 866=>x"7100", 867=>x"7000", 868=>x"6e00",
---- 869=>x"6b00", 870=>x"6800", 871=>x"6200", 872=>x"6f00", 873=>x"7200", 874=>x"7400", 875=>x"7300",
---- 876=>x"6f00", 877=>x"6d00", 878=>x"6a00", 879=>x"6500", 880=>x"6f00", 881=>x"7100", 882=>x"7100",
---- 883=>x"7100", 884=>x"7100", 885=>x"6f00", 886=>x"6d00", 887=>x"6600", 888=>x"6b00", 889=>x"6b00",
---- 890=>x"7200", 891=>x"7500", 892=>x"7100", 893=>x"6d00", 894=>x"7000", 895=>x"6800", 896=>x"7600",
---- 897=>x"7b00", 898=>x"6e00", 899=>x"7600", 900=>x"7100", 901=>x"7200", 902=>x"7000", 903=>x"6d00",
---- 904=>x"a500", 905=>x"7a00", 906=>x"6d00", 907=>x"7500", 908=>x"7100", 909=>x"7100", 910=>x"6f00",
---- 911=>x"6c00", 912=>x"8200", 913=>x"6d00", 914=>x"7400", 915=>x"7300", 916=>x"7300", 917=>x"7200",
---- 918=>x"7300", 919=>x"7400", 920=>x"6c00", 921=>x"7300", 922=>x"7300", 923=>x"7400", 924=>x"7500",
---- 925=>x"7500", 926=>x"7300", 927=>x"7300", 928=>x"7300", 929=>x"7100", 930=>x"7100", 931=>x"7900",
---- 932=>x"7700", 933=>x"7700", 934=>x"7500", 935=>x"7500", 936=>x"7500", 937=>x"7300", 938=>x"7300",
---- 939=>x"7900", 940=>x"7800", 941=>x"7800", 942=>x"7900", 943=>x"7900", 944=>x"7400", 945=>x"7300",
---- 946=>x"7300", 947=>x"7400", 948=>x"7700", 949=>x"7400", 950=>x"7500", 951=>x"7500", 952=>x"8a00",
---- 953=>x"7600", 954=>x"7200", 955=>x"7000", 956=>x"6f00", 957=>x"6e00", 958=>x"6d00", 959=>x"6b00",
---- 960=>x"8c00", 961=>x"7600", 962=>x"7800", 963=>x"7800", 964=>x"7500", 965=>x"7900", 966=>x"7600",
---- 967=>x"7600", 968=>x"8e00", 969=>x"7300", 970=>x"7300", 971=>x"7700", 972=>x"7700", 973=>x"7900",
---- 974=>x"7800", 975=>x"7600", 976=>x"7100", 977=>x"7600", 978=>x"7500", 979=>x"7700", 980=>x"7800",
---- 981=>x"7700", 982=>x"7500", 983=>x"8300", 984=>x"7500", 985=>x"7700", 986=>x"7600", 987=>x"7700",
---- 988=>x"7700", 989=>x"7900", 990=>x"7200", 991=>x"b500", 992=>x"7700", 993=>x"7500", 994=>x"7700",
---- 995=>x"8600", 996=>x"8300", 997=>x"7a00", 998=>x"7900", 999=>x"b300", 1000=>x"7200", 1001=>x"7200",
---- 1002=>x"7600", 1003=>x"7400", 1004=>x"7b00", 1005=>x"8400", 1006=>x"8700", 1007=>x"8d00", 1008=>x"6d00",
---- 1009=>x"7400", 1010=>x"7200", 1011=>x"7900", 1012=>x"8e00", 1013=>x"9a00", 1014=>x"9100", 1015=>x"8700",
---- 1016=>x"6b00", 1017=>x"9300", 1018=>x"7000", 1019=>x"8c00", 1020=>x"9b00", 1021=>x"9d00", 1022=>x"9600",
---- 1023=>x"9000", 1024=>x"6f00", 1025=>x"7900", 1026=>x"8700", 1027=>x"8e00", 1028=>x"9800", 1029=>x"9d00",
---- 1030=>x"9a00", 1031=>x"9700", 1032=>x"6f00", 1033=>x"9f00", 1034=>x"9200", 1035=>x"9100", 1036=>x"9700",
---- 1037=>x"9b00", 1038=>x"9a00", 1039=>x"9800", 1040=>x"c300", 1041=>x"b200", 1042=>x"8100", 1043=>x"9500",
---- 1044=>x"9300", 1045=>x"6800", 1046=>x"9900", 1047=>x"9b00", 1048=>x"d400", 1049=>x"9200", 1050=>x"8200",
---- 1051=>x"9100", 1052=>x"9300", 1053=>x"9800", 1054=>x"9e00", 1055=>x"9000", 1056=>x"b300", 1057=>x"7800",
---- 1058=>x"8800", 1059=>x"9100", 1060=>x"9600", 1061=>x"9b00", 1062=>x"9800", 1063=>x"6900", 1064=>x"b900",
---- 1065=>x"9800", 1066=>x"8a00", 1067=>x"9200", 1068=>x"9500", 1069=>x"9700", 1070=>x"9200", 1071=>x"7200",
---- 1072=>x"7500", 1073=>x"b600", 1074=>x"b700", 1075=>x"9b00", 1076=>x"9400", 1077=>x"9a00", 1078=>x"8600",
---- 1079=>x"6100", 1080=>x"7900", 1081=>x"b000", 1082=>x"cf00", 1083=>x"cf00", 1084=>x"c000", 1085=>x"9400",
---- 1086=>x"4300", 1087=>x"2700", 1088=>x"a900", 1089=>x"be00", 1090=>x"e100", 1091=>x"f900", 1092=>x"bf00",
---- 1093=>x"4f00", 1094=>x"3f00", 1095=>x"2a00", 1096=>x"a000", 1097=>x"d200", 1098=>x"d700", 1099=>x"8800",
---- 1100=>x"3d00", 1101=>x"2d00", 1102=>x"5c00", 1103=>x"3400", 1104=>x"b700", 1105=>x"ae00", 1106=>x"4e00",
---- 1107=>x"2a00", 1108=>x"2e00", 1109=>x"2a00", 1110=>x"5200", 1111=>x"6400", 1112=>x"9300", 1113=>x"4b00",
---- 1114=>x"3a00", 1115=>x"4300", 1116=>x"3500", 1117=>x"3200", 1118=>x"3a00", 1119=>x"7300", 1120=>x"5600",
---- 1121=>x"5000", 1122=>x"3e00", 1123=>x"3000", 1124=>x"2800", 1125=>x"3000", 1126=>x"2500", 1127=>x"4200",
---- 1128=>x"6000", 1129=>x"4d00", 1130=>x"2c00", 1131=>x"2700", 1132=>x"3000", 1133=>x"3400", 1134=>x"2c00",
---- 1135=>x"3300", 1136=>x"5300", 1137=>x"3c00", 1138=>x"2b00", 1139=>x"2600", 1140=>x"4400", 1141=>x"4000",
---- 1142=>x"3800", 1143=>x"4400", 1144=>x"3300", 1145=>x"3700", 1146=>x"2c00", 1147=>x"2f00", 1148=>x"af00",
---- 1149=>x"4700", 1150=>x"4f00", 1151=>x"6c00", 1152=>x"3600", 1153=>x"c900", 1154=>x"cd00", 1155=>x"3900",
---- 1156=>x"6400", 1157=>x"5100", 1158=>x"6700", 1159=>x"7600", 1160=>x"3b00", 1161=>x"4500", 1162=>x"4000",
---- 1163=>x"4400", 1164=>x"6c00", 1165=>x"4c00", 1166=>x"6900", 1167=>x"7600", 1168=>x"3e00", 1169=>x"4200",
---- 1170=>x"3c00", 1171=>x"5100", 1172=>x"6500", 1173=>x"4c00", 1174=>x"6e00", 1175=>x"5a00", 1176=>x"3f00",
---- 1177=>x"3900", 1178=>x"4b00", 1179=>x"5c00", 1180=>x"4f00", 1181=>x"6100", 1182=>x"7000", 1183=>x"7100",
---- 1184=>x"3c00", 1185=>x"5000", 1186=>x"6f00", 1187=>x"4900", 1188=>x"4200", 1189=>x"7200", 1190=>x"8200",
---- 1191=>x"8700", 1192=>x"5700", 1193=>x"7500", 1194=>x"5a00", 1195=>x"3300", 1196=>x"4b00", 1197=>x"8800",
---- 1198=>x"7900", 1199=>x"6500", 1200=>x"7400", 1201=>x"5500", 1202=>x"3000", 1203=>x"3400", 1204=>x"4700",
---- 1205=>x"7500", 1206=>x"7f00", 1207=>x"6000", 1208=>x"4e00", 1209=>x"3200", 1210=>x"3d00", 1211=>x"3d00",
---- 1212=>x"3000", 1213=>x"4a00", 1214=>x"8700", 1215=>x"6200", 1216=>x"2d00", 1217=>x"4c00", 1218=>x"5100",
---- 1219=>x"4800", 1220=>x"3800", 1221=>x"4d00", 1222=>x"8800", 1223=>x"6d00", 1224=>x"2e00", 1225=>x"6800",
---- 1226=>x"5700", 1227=>x"4900", 1228=>x"3900", 1229=>x"8100", 1230=>x"7300", 1231=>x"7700", 1232=>x"4500",
---- 1233=>x"6600", 1234=>x"6300", 1235=>x"6200", 1236=>x"4b00", 1237=>x"8b00", 1238=>x"7000", 1239=>x"7e00",
---- 1240=>x"6400", 1241=>x"5100", 1242=>x"7500", 1243=>x"5200", 1244=>x"5a00", 1245=>x"8000", 1246=>x"6800",
---- 1247=>x"8f00", 1248=>x"5100", 1249=>x"6500", 1250=>x"7900", 1251=>x"4d00", 1252=>x"5f00", 1253=>x"6a00",
---- 1254=>x"6800", 1255=>x"9b00", 1256=>x"3f00", 1257=>x"7900", 1258=>x"5800", 1259=>x"3f00", 1260=>x"6000",
---- 1261=>x"5900", 1262=>x"6200", 1263=>x"9c00", 1264=>x"5400", 1265=>x"8400", 1266=>x"3700", 1267=>x"3400",
---- 1268=>x"7200", 1269=>x"5900", 1270=>x"5a00", 1271=>x"9800", 1272=>x"6f00", 1273=>x"6e00", 1274=>x"2e00",
---- 1275=>x"3500", 1276=>x"8500", 1277=>x"6500", 1278=>x"4b00", 1279=>x"9500", 1280=>x"7e00", 1281=>x"5300",
---- 1282=>x"3300", 1283=>x"2c00", 1284=>x"6a00", 1285=>x"6c00", 1286=>x"3f00", 1287=>x"8100", 1288=>x"7a00",
---- 1289=>x"4800", 1290=>x"4300", 1291=>x"2b00", 1292=>x"5a00", 1293=>x"8c00", 1294=>x"5100", 1295=>x"7300",
---- 1296=>x"5100", 1297=>x"3d00", 1298=>x"5c00", 1299=>x"3500", 1300=>x"5500", 1301=>x"6d00", 1302=>x"5900",
---- 1303=>x"6f00", 1304=>x"4100", 1305=>x"4a00", 1306=>x"6b00", 1307=>x"3500", 1308=>x"4d00", 1309=>x"7900",
---- 1310=>x"5c00", 1311=>x"6c00", 1312=>x"4f00", 1313=>x"5400", 1314=>x"5500", 1315=>x"3d00", 1316=>x"4900",
---- 1317=>x"7e00", 1318=>x"5300", 1319=>x"6300", 1320=>x"5000", 1321=>x"5300", 1322=>x"4500", 1323=>x"5900",
---- 1324=>x"5100", 1325=>x"7200", 1326=>x"5500", 1327=>x"7400", 1328=>x"4b00", 1329=>x"4d00", 1330=>x"4400",
---- 1331=>x"6300", 1332=>x"6b00", 1333=>x"7000", 1334=>x"6800", 1335=>x"7900", 1336=>x"4400", 1337=>x"4d00",
---- 1338=>x"4400", 1339=>x"4d00", 1340=>x"6700", 1341=>x"6100", 1342=>x"6700", 1343=>x"7a00", 1344=>x"4100",
---- 1345=>x"4600", 1346=>x"4800", 1347=>x"4300", 1348=>x"5900", 1349=>x"4800", 1350=>x"5b00", 1351=>x"6f00",
---- 1352=>x"4400", 1353=>x"4300", 1354=>x"4d00", 1355=>x"3e00", 1356=>x"5100", 1357=>x"4800", 1358=>x"5900",
---- 1359=>x"7000", 1360=>x"4700", 1361=>x"3800", 1362=>x"5200", 1363=>x"4600", 1364=>x"4500", 1365=>x"4a00",
---- 1366=>x"4500", 1367=>x"7000", 1368=>x"4600", 1369=>x"3b00", 1370=>x"4a00", 1371=>x"5400", 1372=>x"4100",
---- 1373=>x"4500", 1374=>x"4100", 1375=>x"5d00", 1376=>x"3f00", 1377=>x"5400", 1378=>x"5300", 1379=>x"5300",
---- 1380=>x"4a00", 1381=>x"4000", 1382=>x"4a00", 1383=>x"b100", 1384=>x"4300", 1385=>x"4d00", 1386=>x"6a00",
---- 1387=>x"5600", 1388=>x"6000", 1389=>x"5400", 1390=>x"4f00", 1391=>x"4f00", 1392=>x"3900", 1393=>x"4600",
---- 1394=>x"7800", 1395=>x"5f00", 1396=>x"6400", 1397=>x"6600", 1398=>x"5700", 1399=>x"4b00", 1400=>x"3300",
---- 1401=>x"4e00", 1402=>x"8800", 1403=>x"7700", 1404=>x"6700", 1405=>x"6300", 1406=>x"6900", 1407=>x"5a00",
---- 1408=>x"3500", 1409=>x"4d00", 1410=>x"8800", 1411=>x"7f00", 1412=>x"6700", 1413=>x"5e00", 1414=>x"6600",
---- 1415=>x"6500", 1416=>x"3400", 1417=>x"4a00", 1418=>x"6300", 1419=>x"8600", 1420=>x"5500", 1421=>x"5b00",
---- 1422=>x"6200", 1423=>x"5f00", 1424=>x"3700", 1425=>x"4b00", 1426=>x"aa00", 1427=>x"8400", 1428=>x"4a00",
---- 1429=>x"3d00", 1430=>x"5c00", 1431=>x"6d00", 1432=>x"4500", 1433=>x"5000", 1434=>x"ac00", 1435=>x"8500",
---- 1436=>x"4f00", 1437=>x"3200", 1438=>x"5100", 1439=>x"5a00", 1440=>x"5400", 1441=>x"6b00", 1442=>x"a700",
---- 1443=>x"7900", 1444=>x"8800", 1445=>x"3c00", 1446=>x"4800", 1447=>x"5800", 1448=>x"4e00", 1449=>x"8800",
---- 1450=>x"6800", 1451=>x"5e00", 1452=>x"8100", 1453=>x"9a00", 1454=>x"4c00", 1455=>x"7000", 1456=>x"5200",
---- 1457=>x"9b00", 1458=>x"9900", 1459=>x"5500", 1460=>x"5b00", 1461=>x"8600", 1462=>x"6600", 1463=>x"7d00",
---- 1464=>x"6200", 1465=>x"ad00", 1466=>x"9a00", 1467=>x"6700", 1468=>x"3e00", 1469=>x"8800", 1470=>x"7900",
---- 1471=>x"7b00", 1472=>x"7000", 1473=>x"ad00", 1474=>x"8500", 1475=>x"8d00", 1476=>x"5400", 1477=>x"6700",
---- 1478=>x"9000", 1479=>x"8000", 1480=>x"6d00", 1481=>x"ab00", 1482=>x"8200", 1483=>x"7100", 1484=>x"7b00",
---- 1485=>x"5e00", 1486=>x"9300", 1487=>x"8b00", 1488=>x"5200", 1489=>x"9700", 1490=>x"6c00", 1491=>x"6500",
---- 1492=>x"7500", 1493=>x"6d00", 1494=>x"7600", 1495=>x"9500", 1496=>x"5300", 1497=>x"8f00", 1498=>x"6000",
---- 1499=>x"5e00", 1500=>x"6d00", 1501=>x"7700", 1502=>x"6e00", 1503=>x"8400", 1504=>x"5b00", 1505=>x"7e00",
---- 1506=>x"6700", 1507=>x"4e00", 1508=>x"3e00", 1509=>x"5200", 1510=>x"7300", 1511=>x"7b00", 1512=>x"6600",
---- 1513=>x"8300", 1514=>x"6300", 1515=>x"4900", 1516=>x"3200", 1517=>x"3600", 1518=>x"4600", 1519=>x"6e00",
---- 1520=>x"6600", 1521=>x"8a00", 1522=>x"7e00", 1523=>x"5c00", 1524=>x"2f00", 1525=>x"4200", 1526=>x"4300",
---- 1527=>x"a400", 1528=>x"5300", 1529=>x"9200", 1530=>x"8100", 1531=>x"7100", 1532=>x"3600", 1533=>x"4800",
---- 1534=>x"5000", 1535=>x"5a00", 1536=>x"4000", 1537=>x"9900", 1538=>x"8400", 1539=>x"7d00", 1540=>x"4000",
---- 1541=>x"4300", 1542=>x"5200", 1543=>x"4400", 1544=>x"3700", 1545=>x"9000", 1546=>x"9000", 1547=>x"9000",
---- 1548=>x"5f00", 1549=>x"5600", 1550=>x"5f00", 1551=>x"3f00", 1552=>x"3400", 1553=>x"8500", 1554=>x"8300",
---- 1555=>x"9200", 1556=>x"8900", 1557=>x"5800", 1558=>x"5700", 1559=>x"4300", 1560=>x"4000", 1561=>x"8500",
---- 1562=>x"7800", 1563=>x"7b00", 1564=>x"9300", 1565=>x"5f00", 1566=>x"4c00", 1567=>x"4e00", 1568=>x"4200",
---- 1569=>x"7e00", 1570=>x"8200", 1571=>x"6f00", 1572=>x"8100", 1573=>x"9400", 1574=>x"5f00", 1575=>x"3f00",
---- 1576=>x"3800", 1577=>x"5600", 1578=>x"7b00", 1579=>x"8300", 1580=>x"6c00", 1581=>x"7f00", 1582=>x"8b00",
---- 1583=>x"5100", 1584=>x"3a00", 1585=>x"3500", 1586=>x"4a00", 1587=>x"8700", 1588=>x"7b00", 1589=>x"ab00",
---- 1590=>x"7e00", 1591=>x"8400", 1592=>x"4a00", 1593=>x"3200", 1594=>x"2100", 1595=>x"6b00", 1596=>x"8e00",
---- 1597=>x"6e00", 1598=>x"5500", 1599=>x"4500", 1600=>x"5d00", 1601=>x"2d00", 1602=>x"1f00", 1603=>x"3800",
---- 1604=>x"7400", 1605=>x"8b00", 1606=>x"7800", 1607=>x"5000", 1608=>x"6a00", 1609=>x"2e00", 1610=>x"2900",
---- 1611=>x"2500", 1612=>x"4000", 1613=>x"7600", 1614=>x"8300", 1615=>x"8a00", 1616=>x"4900", 1617=>x"3300",
---- 1618=>x"2c00", 1619=>x"2e00", 1620=>x"5b00", 1621=>x"5300", 1622=>x"3c00", 1623=>x"6000", 1624=>x"4c00",
---- 1625=>x"3200", 1626=>x"2a00", 1627=>x"6000", 1628=>x"6f00", 1629=>x"4200", 1630=>x"3800", 1631=>x"5200",
---- 1632=>x"4800", 1633=>x"4300", 1634=>x"6700", 1635=>x"8000", 1636=>x"4500", 1637=>x"2c00", 1638=>x"3a00",
---- 1639=>x"7a00", 1640=>x"a500", 1641=>x"6700", 1642=>x"6600", 1643=>x"4c00", 1644=>x"2900", 1645=>x"2000",
---- 1646=>x"5400", 1647=>x"9200", 1648=>x"3a00", 1649=>x"3100", 1650=>x"2f00", 1651=>x"3500", 1652=>x"2e00",
---- 1653=>x"2b00", 1654=>x"9e00", 1655=>x"8b00", 1656=>x"2d00", 1657=>x"2800", 1658=>x"2a00", 1659=>x"4000",
---- 1660=>x"4000", 1661=>x"2900", 1662=>x"3900", 1663=>x"5700", 1664=>x"3500", 1665=>x"2800", 1666=>x"2800",
---- 1667=>x"4500", 1668=>x"5b00", 1669=>x"2700", 1670=>x"2700", 1671=>x"3e00", 1672=>x"4800", 1673=>x"2900",
---- 1674=>x"2700", 1675=>x"3700", 1676=>x"6a00", 1677=>x"3800", 1678=>x"2700", 1679=>x"3800", 1680=>x"4900",
---- 1681=>x"2a00", 1682=>x"2500", 1683=>x"2700", 1684=>x"5f00", 1685=>x"5800", 1686=>x"2700", 1687=>x"2d00",
---- 1688=>x"4600", 1689=>x"3200", 1690=>x"2600", 1691=>x"2300", 1692=>x"3600", 1693=>x"5c00", 1694=>x"4b00",
---- 1695=>x"2600", 1696=>x"5200", 1697=>x"3a00", 1698=>x"2400", 1699=>x"2600", 1700=>x"2700", 1701=>x"3100",
---- 1702=>x"6000", 1703=>x"5100", 1704=>x"5200", 1705=>x"3800", 1706=>x"2400", 1707=>x"2700", 1708=>x"3300",
---- 1709=>x"2900", 1710=>x"3e00", 1711=>x"5800", 1712=>x"4b00", 1713=>x"4700", 1714=>x"2600", 1715=>x"2e00",
---- 1716=>x"3b00", 1717=>x"2b00", 1718=>x"3800", 1719=>x"3600", 1720=>x"3e00", 1721=>x"4d00", 1722=>x"2800",
---- 1723=>x"3500", 1724=>x"4200", 1725=>x"2d00", 1726=>x"3f00", 1727=>x"3a00", 1728=>x"3000", 1729=>x"3f00",
---- 1730=>x"2900", 1731=>x"3e00", 1732=>x"4400", 1733=>x"3000", 1734=>x"3600", 1735=>x"3b00", 1736=>x"2b00",
---- 1737=>x"3700", 1738=>x"3000", 1739=>x"4100", 1740=>x"3b00", 1741=>x"3600", 1742=>x"2e00", 1743=>x"3200",
---- 1744=>x"2900", 1745=>x"2e00", 1746=>x"3a00", 1747=>x"4500", 1748=>x"2f00", 1749=>x"3500", 1750=>x"2700",
---- 1751=>x"2700", 1752=>x"2e00", 1753=>x"3200", 1754=>x"4500", 1755=>x"4a00", 1756=>x"2a00", 1757=>x"3500",
---- 1758=>x"2d00", 1759=>x"2600", 1760=>x"2d00", 1761=>x"3300", 1762=>x"4f00", 1763=>x"4300", 1764=>x"2d00",
---- 1765=>x"2d00", 1766=>x"3000", 1767=>x"2700", 1768=>x"2800", 1769=>x"3600", 1770=>x"4600", 1771=>x"3a00",
---- 1772=>x"3500", 1773=>x"2900", 1774=>x"2e00", 1775=>x"2a00", 1776=>x"3400", 1777=>x"3e00", 1778=>x"2f00",
---- 1779=>x"3700", 1780=>x"3800", 1781=>x"2e00", 1782=>x"3300", 1783=>x"3100", 1784=>x"3c00", 1785=>x"3d00",
---- 1786=>x"2c00", 1787=>x"3500", 1788=>x"3d00", 1789=>x"3000", 1790=>x"3200", 1791=>x"2c00", 1792=>x"3a00",
---- 1793=>x"3000", 1794=>x"2f00", 1795=>x"3c00", 1796=>x"4500", 1797=>x"2e00", 1798=>x"2a00", 1799=>x"2600",
---- 1800=>x"2b00", 1801=>x"2d00", 1802=>x"2e00", 1803=>x"3500", 1804=>x"4c00", 1805=>x"3700", 1806=>x"2500",
---- 1807=>x"2b00", 1808=>x"3000", 1809=>x"3200", 1810=>x"3300", 1811=>x"2f00", 1812=>x"4100", 1813=>x"3d00",
---- 1814=>x"2500", 1815=>x"2b00", 1816=>x"c600", 1817=>x"3800", 1818=>x"3800", 1819=>x"2f00", 1820=>x"3500",
---- 1821=>x"5100", 1822=>x"2a00", 1823=>x"3200", 1824=>x"3f00", 1825=>x"4500", 1826=>x"4100", 1827=>x"3300",
---- 1828=>x"2900", 1829=>x"4200", 1830=>x"3c00", 1831=>x"3c00", 1832=>x"3f00", 1833=>x"3a00", 1834=>x"3d00",
---- 1835=>x"3b00", 1836=>x"3500", 1837=>x"4000", 1838=>x"3e00", 1839=>x"2e00", 1840=>x"4500", 1841=>x"3000",
---- 1842=>x"3100", 1843=>x"3200", 1844=>x"3c00", 1845=>x"3700", 1846=>x"2c00", 1847=>x"2700", 1848=>x"4900",
---- 1849=>x"2f00", 1850=>x"2a00", 1851=>x"2b00", 1852=>x"3100", 1853=>x"3400", 1854=>x"2f00", 1855=>x"2900",
---- 1856=>x"4900", 1857=>x"3500", 1858=>x"3000", 1859=>x"2c00", 1860=>x"2e00", 1861=>x"2b00", 1862=>x"3100",
---- 1863=>x"2800", 1864=>x"4300", 1865=>x"3700", 1866=>x"3400", 1867=>x"2f00", 1868=>x"2b00", 1869=>x"2b00",
---- 1870=>x"3200", 1871=>x"3300", 1872=>x"4200", 1873=>x"3900", 1874=>x"3d00", 1875=>x"3900", 1876=>x"2a00",
---- 1877=>x"2b00", 1878=>x"3100", 1879=>x"3500", 1880=>x"4300", 1881=>x"4000", 1882=>x"4100", 1883=>x"3a00",
---- 1884=>x"3200", 1885=>x"2800", 1886=>x"3500", 1887=>x"3200", 1888=>x"3b00", 1889=>x"3b00", 1890=>x"3900",
---- 1891=>x"3600", 1892=>x"3a00", 1893=>x"3700", 1894=>x"3400", 1895=>x"2e00", 1896=>x"3b00", 1897=>x"3a00",
---- 1898=>x"3a00", 1899=>x"3800", 1900=>x"3400", 1901=>x"3c00", 1902=>x"2d00", 1903=>x"2a00", 1904=>x"4200",
---- 1905=>x"3600", 1906=>x"3f00", 1907=>x"3d00", 1908=>x"3100", 1909=>x"2f00", 1910=>x"2a00", 1911=>x"2c00",
---- 1912=>x"4700", 1913=>x"3c00", 1914=>x"4000", 1915=>x"3e00", 1916=>x"2d00", 1917=>x"2f00", 1918=>x"2f00",
---- 1919=>x"2a00", 1920=>x"4800", 1921=>x"3b00", 1922=>x"3a00", 1923=>x"3a00", 1924=>x"3b00", 1925=>x"2e00",
---- 1926=>x"2c00", 1927=>x"2c00", 1928=>x"4200", 1929=>x"3500", 1930=>x"3000", 1931=>x"3f00", 1932=>x"5400",
---- 1933=>x"3700", 1934=>x"3100", 1935=>x"3100", 1936=>x"4500", 1937=>x"3100", 1938=>x"3000", 1939=>x"4b00",
---- 1940=>x"5b00", 1941=>x"3900", 1942=>x"2a00", 1943=>x"3400", 1944=>x"5400", 1945=>x"3000", 1946=>x"3800",
---- 1947=>x"4b00", 1948=>x"5b00", 1949=>x"4d00", 1950=>x"2a00", 1951=>x"2e00", 1952=>x"6300", 1953=>x"2f00",
---- 1954=>x"c900", 1955=>x"5100", 1956=>x"5f00", 1957=>x"5800", 1958=>x"3d00", 1959=>x"2600", 1960=>x"6200",
---- 1961=>x"2900", 1962=>x"3500", 1963=>x"5000", 1964=>x"6500", 1965=>x"6100", 1966=>x"5b00", 1967=>x"3200",
---- 1968=>x"5600", 1969=>x"2800", 1970=>x"3500", 1971=>x"5600", 1972=>x"6c00", 1973=>x"7300", 1974=>x"6b00",
---- 1975=>x"4a00", 1976=>x"4c00", 1977=>x"2700", 1978=>x"2e00", 1979=>x"5100", 1980=>x"6900", 1981=>x"7000",
---- 1982=>x"6c00", 1983=>x"5200", 1984=>x"3a00", 1985=>x"2a00", 1986=>x"2900", 1987=>x"4800", 1988=>x"6500",
---- 1989=>x"5d00", 1990=>x"7f00", 1991=>x"9e00", 1992=>x"2a00", 1993=>x"2c00", 1994=>x"2700", 1995=>x"4400",
---- 1996=>x"7000", 1997=>x"4700", 1998=>x"7000", 1999=>x"8000", 2000=>x"2f00", 2001=>x"2c00", 2002=>x"2b00",
---- 2003=>x"4200", 2004=>x"7700", 2005=>x"4600", 2006=>x"5100", 2007=>x"8e00", 2008=>x"2d00", 2009=>x"3000",
---- 2010=>x"2f00", 2011=>x"4700", 2012=>x"7900", 2013=>x"5000", 2014=>x"4200", 2015=>x"8800", 2016=>x"3100",
---- 2017=>x"2f00", 2018=>x"2c00", 2019=>x"5000", 2020=>x"7e00", 2021=>x"4c00", 2022=>x"4600", 2023=>x"6700",
---- 2024=>x"3a00", 2025=>x"2e00", 2026=>x"3700", 2027=>x"5300", 2028=>x"7700", 2029=>x"3d00", 2030=>x"4c00",
---- 2031=>x"4a00", 2032=>x"3d00", 2033=>x"3400", 2034=>x"3c00", 2035=>x"4f00", 2036=>x"7d00", 2037=>x"3800",
---- 2038=>x"4300", 2039=>x"5300", 2040=>x"4500", 2041=>x"3200", 2042=>x"3600", 2043=>x"4e00", 2044=>x"7a00",
---- 2045=>x"3b00", 2046=>x"3300", 2047=>x"5300"),
---- 8  => (0=>x"7c00", 1=>x"8300", 2=>x"8000", 3=>x"8100", 4=>x"8500", 5=>x"8600", 6=>x"8300", 7=>x"8000",
---- 8=>x"8300", 9=>x"8300", 10=>x"8100", 11=>x"8100", 12=>x"8500", 13=>x"8600", 14=>x"8400",
---- 15=>x"8100", 16=>x"8200", 17=>x"8300", 18=>x"8200", 19=>x"8100", 20=>x"8400", 21=>x"8500",
---- 22=>x"8400", 23=>x"8200", 24=>x"7c00", 25=>x"8100", 26=>x"8400", 27=>x"8000", 28=>x"8100",
---- 29=>x"8200", 30=>x"8400", 31=>x"8100", 32=>x"7e00", 33=>x"8000", 34=>x"8000", 35=>x"8200",
---- 36=>x"8300", 37=>x"8200", 38=>x"8200", 39=>x"8200", 40=>x"7f00", 41=>x"8300", 42=>x"7f00",
---- 43=>x"8000", 44=>x"8100", 45=>x"8100", 46=>x"8000", 47=>x"8300", 48=>x"7e00", 49=>x"7e00",
---- 50=>x"7f00", 51=>x"8300", 52=>x"7e00", 53=>x"8200", 54=>x"8100", 55=>x"8400", 56=>x"7e00",
---- 57=>x"7d00", 58=>x"8000", 59=>x"8000", 60=>x"7d00", 61=>x"8300", 62=>x"8300", 63=>x"8300",
---- 64=>x"7f00", 65=>x"8100", 66=>x"7f00", 67=>x"8300", 68=>x"7f00", 69=>x"8200", 70=>x"8200",
---- 71=>x"8200", 72=>x"8000", 73=>x"8000", 74=>x"8000", 75=>x"8200", 76=>x"8100", 77=>x"8100",
---- 78=>x"8500", 79=>x"8400", 80=>x"7d00", 81=>x"7f00", 82=>x"8000", 83=>x"8100", 84=>x"8100",
---- 85=>x"8100", 86=>x"8300", 87=>x"8100", 88=>x"7c00", 89=>x"8000", 90=>x"8000", 91=>x"8200",
---- 92=>x"8200", 93=>x"8000", 94=>x"8300", 95=>x"8100", 96=>x"8000", 97=>x"8300", 98=>x"7f00",
---- 99=>x"7e00", 100=>x"8000", 101=>x"8300", 102=>x"8100", 103=>x"8200", 104=>x"7f00", 105=>x"8100",
---- 106=>x"8000", 107=>x"7d00", 108=>x"7f00", 109=>x"8100", 110=>x"8100", 111=>x"8200", 112=>x"8000",
---- 113=>x"7e00", 114=>x"7d00", 115=>x"7e00", 116=>x"8100", 117=>x"7e00", 118=>x"7e00", 119=>x"8100",
---- 120=>x"7e00", 121=>x"7e00", 122=>x"8000", 123=>x"7f00", 124=>x"7f00", 125=>x"8000", 126=>x"7f00",
---- 127=>x"7e00", 128=>x"7e00", 129=>x"7e00", 130=>x"8100", 131=>x"7d00", 132=>x"7e00", 133=>x"8100",
---- 134=>x"8000", 135=>x"7f00", 136=>x"7d00", 137=>x"7d00", 138=>x"7f00", 139=>x"8100", 140=>x"8000",
---- 141=>x"7f00", 142=>x"8000", 143=>x"8200", 144=>x"7a00", 145=>x"7c00", 146=>x"7f00", 147=>x"8000",
---- 148=>x"7f00", 149=>x"7d00", 150=>x"8200", 151=>x"8100", 152=>x"7c00", 153=>x"7d00", 154=>x"7e00",
---- 155=>x"7e00", 156=>x"7b00", 157=>x"7b00", 158=>x"8100", 159=>x"8100", 160=>x"7c00", 161=>x"7a00",
---- 162=>x"7900", 163=>x"7e00", 164=>x"7e00", 165=>x"7d00", 166=>x"7d00", 167=>x"7e00", 168=>x"7c00",
---- 169=>x"7d00", 170=>x"7800", 171=>x"7c00", 172=>x"7c00", 173=>x"8000", 174=>x"7e00", 175=>x"7a00",
---- 176=>x"7d00", 177=>x"7d00", 178=>x"7c00", 179=>x"7b00", 180=>x"8200", 181=>x"7e00", 182=>x"7d00",
---- 183=>x"7c00", 184=>x"7b00", 185=>x"7c00", 186=>x"7b00", 187=>x"7e00", 188=>x"7e00", 189=>x"7f00",
---- 190=>x"7d00", 191=>x"7b00", 192=>x"7b00", 193=>x"7d00", 194=>x"7c00", 195=>x"7f00", 196=>x"7f00",
---- 197=>x"7f00", 198=>x"8000", 199=>x"7f00", 200=>x"7f00", 201=>x"7c00", 202=>x"8400", 203=>x"7e00",
---- 204=>x"7d00", 205=>x"7e00", 206=>x"7d00", 207=>x"7f00", 208=>x"7f00", 209=>x"8000", 210=>x"7d00",
---- 211=>x"7d00", 212=>x"7b00", 213=>x"7d00", 214=>x"7d00", 215=>x"7d00", 216=>x"8200", 217=>x"7e00",
---- 218=>x"7f00", 219=>x"7c00", 220=>x"7c00", 221=>x"7c00", 222=>x"8000", 223=>x"8100", 224=>x"7f00",
---- 225=>x"7c00", 226=>x"7c00", 227=>x"7d00", 228=>x"7e00", 229=>x"7d00", 230=>x"8000", 231=>x"8000",
---- 232=>x"7c00", 233=>x"7900", 234=>x"7a00", 235=>x"7b00", 236=>x"7700", 237=>x"7e00", 238=>x"7e00",
---- 239=>x"7b00", 240=>x"7800", 241=>x"7a00", 242=>x"7d00", 243=>x"7a00", 244=>x"7b00", 245=>x"7900",
---- 246=>x"7e00", 247=>x"7e00", 248=>x"7a00", 249=>x"7a00", 250=>x"7d00", 251=>x"7b00", 252=>x"8300",
---- 253=>x"7c00", 254=>x"7c00", 255=>x"7d00", 256=>x"7b00", 257=>x"7900", 258=>x"7b00", 259=>x"7b00",
---- 260=>x"7800", 261=>x"7a00", 262=>x"7c00", 263=>x"7e00", 264=>x"7c00", 265=>x"7c00", 266=>x"7a00",
---- 267=>x"7c00", 268=>x"7b00", 269=>x"7b00", 270=>x"7c00", 271=>x"7c00", 272=>x"7900", 273=>x"7c00",
---- 274=>x"7800", 275=>x"7900", 276=>x"7a00", 277=>x"7d00", 278=>x"7a00", 279=>x"7b00", 280=>x"7600",
---- 281=>x"7700", 282=>x"7700", 283=>x"7700", 284=>x"7b00", 285=>x"7b00", 286=>x"7a00", 287=>x"7e00",
---- 288=>x"7700", 289=>x"7700", 290=>x"7500", 291=>x"7800", 292=>x"7900", 293=>x"7600", 294=>x"7b00",
---- 295=>x"7b00", 296=>x"7900", 297=>x"7900", 298=>x"7700", 299=>x"7700", 300=>x"7900", 301=>x"8500",
---- 302=>x"7a00", 303=>x"7c00", 304=>x"8800", 305=>x"7500", 306=>x"7700", 307=>x"7600", 308=>x"7800",
---- 309=>x"7b00", 310=>x"7800", 311=>x"7900", 312=>x"7800", 313=>x"7900", 314=>x"7800", 315=>x"7800",
---- 316=>x"7c00", 317=>x"7a00", 318=>x"7900", 319=>x"7900", 320=>x"7b00", 321=>x"7900", 322=>x"7d00",
---- 323=>x"7900", 324=>x"7b00", 325=>x"7d00", 326=>x"7600", 327=>x"7700", 328=>x"7900", 329=>x"7600",
---- 330=>x"7a00", 331=>x"7a00", 332=>x"7a00", 333=>x"7700", 334=>x"7900", 335=>x"7b00", 336=>x"7900",
---- 337=>x"7900", 338=>x"7900", 339=>x"7800", 340=>x"7c00", 341=>x"7900", 342=>x"7d00", 343=>x"7b00",
---- 344=>x"7800", 345=>x"7800", 346=>x"7800", 347=>x"7800", 348=>x"7b00", 349=>x"7a00", 350=>x"7e00",
---- 351=>x"7b00", 352=>x"7900", 353=>x"7700", 354=>x"7900", 355=>x"7900", 356=>x"7a00", 357=>x"7b00",
---- 358=>x"7b00", 359=>x"8100", 360=>x"7a00", 361=>x"7a00", 362=>x"7800", 363=>x"7c00", 364=>x"7800",
---- 365=>x"7700", 366=>x"8100", 367=>x"8100", 368=>x"7900", 369=>x"7c00", 370=>x"7800", 371=>x"7800",
---- 372=>x"8400", 373=>x"7b00", 374=>x"7f00", 375=>x"7200", 376=>x"7600", 377=>x"7800", 378=>x"7b00",
---- 379=>x"7c00", 380=>x"7b00", 381=>x"7f00", 382=>x"7900", 383=>x"7000", 384=>x"7700", 385=>x"7700",
---- 386=>x"7800", 387=>x"7a00", 388=>x"7f00", 389=>x"7e00", 390=>x"7400", 391=>x"7500", 392=>x"8500",
---- 393=>x"7900", 394=>x"7800", 395=>x"7a00", 396=>x"8900", 397=>x"7800", 398=>x"6f00", 399=>x"7100",
---- 400=>x"7b00", 401=>x"7700", 402=>x"7800", 403=>x"8500", 404=>x"8900", 405=>x"6f00", 406=>x"6b00",
---- 407=>x"6c00", 408=>x"7900", 409=>x"7600", 410=>x"7a00", 411=>x"8900", 412=>x"7b00", 413=>x"6d00",
---- 414=>x"6e00", 415=>x"6900", 416=>x"7300", 417=>x"7400", 418=>x"9400", 419=>x"8500", 420=>x"6d00",
---- 421=>x"6900", 422=>x"6700", 423=>x"6500", 424=>x"6f00", 425=>x"8700", 426=>x"b600", 427=>x"7b00",
---- 428=>x"6400", 429=>x"6500", 430=>x"6800", 431=>x"6700", 432=>x"6c00", 433=>x"9f00", 434=>x"b300",
---- 435=>x"7400", 436=>x"5f00", 437=>x"6700", 438=>x"6b00", 439=>x"6c00", 440=>x"7400", 441=>x"c000",
---- 442=>x"a900", 443=>x"6900", 444=>x"6200", 445=>x"6700", 446=>x"6d00", 447=>x"6900", 448=>x"9800",
---- 449=>x"cf00", 450=>x"9400", 451=>x"6400", 452=>x"6600", 453=>x"6900", 454=>x"6700", 455=>x"6900",
---- 456=>x"be00", 457=>x"c700", 458=>x"8a00", 459=>x"6100", 460=>x"6600", 461=>x"6b00", 462=>x"6700",
---- 463=>x"6700", 464=>x"d600", 465=>x"b600", 466=>x"7a00", 467=>x"6000", 468=>x"6700", 469=>x"6800",
---- 470=>x"6600", 471=>x"6a00", 472=>x"d900", 473=>x"a000", 474=>x"7b00", 475=>x"6600", 476=>x"6300",
---- 477=>x"6700", 478=>x"6700", 479=>x"6a00", 480=>x"c800", 481=>x"a700", 482=>x"8400", 483=>x"6700",
---- 484=>x"6100", 485=>x"6800", 486=>x"6800", 487=>x"6a00", 488=>x"c300", 489=>x"a200", 490=>x"7a00",
---- 491=>x"6600", 492=>x"9a00", 493=>x"6200", 494=>x"6400", 495=>x"6a00", 496=>x"be00", 497=>x"9600",
---- 498=>x"7300", 499=>x"6000", 500=>x"6100", 501=>x"6600", 502=>x"6900", 503=>x"6800", 504=>x"b800",
---- 505=>x"9600", 506=>x"6e00", 507=>x"5c00", 508=>x"6000", 509=>x"6700", 510=>x"6600", 511=>x"6800",
---- 512=>x"b100", 513=>x"5e00", 514=>x"7200", 515=>x"5b00", 516=>x"6400", 517=>x"6700", 518=>x"6600",
---- 519=>x"6d00", 520=>x"b100", 521=>x"8d00", 522=>x"7100", 523=>x"6200", 524=>x"6800", 525=>x"6700",
---- 526=>x"6700", 527=>x"6b00", 528=>x"a800", 529=>x"8300", 530=>x"6f00", 531=>x"6200", 532=>x"6100",
---- 533=>x"6200", 534=>x"6500", 535=>x"6700", 536=>x"9b00", 537=>x"7b00", 538=>x"7000", 539=>x"6400",
---- 540=>x"5d00", 541=>x"6100", 542=>x"6400", 543=>x"9a00", 544=>x"9300", 545=>x"7400", 546=>x"7500",
---- 547=>x"6a00", 548=>x"5f00", 549=>x"6000", 550=>x"6400", 551=>x"6b00", 552=>x"8900", 553=>x"8300",
---- 554=>x"7800", 555=>x"6c00", 556=>x"6400", 557=>x"6400", 558=>x"6800", 559=>x"6c00", 560=>x"9200",
---- 561=>x"8200", 562=>x"7c00", 563=>x"6c00", 564=>x"6900", 565=>x"6800", 566=>x"6900", 567=>x"6700",
---- 568=>x"9200", 569=>x"8200", 570=>x"7e00", 571=>x"6b00", 572=>x"6600", 573=>x"6d00", 574=>x"6800",
---- 575=>x"6900", 576=>x"9e00", 577=>x"8600", 578=>x"7f00", 579=>x"7100", 580=>x"9800", 581=>x"6800",
---- 582=>x"6200", 583=>x"6b00", 584=>x"9d00", 585=>x"8b00", 586=>x"8000", 587=>x"7400", 588=>x"6a00",
---- 589=>x"6300", 590=>x"6c00", 591=>x"6d00", 592=>x"9d00", 593=>x"9100", 594=>x"7a00", 595=>x"7700",
---- 596=>x"7000", 597=>x"7000", 598=>x"6f00", 599=>x"6900", 600=>x"9f00", 601=>x"9400", 602=>x"8a00",
---- 603=>x"8200", 604=>x"7b00", 605=>x"7e00", 606=>x"6f00", 607=>x"6e00", 608=>x"9900", 609=>x"9000",
---- 610=>x"8b00", 611=>x"8800", 612=>x"7a00", 613=>x"8000", 614=>x"7700", 615=>x"7300", 616=>x"a000",
---- 617=>x"9d00", 618=>x"8800", 619=>x"9000", 620=>x"8100", 621=>x"8300", 622=>x"8100", 623=>x"6c00",
---- 624=>x"aa00", 625=>x"a400", 626=>x"9a00", 627=>x"8b00", 628=>x"9300", 629=>x"8200", 630=>x"7e00",
---- 631=>x"6f00", 632=>x"9c00", 633=>x"a000", 634=>x"9500", 635=>x"8f00", 636=>x"8d00", 637=>x"8800",
---- 638=>x"8400", 639=>x"7f00", 640=>x"a900", 641=>x"9c00", 642=>x"ad00", 643=>x"9200", 644=>x"8e00",
---- 645=>x"8700", 646=>x"8e00", 647=>x"8200", 648=>x"a200", 649=>x"a000", 650=>x"9600", 651=>x"9400",
---- 652=>x"8e00", 653=>x"8900", 654=>x"8c00", 655=>x"8400", 656=>x"b000", 657=>x"9700", 658=>x"9800",
---- 659=>x"9600", 660=>x"9000", 661=>x"7d00", 662=>x"8b00", 663=>x"8400", 664=>x"ae00", 665=>x"a300",
---- 666=>x"9400", 667=>x"9e00", 668=>x"9400", 669=>x"8b00", 670=>x"8d00", 671=>x"8e00", 672=>x"b500",
---- 673=>x"a800", 674=>x"a200", 675=>x"9d00", 676=>x"9a00", 677=>x"8f00", 678=>x"8c00", 679=>x"9100",
---- 680=>x"b700", 681=>x"a900", 682=>x"aa00", 683=>x"5d00", 684=>x"9b00", 685=>x"8c00", 686=>x"9100",
---- 687=>x"9800", 688=>x"b300", 689=>x"ac00", 690=>x"a100", 691=>x"a900", 692=>x"9800", 693=>x"a500",
---- 694=>x"9200", 695=>x"9c00", 696=>x"bc00", 697=>x"a400", 698=>x"a800", 699=>x"9f00", 700=>x"a000",
---- 701=>x"9200", 702=>x"9f00", 703=>x"9400", 704=>x"ba00", 705=>x"b600", 706=>x"a600", 707=>x"a600",
---- 708=>x"9100", 709=>x"9b00", 710=>x"8e00", 711=>x"a000", 712=>x"c500", 713=>x"b600", 714=>x"b600",
---- 715=>x"a300", 716=>x"9800", 717=>x"8400", 718=>x"6f00", 719=>x"9200", 720=>x"bd00", 721=>x"c600",
---- 722=>x"b100", 723=>x"a900", 724=>x"8c00", 725=>x"7900", 726=>x"7b00", 727=>x"8f00", 728=>x"d000",
---- 729=>x"c200", 730=>x"b900", 731=>x"9e00", 732=>x"9200", 733=>x"7c00", 734=>x"7a00", 735=>x"8900",
---- 736=>x"c400", 737=>x"ca00", 738=>x"4600", 739=>x"ac00", 740=>x"8700", 741=>x"7400", 742=>x"6f00",
---- 743=>x"7b00", 744=>x"ca00", 745=>x"c600", 746=>x"bf00", 747=>x"a200", 748=>x"9300", 749=>x"8800",
---- 750=>x"6c00", 751=>x"9c00", 752=>x"c500", 753=>x"d100", 754=>x"c000", 755=>x"a200", 756=>x"8800",
---- 757=>x"7c00", 758=>x"8a00", 759=>x"9400", 760=>x"c700", 761=>x"c300", 762=>x"c400", 763=>x"a200",
---- 764=>x"9400", 765=>x"8400", 766=>x"8700", 767=>x"8a00", 768=>x"c000", 769=>x"c500", 770=>x"be00",
---- 771=>x"b700", 772=>x"9b00", 773=>x"8600", 774=>x"7400", 775=>x"9700", 776=>x"c800", 777=>x"bd00",
---- 778=>x"ca00", 779=>x"b700", 780=>x"a800", 781=>x"a000", 782=>x"8700", 783=>x"8600", 784=>x"c100",
---- 785=>x"c900", 786=>x"c100", 787=>x"c600", 788=>x"ba00", 789=>x"9c00", 790=>x"a900", 791=>x"8e00",
---- 792=>x"cd00", 793=>x"c500", 794=>x"c600", 795=>x"c500", 796=>x"a300", 797=>x"ac00", 798=>x"aa00",
---- 799=>x"a400", 800=>x"cf00", 801=>x"cd00", 802=>x"cc00", 803=>x"b400", 804=>x"9f00", 805=>x"af00",
---- 806=>x"b400", 807=>x"a400", 808=>x"de00", 809=>x"d100", 810=>x"c900", 811=>x"c100", 812=>x"9d00",
---- 813=>x"a500", 814=>x"b400", 815=>x"b300", 816=>x"d100", 817=>x"d200", 818=>x"d400", 819=>x"c300",
---- 820=>x"b400", 821=>x"a800", 822=>x"b100", 823=>x"bf00", 824=>x"9900", 825=>x"e100", 826=>x"cf00",
---- 827=>x"bf00", 828=>x"c400", 829=>x"bb00", 830=>x"ba00", 831=>x"af00", 832=>x"6600", 833=>x"ca00",
---- 834=>x"d200", 835=>x"c200", 836=>x"c100", 837=>x"bf00", 838=>x"c700", 839=>x"9600", 840=>x"5100",
---- 841=>x"9f00", 842=>x"e100", 843=>x"cc00", 844=>x"c200", 845=>x"bf00", 846=>x"ca00", 847=>x"9a00",
---- 848=>x"5200", 849=>x"8d00", 850=>x"df00", 851=>x"d900", 852=>x"c900", 853=>x"c700", 854=>x"c600",
---- 855=>x"b000", 856=>x"5100", 857=>x"8a00", 858=>x"dd00", 859=>x"d500", 860=>x"d300", 861=>x"c800",
---- 862=>x"c600", 863=>x"b100", 864=>x"5300", 865=>x"8800", 866=>x"e000", 867=>x"d500", 868=>x"2800",
---- 869=>x"d200", 870=>x"c500", 871=>x"8f00", 872=>x"5200", 873=>x"8800", 874=>x"db00", 875=>x"d800",
---- 876=>x"d200", 877=>x"d900", 878=>x"b100", 879=>x"6f00", 880=>x"5900", 881=>x"7900", 882=>x"d900",
---- 883=>x"da00", 884=>x"d500", 885=>x"d400", 886=>x"9400", 887=>x"6200", 888=>x"6100", 889=>x"6600",
---- 890=>x"c600", 891=>x"dd00", 892=>x"da00", 893=>x"c500", 894=>x"7300", 895=>x"6900", 896=>x"6500",
---- 897=>x"5b00", 898=>x"a600", 899=>x"e100", 900=>x"dd00", 901=>x"b700", 902=>x"6d00", 903=>x"6e00",
---- 904=>x"6b00", 905=>x"6100", 906=>x"8500", 907=>x"dd00", 908=>x"e300", 909=>x"a400", 910=>x"6f00",
---- 911=>x"6f00", 912=>x"7000", 913=>x"6b00", 914=>x"6c00", 915=>x"b900", 916=>x"e900", 917=>x"a800",
---- 918=>x"6c00", 919=>x"7400", 920=>x"7300", 921=>x"6f00", 922=>x"6600", 923=>x"8800", 924=>x"e300",
---- 925=>x"c000", 926=>x"7400", 927=>x"7500", 928=>x"7500", 929=>x"7300", 930=>x"6e00", 931=>x"6f00",
---- 932=>x"c100", 933=>x"d100", 934=>x"8100", 935=>x"7700", 936=>x"7900", 937=>x"7400", 938=>x"7400",
---- 939=>x"7000", 940=>x"9000", 941=>x"c700", 942=>x"8600", 943=>x"7900", 944=>x"7600", 945=>x"7400",
---- 946=>x"7700", 947=>x"8000", 948=>x"7f00", 949=>x"9400", 950=>x"7a00", 951=>x"7500", 952=>x"6800",
---- 953=>x"6a00", 954=>x"8400", 955=>x"8800", 956=>x"5c00", 957=>x"6400", 958=>x"7500", 959=>x"6800",
---- 960=>x"7700", 961=>x"7a00", 962=>x"8d00", 963=>x"5f00", 964=>x"6000", 965=>x"8300", 966=>x"9500",
---- 967=>x"7300", 968=>x"7400", 969=>x"7500", 970=>x"a200", 971=>x"8a00", 972=>x"7b00", 973=>x"9400",
---- 974=>x"bc00", 975=>x"9700", 976=>x"ac00", 977=>x"9e00", 978=>x"9500", 979=>x"5000", 980=>x"3d00",
---- 981=>x"4a00", 982=>x"5a00", 983=>x"7700", 984=>x"c900", 985=>x"7a00", 986=>x"5500", 987=>x"2100",
---- 988=>x"2000", 989=>x"2200", 990=>x"2800", 991=>x"7400", 992=>x"b100", 993=>x"5600", 994=>x"3200",
---- 995=>x"3400", 996=>x"2a00", 997=>x"2a00", 998=>x"5200", 999=>x"7000", 1000=>x"6100", 1001=>x"8600",
---- 1002=>x"4400", 1003=>x"3100", 1004=>x"2400", 1005=>x"2700", 1006=>x"5300", 1007=>x"8f00", 1008=>x"9500",
---- 1009=>x"8200", 1010=>x"3100", 1011=>x"3d00", 1012=>x"3e00", 1013=>x"1d00", 1014=>x"4e00", 1015=>x"8600",
---- 1016=>x"9800", 1017=>x"af00", 1018=>x"7100", 1019=>x"7600", 1020=>x"8d00", 1021=>x"4e00", 1022=>x"6800",
---- 1023=>x"8100", 1024=>x"9700", 1025=>x"b500", 1026=>x"ad00", 1027=>x"a400", 1028=>x"ab00", 1029=>x"8900",
---- 1030=>x"6600", 1031=>x"5200", 1032=>x"9a00", 1033=>x"9a00", 1034=>x"7b00", 1035=>x"7d00", 1036=>x"9900",
---- 1037=>x"6f00", 1038=>x"3000", 1039=>x"2b00", 1040=>x"9d00", 1041=>x"9100", 1042=>x"6c00", 1043=>x"4000",
---- 1044=>x"5600", 1045=>x"5d00", 1046=>x"2c00", 1047=>x"2400", 1048=>x"8800", 1049=>x"8300", 1050=>x"5800",
---- 1051=>x"3b00", 1052=>x"4300", 1053=>x"3200", 1054=>x"2600", 1055=>x"1c00", 1056=>x"7800", 1057=>x"8500",
---- 1058=>x"5300", 1059=>x"4c00", 1060=>x"2d00", 1061=>x"2700", 1062=>x"2a00", 1063=>x"3500", 1064=>x"9900",
---- 1065=>x"7d00", 1066=>x"3700", 1067=>x"3e00", 1068=>x"2500", 1069=>x"2c00", 1070=>x"4b00", 1071=>x"6400",
---- 1072=>x"6a00", 1073=>x"4200", 1074=>x"2400", 1075=>x"2800", 1076=>x"2500", 1077=>x"4700", 1078=>x"7300",
---- 1079=>x"4800", 1080=>x"2800", 1081=>x"2b00", 1082=>x"2700", 1083=>x"2a00", 1084=>x"4100", 1085=>x"5f00",
---- 1086=>x"4500", 1087=>x"3600", 1088=>x"2b00", 1089=>x"2500", 1090=>x"2200", 1091=>x"3600", 1092=>x"6000",
---- 1093=>x"5400", 1094=>x"4900", 1095=>x"4b00", 1096=>x"2500", 1097=>x"3200", 1098=>x"4c00", 1099=>x"7700",
---- 1100=>x"7a00", 1101=>x"6500", 1102=>x"3900", 1103=>x"2a00", 1104=>x"5200", 1105=>x"6a00", 1106=>x"7600",
---- 1107=>x"5a00", 1108=>x"5a00", 1109=>x"4e00", 1110=>x"2000", 1111=>x"2500", 1112=>x"7e00", 1113=>x"4800",
---- 1114=>x"3000", 1115=>x"4800", 1116=>x"6b00", 1117=>x"2c00", 1118=>x"2300", 1119=>x"2c00", 1120=>x"8f00",
---- 1121=>x"7a00", 1122=>x"5600", 1123=>x"8300", 1124=>x"6e00", 1125=>x"af00", 1126=>x"4300", 1127=>x"3100",
---- 1128=>x"4600", 1129=>x"8d00", 1130=>x"8f00", 1131=>x"8600", 1132=>x"7a00", 1133=>x"7600", 1134=>x"4b00",
---- 1135=>x"3200", 1136=>x"4a00", 1137=>x"6800", 1138=>x"6a00", 1139=>x"6300", 1140=>x"6700", 1141=>x"5300",
---- 1142=>x"3200", 1143=>x"2b00", 1144=>x"7300", 1145=>x"6900", 1146=>x"3400", 1147=>x"3a00", 1148=>x"6600",
---- 1149=>x"5000", 1150=>x"2800", 1151=>x"2600", 1152=>x"6f00", 1153=>x"5b00", 1154=>x"3c00", 1155=>x"6800",
---- 1156=>x"7100", 1157=>x"3200", 1158=>x"2100", 1159=>x"2a00", 1160=>x"5e00", 1161=>x"6100", 1162=>x"6d00",
---- 1163=>x"7600", 1164=>x"4400", 1165=>x"2400", 1166=>x"2700", 1167=>x"2700", 1168=>x"6300", 1169=>x"7f00",
---- 1170=>x"7600", 1171=>x"4f00", 1172=>x"2d00", 1173=>x"2d00", 1174=>x"2e00", 1175=>x"2700", 1176=>x"8a00",
---- 1177=>x"8500", 1178=>x"4900", 1179=>x"2f00", 1180=>x"3500", 1181=>x"3400", 1182=>x"2e00", 1183=>x"2f00",
---- 1184=>x"5700", 1185=>x"4d00", 1186=>x"4d00", 1187=>x"2e00", 1188=>x"3700", 1189=>x"2e00", 1190=>x"2e00",
---- 1191=>x"2e00", 1192=>x"4600", 1193=>x"4000", 1194=>x"5800", 1195=>x"3400", 1196=>x"2f00", 1197=>x"2b00",
---- 1198=>x"2d00", 1199=>x"3500", 1200=>x"5d00", 1201=>x"4000", 1202=>x"4600", 1203=>x"3500", 1204=>x"2900",
---- 1205=>x"2e00", 1206=>x"3700", 1207=>x"3300", 1208=>x"6400", 1209=>x"3800", 1210=>x"3a00", 1211=>x"3c00",
---- 1212=>x"3300", 1213=>x"3300", 1214=>x"3b00", 1215=>x"3000", 1216=>x"7600", 1217=>x"5000", 1218=>x"3100",
---- 1219=>x"3d00", 1220=>x"3a00", 1221=>x"3600", 1222=>x"3e00", 1223=>x"3400", 1224=>x"6800", 1225=>x"6e00",
---- 1226=>x"3000", 1227=>x"3500", 1228=>x"3e00", 1229=>x"3e00", 1230=>x"3b00", 1231=>x"3100", 1232=>x"5600",
---- 1233=>x"8100", 1234=>x"4200", 1235=>x"c600", 1236=>x"4000", 1237=>x"3a00", 1238=>x"3700", 1239=>x"3100",
---- 1240=>x"5d00", 1241=>x"7c00", 1242=>x"5700", 1243=>x"2e00", 1244=>x"3100", 1245=>x"c600", 1246=>x"3800",
---- 1247=>x"3000", 1248=>x"6200", 1249=>x"5000", 1250=>x"5600", 1251=>x"1f00", 1252=>x"2b00", 1253=>x"2e00",
---- 1254=>x"3500", 1255=>x"3200", 1256=>x"6c00", 1257=>x"3e00", 1258=>x"6b00", 1259=>x"2500", 1260=>x"2a00",
---- 1261=>x"3200", 1262=>x"2b00", 1263=>x"3000", 1264=>x"7e00", 1265=>x"3500", 1266=>x"6f00", 1267=>x"3f00",
---- 1268=>x"2200", 1269=>x"3000", 1270=>x"2f00", 1271=>x"4400", 1272=>x"8700", 1273=>x"3000", 1274=>x"5a00",
---- 1275=>x"5700", 1276=>x"2800", 1277=>x"3b00", 1278=>x"4500", 1279=>x"3600", 1280=>x"6400", 1281=>x"3a00",
---- 1282=>x"4d00", 1283=>x"7f00", 1284=>x"2f00", 1285=>x"3a00", 1286=>x"3600", 1287=>x"2900", 1288=>x"b100",
---- 1289=>x"5d00", 1290=>x"3d00", 1291=>x"9200", 1292=>x"4100", 1293=>x"2700", 1294=>x"3000", 1295=>x"3f00",
---- 1296=>x"a600", 1297=>x"8300", 1298=>x"3000", 1299=>x"8400", 1300=>x"4d00", 1301=>x"2600", 1302=>x"3000",
---- 1303=>x"4900", 1304=>x"8900", 1305=>x"9600", 1306=>x"3b00", 1307=>x"8200", 1308=>x"6300", 1309=>x"1900",
---- 1310=>x"2600", 1311=>x"2f00", 1312=>x"7800", 1313=>x"9c00", 1314=>x"6200", 1315=>x"7700", 1316=>x"7400",
---- 1317=>x"1c00", 1318=>x"2100", 1319=>x"3400", 1320=>x"6800", 1321=>x"8100", 1322=>x"8200", 1323=>x"7900",
---- 1324=>x"8400", 1325=>x"3500", 1326=>x"2000", 1327=>x"3600", 1328=>x"5100", 1329=>x"6400", 1330=>x"8c00",
---- 1331=>x"7c00", 1332=>x"9200", 1333=>x"5800", 1334=>x"2600", 1335=>x"3300", 1336=>x"5f00", 1337=>x"a600",
---- 1338=>x"9200", 1339=>x"6900", 1340=>x"8e00", 1341=>x"7500", 1342=>x"4500", 1343=>x"3d00", 1344=>x"6900",
---- 1345=>x"4d00", 1346=>x"7600", 1347=>x"6a00", 1348=>x"8900", 1349=>x"8000", 1350=>x"5600", 1351=>x"4600",
---- 1352=>x"5100", 1353=>x"4a00", 1354=>x"6800", 1355=>x"7c00", 1356=>x"8400", 1357=>x"8b00", 1358=>x"9e00",
---- 1359=>x"3500", 1360=>x"4800", 1361=>x"4100", 1362=>x"6e00", 1363=>x"8600", 1364=>x"7600", 1365=>x"7b00",
---- 1366=>x"7a00", 1367=>x"4900", 1368=>x"6000", 1369=>x"3700", 1370=>x"3c00", 1371=>x"7000", 1372=>x"8600",
---- 1373=>x"6e00", 1374=>x"7b00", 1375=>x"8600", 1376=>x"5e00", 1377=>x"5900", 1378=>x"2e00", 1379=>x"3f00",
---- 1380=>x"8100", 1381=>x"8300", 1382=>x"7a00", 1383=>x"9a00", 1384=>x"4300", 1385=>x"6900", 1386=>x"5800",
---- 1387=>x"3200", 1388=>x"4600", 1389=>x"5d00", 1390=>x"7000", 1391=>x"8800", 1392=>x"4400", 1393=>x"4700",
---- 1394=>x"7000", 1395=>x"5300", 1396=>x"3b00", 1397=>x"5d00", 1398=>x"6400", 1399=>x"7c00", 1400=>x"b200",
---- 1401=>x"3e00", 1402=>x"4900", 1403=>x"6e00", 1404=>x"6f00", 1405=>x"6e00", 1406=>x"4200", 1407=>x"6200",
---- 1408=>x"6a00", 1409=>x"5900", 1410=>x"4a00", 1411=>x"5800", 1412=>x"8e00", 1413=>x"7700", 1414=>x"3800",
---- 1415=>x"4900", 1416=>x"6600", 1417=>x"6a00", 1418=>x"6300", 1419=>x"5f00", 1420=>x"5b00", 1421=>x"5e00",
---- 1422=>x"5c00", 1423=>x"4300", 1424=>x"6f00", 1425=>x"5f00", 1426=>x"5100", 1427=>x"5e00", 1428=>x"3b00",
---- 1429=>x"3b00", 1430=>x"6d00", 1431=>x"6000", 1432=>x"6600", 1433=>x"7700", 1434=>x"6300", 1435=>x"5800",
---- 1436=>x"4500", 1437=>x"4200", 1438=>x"5200", 1439=>x"6300", 1440=>x"4000", 1441=>x"5c00", 1442=>x"8200",
---- 1443=>x"6500", 1444=>x"6a00", 1445=>x"5600", 1446=>x"6000", 1447=>x"6000", 1448=>x"5200", 1449=>x"3b00",
---- 1450=>x"5d00", 1451=>x"8200", 1452=>x"7000", 1453=>x"7200", 1454=>x"8a00", 1455=>x"6e00", 1456=>x"6300",
---- 1457=>x"4100", 1458=>x"3900", 1459=>x"5d00", 1460=>x"8200", 1461=>x"8600", 1462=>x"6d00", 1463=>x"7f00",
---- 1464=>x"6a00", 1465=>x"4900", 1466=>x"4700", 1467=>x"5000", 1468=>x"8800", 1469=>x"8a00", 1470=>x"7200",
---- 1471=>x"6f00", 1472=>x"7000", 1473=>x"5f00", 1474=>x"7300", 1475=>x"7200", 1476=>x"5b00", 1477=>x"7400",
---- 1478=>x"8400", 1479=>x"6b00", 1480=>x"6b00", 1481=>x"6d00", 1482=>x"7f00", 1483=>x"5000", 1484=>x"4e00",
---- 1485=>x"7000", 1486=>x"8300", 1487=>x"7500", 1488=>x"7000", 1489=>x"7300", 1490=>x"6400", 1491=>x"5100",
---- 1492=>x"ac00", 1493=>x"5500", 1494=>x"7c00", 1495=>x"7c00", 1496=>x"7c00", 1497=>x"7500", 1498=>x"7200",
---- 1499=>x"6800", 1500=>x"5200", 1501=>x"4600", 1502=>x"7c00", 1503=>x"7e00", 1504=>x"8200", 1505=>x"8500",
---- 1506=>x"7d00", 1507=>x"7a00", 1508=>x"6800", 1509=>x"4700", 1510=>x"7800", 1511=>x"8a00", 1512=>x"8700",
---- 1513=>x"8e00", 1514=>x"7200", 1515=>x"7b00", 1516=>x"8200", 1517=>x"6700", 1518=>x"7300", 1519=>x"9100",
---- 1520=>x"6a00", 1521=>x"7a00", 1522=>x"7700", 1523=>x"8400", 1524=>x"8c00", 1525=>x"7300", 1526=>x"6c00",
---- 1527=>x"7a00", 1528=>x"6700", 1529=>x"6700", 1530=>x"7400", 1531=>x"7b00", 1532=>x"8f00", 1533=>x"8a00",
---- 1534=>x"8800", 1535=>x"7500", 1536=>x"5800", 1537=>x"7100", 1538=>x"7500", 1539=>x"5f00", 1540=>x"6d00",
---- 1541=>x"9600", 1542=>x"7800", 1543=>x"7800", 1544=>x"4400", 1545=>x"7400", 1546=>x"7a00", 1547=>x"6c00",
---- 1548=>x"4f00", 1549=>x"7600", 1550=>x"5e00", 1551=>x"7b00", 1552=>x"3800", 1553=>x"5b00", 1554=>x"8c00",
---- 1555=>x"6f00", 1556=>x"3e00", 1557=>x"6b00", 1558=>x"8100", 1559=>x"a300", 1560=>x"3500", 1561=>x"3a00",
---- 1562=>x"5a00", 1563=>x"5b00", 1564=>x"5300", 1565=>x"8c00", 1566=>x"6600", 1567=>x"5800", 1568=>x"2d00",
---- 1569=>x"2e00", 1570=>x"5700", 1571=>x"7500", 1572=>x"7400", 1573=>x"9e00", 1574=>x"7600", 1575=>x"5800",
---- 1576=>x"2e00", 1577=>x"4000", 1578=>x"5f00", 1579=>x"7f00", 1580=>x"9200", 1581=>x"9500", 1582=>x"4e00",
---- 1583=>x"5a00", 1584=>x"7700", 1585=>x"7b00", 1586=>x"7b00", 1587=>x"9100", 1588=>x"a300", 1589=>x"6000",
---- 1590=>x"4a00", 1591=>x"4f00", 1592=>x"6100", 1593=>x"7300", 1594=>x"7d00", 1595=>x"9f00", 1596=>x"7a00",
---- 1597=>x"4300", 1598=>x"5400", 1599=>x"6500", 1600=>x"4a00", 1601=>x"5000", 1602=>x"5300", 1603=>x"8c00",
---- 1604=>x"4600", 1605=>x"5900", 1606=>x"6c00", 1607=>x"6100", 1608=>x"6e00", 1609=>x"5a00", 1610=>x"7a00",
---- 1611=>x"8100", 1612=>x"4100", 1613=>x"4400", 1614=>x"8d00", 1615=>x"7200", 1616=>x"7000", 1617=>x"8000",
---- 1618=>x"8200", 1619=>x"4e00", 1620=>x"4400", 1621=>x"4b00", 1622=>x"4700", 1623=>x"7600", 1624=>x"8100",
---- 1625=>x"6c00", 1626=>x"4b00", 1627=>x"3900", 1628=>x"4500", 1629=>x"5300", 1630=>x"4c00", 1631=>x"5100",
---- 1632=>x"6700", 1633=>x"3700", 1634=>x"4200", 1635=>x"4000", 1636=>x"3700", 1637=>x"4f00", 1638=>x"6500",
---- 1639=>x"4e00", 1640=>x"3f00", 1641=>x"3300", 1642=>x"4200", 1643=>x"4a00", 1644=>x"3d00", 1645=>x"3e00",
---- 1646=>x"5f00", 1647=>x"9900", 1648=>x"5100", 1649=>x"2b00", 1650=>x"3d00", 1651=>x"5000", 1652=>x"4d00",
---- 1653=>x"4400", 1654=>x"4700", 1655=>x"9300", 1656=>x"6d00", 1657=>x"3c00", 1658=>x"3000", 1659=>x"4600",
---- 1660=>x"4200", 1661=>x"4c00", 1662=>x"4b00", 1663=>x"5300", 1664=>x"6800", 1665=>x"6400", 1666=>x"3500",
---- 1667=>x"3300", 1668=>x"4600", 1669=>x"4a00", 1670=>x"4700", 1671=>x"4500", 1672=>x"5a00", 1673=>x"5400",
---- 1674=>x"5a00", 1675=>x"3700", 1676=>x"4100", 1677=>x"5000", 1678=>x"4c00", 1679=>x"b700", 1680=>x"a300",
---- 1681=>x"4200", 1682=>x"5200", 1683=>x"5d00", 1684=>x"3900", 1685=>x"5800", 1686=>x"6100", 1687=>x"4c00",
---- 1688=>x"5400", 1689=>x"4700", 1690=>x"3900", 1691=>x"6300", 1692=>x"5800", 1693=>x"4f00", 1694=>x"6900",
---- 1695=>x"6500", 1696=>x"4a00", 1697=>x"5000", 1698=>x"3100", 1699=>x"4b00", 1700=>x"5b00", 1701=>x"5400",
---- 1702=>x"5d00", 1703=>x"7400", 1704=>x"6100", 1705=>x"5c00", 1706=>x"3400", 1707=>x"4200", 1708=>x"4400",
---- 1709=>x"5d00", 1710=>x"5700", 1711=>x"7200", 1712=>x"3a00", 1713=>x"4600", 1714=>x"cf00", 1715=>x"4b00",
---- 1716=>x"4500", 1717=>x"5400", 1718=>x"5f00", 1719=>x"6400", 1720=>x"2100", 1721=>x"3200", 1722=>x"cc00",
---- 1723=>x"c000", 1724=>x"5200", 1725=>x"4500", 1726=>x"6700", 1727=>x"6000", 1728=>x"2e00", 1729=>x"2f00",
---- 1730=>x"3100", 1731=>x"3200", 1732=>x"4c00", 1733=>x"4300", 1734=>x"5900", 1735=>x"5c00", 1736=>x"3000",
---- 1737=>x"3400", 1738=>x"3300", 1739=>x"2c00", 1740=>x"4100", 1741=>x"4400", 1742=>x"4d00", 1743=>x"4f00",
---- 1744=>x"2b00", 1745=>x"3a00", 1746=>x"3d00", 1747=>x"2b00", 1748=>x"3b00", 1749=>x"4400", 1750=>x"3b00",
---- 1751=>x"3700", 1752=>x"2c00", 1753=>x"c500", 1754=>x"4100", 1755=>x"2600", 1756=>x"3600", 1757=>x"4b00",
---- 1758=>x"3700", 1759=>x"4300", 1760=>x"2a00", 1761=>x"3a00", 1762=>x"4500", 1763=>x"2500", 1764=>x"2f00",
---- 1765=>x"5c00", 1766=>x"3900", 1767=>x"3700", 1768=>x"2e00", 1769=>x"4100", 1770=>x"3a00", 1771=>x"2b00",
---- 1772=>x"3500", 1773=>x"5c00", 1774=>x"4300", 1775=>x"2d00", 1776=>x"2f00", 1777=>x"3c00", 1778=>x"4000",
---- 1779=>x"2d00", 1780=>x"4d00", 1781=>x"5d00", 1782=>x"3b00", 1783=>x"3500", 1784=>x"2700", 1785=>x"3800",
---- 1786=>x"3f00", 1787=>x"2900", 1788=>x"5800", 1789=>x"6300", 1790=>x"2700", 1791=>x"4000", 1792=>x"2700",
---- 1793=>x"3f00", 1794=>x"3300", 1795=>x"2a00", 1796=>x"5900", 1797=>x"6100", 1798=>x"2500", 1799=>x"3200",
---- 1800=>x"2f00", 1801=>x"4000", 1802=>x"2500", 1803=>x"3800", 1804=>x"5700", 1805=>x"4a00", 1806=>x"5300",
---- 1807=>x"2800", 1808=>x"3300", 1809=>x"4000", 1810=>x"2500", 1811=>x"4f00", 1812=>x"5600", 1813=>x"3400",
---- 1814=>x"6000", 1815=>x"5300", 1816=>x"3400", 1817=>x"3900", 1818=>x"3900", 1819=>x"4c00", 1820=>x"4300",
---- 1821=>x"3b00", 1822=>x"4c00", 1823=>x"6900", 1824=>x"2c00", 1825=>x"3400", 1826=>x"6200", 1827=>x"4300",
---- 1828=>x"2d00", 1829=>x"3700", 1830=>x"3600", 1831=>x"6400", 1832=>x"2400", 1833=>x"3d00", 1834=>x"6700",
---- 1835=>x"3c00", 1836=>x"2600", 1837=>x"2e00", 1838=>x"3b00", 1839=>x"6400", 1840=>x"2300", 1841=>x"4a00",
---- 1842=>x"4f00", 1843=>x"3000", 1844=>x"2f00", 1845=>x"2b00", 1846=>x"4c00", 1847=>x"7800", 1848=>x"2800",
---- 1849=>x"4d00", 1850=>x"3600", 1851=>x"2e00", 1852=>x"4200", 1853=>x"3100", 1854=>x"3b00", 1855=>x"7000",
---- 1856=>x"2b00", 1857=>x"3c00", 1858=>x"3000", 1859=>x"3500", 1860=>x"4800", 1861=>x"6100", 1862=>x"5800",
---- 1863=>x"6100", 1864=>x"3100", 1865=>x"2b00", 1866=>x"3400", 1867=>x"5c00", 1868=>x"2700", 1869=>x"5300",
---- 1870=>x"7a00", 1871=>x"5d00", 1872=>x"3400", 1873=>x"2e00", 1874=>x"3800", 1875=>x"4600", 1876=>x"1e00",
---- 1877=>x"2900", 1878=>x"5e00", 1879=>x"5100", 1880=>x"3800", 1881=>x"3800", 1882=>x"3000", 1883=>x"2500",
---- 1884=>x"2b00", 1885=>x"2e00", 1886=>x"2f00", 1887=>x"5800", 1888=>x"2b00", 1889=>x"3900", 1890=>x"3b00",
---- 1891=>x"2e00", 1892=>x"3400", 1893=>x"cc00", 1894=>x"2300", 1895=>x"3300", 1896=>x"2700", 1897=>x"2800",
---- 1898=>x"4100", 1899=>x"3a00", 1900=>x"2b00", 1901=>x"3a00", 1902=>x"2e00", 1903=>x"2b00", 1904=>x"3000",
---- 1905=>x"2800", 1906=>x"2e00", 1907=>x"3900", 1908=>x"3100", 1909=>x"4a00", 1910=>x"3c00", 1911=>x"3100",
---- 1912=>x"3200", 1913=>x"3500", 1914=>x"2200", 1915=>x"3400", 1916=>x"4600", 1917=>x"3f00", 1918=>x"4000",
---- 1919=>x"3000", 1920=>x"2d00", 1921=>x"3e00", 1922=>x"3700", 1923=>x"2700", 1924=>x"3d00", 1925=>x"4400",
---- 1926=>x"4000", 1927=>x"3700", 1928=>x"2500", 1929=>x"3a00", 1930=>x"4f00", 1931=>x"3900", 1932=>x"2800",
---- 1933=>x"3c00", 1934=>x"4c00", 1935=>x"3400", 1936=>x"2500", 1937=>x"3300", 1938=>x"5a00", 1939=>x"5b00",
---- 1940=>x"cb00", 1941=>x"3000", 1942=>x"5300", 1943=>x"3e00", 1944=>x"2b00", 1945=>x"3100", 1946=>x"5400",
---- 1947=>x"4f00", 1948=>x"4600", 1949=>x"3800", 1950=>x"4100", 1951=>x"5500", 1952=>x"3300", 1953=>x"2c00",
---- 1954=>x"5500", 1955=>x"4800", 1956=>x"2d00", 1957=>x"3400", 1958=>x"2f00", 1959=>x"6f00", 1960=>x"3100",
---- 1961=>x"2b00", 1962=>x"3d00", 1963=>x"6400", 1964=>x"2b00", 1965=>x"2c00", 1966=>x"3a00", 1967=>x"5500",
---- 1968=>x"3300", 1969=>x"3500", 1970=>x"2d00", 1971=>x"6000", 1972=>x"4700", 1973=>x"2a00", 1974=>x"3300",
---- 1975=>x"3600", 1976=>x"2900", 1977=>x"2900", 1978=>x"4500", 1979=>x"5700", 1980=>x"7100", 1981=>x"2a00",
---- 1982=>x"1e00", 1983=>x"3d00", 1984=>x"2900", 1985=>x"2400", 1986=>x"3900", 1987=>x"5e00", 1988=>x"7a00",
---- 1989=>x"5200", 1990=>x"1c00", 1991=>x"3100", 1992=>x"3c00", 1993=>x"2100", 1994=>x"2700", 1995=>x"5600",
---- 1996=>x"7800", 1997=>x"7000", 1998=>x"2e00", 1999=>x"1c00", 2000=>x"6200", 2001=>x"3400", 2002=>x"2a00",
---- 2003=>x"4900", 2004=>x"7100", 2005=>x"6e00", 2006=>x"4800", 2007=>x"2800", 2008=>x"8600", 2009=>x"4400",
---- 2010=>x"2800", 2011=>x"2d00", 2012=>x"5300", 2013=>x"6d00", 2014=>x"4200", 2015=>x"3f00", 2016=>x"9100",
---- 2017=>x"5800", 2018=>x"2600", 2019=>x"2800", 2020=>x"3500", 2021=>x"6c00", 2022=>x"4b00", 2023=>x"3800",
---- 2024=>x"7d00", 2025=>x"8500", 2026=>x"3600", 2027=>x"2700", 2028=>x"3b00", 2029=>x"6e00", 2030=>x"6d00",
---- 2031=>x"3400", 2032=>x"5200", 2033=>x"7f00", 2034=>x"6400", 2035=>x"2b00", 2036=>x"3900", 2037=>x"7400",
---- 2038=>x"7800", 2039=>x"4000", 2040=>x"4300", 2041=>x"5300", 2042=>x"8400", 2043=>x"5500", 2044=>x"2e00",
---- 2045=>x"7700", 2046=>x"7000", 2047=>x"3100"),
---- 9  => (0=>x"8300", 1=>x"7f00", 2=>x"8400", 3=>x"8200", 4=>x"8300", 5=>x"8100", 6=>x"8500", 7=>x"8700",
---- 8=>x"8200", 9=>x"7f00", 10=>x"8300", 11=>x"8200", 12=>x"8200", 13=>x"8000", 14=>x"8600",
---- 15=>x"8700", 16=>x"8300", 17=>x"7e00", 18=>x"8300", 19=>x"8200", 20=>x"8100", 21=>x"8100",
---- 22=>x"8600", 23=>x"8700", 24=>x"8100", 25=>x"8300", 26=>x"7b00", 27=>x"8200", 28=>x"8000",
---- 29=>x"8400", 30=>x"8300", 31=>x"8300", 32=>x"8300", 33=>x"8200", 34=>x"8300", 35=>x"8200",
---- 36=>x"8200", 37=>x"8200", 38=>x"8200", 39=>x"8300", 40=>x"8300", 41=>x"8300", 42=>x"8300",
---- 43=>x"8000", 44=>x"8200", 45=>x"8200", 46=>x"8000", 47=>x"8300", 48=>x"8400", 49=>x"8400",
---- 50=>x"8200", 51=>x"8100", 52=>x"8300", 53=>x"7d00", 54=>x"8100", 55=>x"8600", 56=>x"8200",
---- 57=>x"7c00", 58=>x"8200", 59=>x"8100", 60=>x"8200", 61=>x"8100", 62=>x"8300", 63=>x"8300",
---- 64=>x"8300", 65=>x"8300", 66=>x"8200", 67=>x"8300", 68=>x"8300", 69=>x"8300", 70=>x"8000",
---- 71=>x"8200", 72=>x"8100", 73=>x"8300", 74=>x"8500", 75=>x"8400", 76=>x"8500", 77=>x"8300",
---- 78=>x"8100", 79=>x"8200", 80=>x"8000", 81=>x"8500", 82=>x"8200", 83=>x"8300", 84=>x"8400",
---- 85=>x"8300", 86=>x"8200", 87=>x"8300", 88=>x"8100", 89=>x"8200", 90=>x"8200", 91=>x"8000",
---- 92=>x"8100", 93=>x"8000", 94=>x"8200", 95=>x"8200", 96=>x"8200", 97=>x"8100", 98=>x"8200",
---- 99=>x"8400", 100=>x"8000", 101=>x"8000", 102=>x"8100", 103=>x"8100", 104=>x"8000", 105=>x"8000",
---- 106=>x"7f00", 107=>x"8100", 108=>x"8000", 109=>x"8200", 110=>x"8400", 111=>x"8000", 112=>x"7f00",
---- 113=>x"7f00", 114=>x"8200", 115=>x"8000", 116=>x"8300", 117=>x"8200", 118=>x"8100", 119=>x"8300",
---- 120=>x"7f00", 121=>x"7d00", 122=>x"8000", 123=>x"8000", 124=>x"8000", 125=>x"8200", 126=>x"8100",
---- 127=>x"8000", 128=>x"7e00", 129=>x"7c00", 130=>x"7f00", 131=>x"8100", 132=>x"7f00", 133=>x"8300",
---- 134=>x"8100", 135=>x"8100", 136=>x"7f00", 137=>x"8100", 138=>x"7f00", 139=>x"7f00", 140=>x"7e00",
---- 141=>x"7f00", 142=>x"8100", 143=>x"8300", 144=>x"7f00", 145=>x"8000", 146=>x"7c00", 147=>x"7e00",
---- 148=>x"7b00", 149=>x"7d00", 150=>x"8100", 151=>x"8100", 152=>x"7d00", 153=>x"7d00", 154=>x"7a00",
---- 155=>x"7e00", 156=>x"7e00", 157=>x"7f00", 158=>x"7f00", 159=>x"8000", 160=>x"8000", 161=>x"7c00",
---- 162=>x"7b00", 163=>x"7c00", 164=>x"7d00", 165=>x"7d00", 166=>x"8100", 167=>x"7f00", 168=>x"7c00",
---- 169=>x"7d00", 170=>x"7e00", 171=>x"7e00", 172=>x"7f00", 173=>x"7f00", 174=>x"8100", 175=>x"7f00",
---- 176=>x"7c00", 177=>x"7d00", 178=>x"7d00", 179=>x"8000", 180=>x"8000", 181=>x"8200", 182=>x"8300",
---- 183=>x"8000", 184=>x"7e00", 185=>x"8000", 186=>x"7f00", 187=>x"8300", 188=>x"8000", 189=>x"7f00",
---- 190=>x"8300", 191=>x"8100", 192=>x"7d00", 193=>x"7e00", 194=>x"7f00", 195=>x"8100", 196=>x"7f00",
---- 197=>x"8200", 198=>x"8000", 199=>x"7e00", 200=>x"7e00", 201=>x"8100", 202=>x"8200", 203=>x"8000",
---- 204=>x"8100", 205=>x"8200", 206=>x"8200", 207=>x"7c00", 208=>x"7e00", 209=>x"8400", 210=>x"8100",
---- 211=>x"8000", 212=>x"8000", 213=>x"8100", 214=>x"8100", 215=>x"7d00", 216=>x"8300", 217=>x"8200",
---- 218=>x"7e00", 219=>x"7e00", 220=>x"7e00", 221=>x"8000", 222=>x"8300", 223=>x"8100", 224=>x"7f00",
---- 225=>x"7d00", 226=>x"8100", 227=>x"7e00", 228=>x"8000", 229=>x"8100", 230=>x"8000", 231=>x"8000",
---- 232=>x"7d00", 233=>x"7f00", 234=>x"7d00", 235=>x"7e00", 236=>x"7f00", 237=>x"8000", 238=>x"8000",
---- 239=>x"8000", 240=>x"7c00", 241=>x"8000", 242=>x"7e00", 243=>x"8000", 244=>x"7f00", 245=>x"7f00",
---- 246=>x"7b00", 247=>x"7b00", 248=>x"7f00", 249=>x"7e00", 250=>x"7e00", 251=>x"7d00", 252=>x"7d00",
---- 253=>x"7f00", 254=>x"7800", 255=>x"8500", 256=>x"7d00", 257=>x"7a00", 258=>x"7d00", 259=>x"7c00",
---- 260=>x"7b00", 261=>x"7b00", 262=>x"7b00", 263=>x"a900", 264=>x"7d00", 265=>x"8300", 266=>x"7d00",
---- 267=>x"7a00", 268=>x"7900", 269=>x"7600", 270=>x"9b00", 271=>x"a800", 272=>x"7c00", 273=>x"7c00",
---- 274=>x"7c00", 275=>x"7c00", 276=>x"7d00", 277=>x"7500", 278=>x"6400", 279=>x"8e00", 280=>x"7f00",
---- 281=>x"7a00", 282=>x"7e00", 283=>x"7f00", 284=>x"7d00", 285=>x"8600", 286=>x"7400", 287=>x"6a00",
---- 288=>x"7d00", 289=>x"7900", 290=>x"7a00", 291=>x"7700", 292=>x"8100", 293=>x"9100", 294=>x"7000",
---- 295=>x"6f00", 296=>x"7c00", 297=>x"7b00", 298=>x"7a00", 299=>x"7900", 300=>x"ac00", 301=>x"8900",
---- 302=>x"6a00", 303=>x"7300", 304=>x"7d00", 305=>x"7d00", 306=>x"7600", 307=>x"8a00", 308=>x"a500",
---- 309=>x"7400", 310=>x"7200", 311=>x"7300", 312=>x"7c00", 313=>x"7c00", 314=>x"7900", 315=>x"9500",
---- 316=>x"8400", 317=>x"7000", 318=>x"7300", 319=>x"6b00", 320=>x"7c00", 321=>x"7e00", 322=>x"8300",
---- 323=>x"8500", 324=>x"7700", 325=>x"7000", 326=>x"6c00", 327=>x"6d00", 328=>x"7c00", 329=>x"7d00",
---- 330=>x"8200", 331=>x"7b00", 332=>x"6d00", 333=>x"6d00", 334=>x"6c00", 335=>x"6e00", 336=>x"7c00",
---- 337=>x"8400", 338=>x"7c00", 339=>x"6d00", 340=>x"6d00", 341=>x"6a00", 342=>x"6f00", 343=>x"6d00",
---- 344=>x"7e00", 345=>x"8000", 346=>x"7000", 347=>x"6800", 348=>x"6a00", 349=>x"6c00", 350=>x"6f00",
---- 351=>x"7000", 352=>x"7c00", 353=>x"7200", 354=>x"6e00", 355=>x"6c00", 356=>x"6a00", 357=>x"6b00",
---- 358=>x"6f00", 359=>x"7300", 360=>x"7000", 361=>x"6c00", 362=>x"6a00", 363=>x"6b00", 364=>x"6d00",
---- 365=>x"6d00", 366=>x"6f00", 367=>x"7300", 368=>x"6a00", 369=>x"6e00", 370=>x"6b00", 371=>x"6e00",
---- 372=>x"7300", 373=>x"7100", 374=>x"7100", 375=>x"6f00", 376=>x"6d00", 377=>x"6900", 378=>x"6f00",
---- 379=>x"7500", 380=>x"6f00", 381=>x"6f00", 382=>x"7400", 383=>x"7000", 384=>x"6f00", 385=>x"7000",
---- 386=>x"6e00", 387=>x"7100", 388=>x"7200", 389=>x"7000", 390=>x"7000", 391=>x"7400", 392=>x"7200",
---- 393=>x"7500", 394=>x"6e00", 395=>x"9200", 396=>x"6e00", 397=>x"7000", 398=>x"7100", 399=>x"7400",
---- 400=>x"6d00", 401=>x"7400", 402=>x"7400", 403=>x"6d00", 404=>x"6d00", 405=>x"6e00", 406=>x"7100",
---- 407=>x"7100", 408=>x"6b00", 409=>x"7100", 410=>x"7400", 411=>x"7100", 412=>x"7200", 413=>x"7000",
---- 414=>x"7000", 415=>x"6f00", 416=>x"6700", 417=>x"6c00", 418=>x"7600", 419=>x"7400", 420=>x"7300",
---- 421=>x"7100", 422=>x"7100", 423=>x"7500", 424=>x"6900", 425=>x"6c00", 426=>x"7000", 427=>x"7100",
---- 428=>x"7300", 429=>x"7000", 430=>x"6e00", 431=>x"6f00", 432=>x"6800", 433=>x"7200", 434=>x"6f00",
---- 435=>x"7000", 436=>x"6f00", 437=>x"7100", 438=>x"7100", 439=>x"7200", 440=>x"6c00", 441=>x"6d00",
---- 442=>x"6d00", 443=>x"7100", 444=>x"6c00", 445=>x"7000", 446=>x"7300", 447=>x"7100", 448=>x"6c00",
---- 449=>x"6d00", 450=>x"6b00", 451=>x"6f00", 452=>x"6e00", 453=>x"8e00", 454=>x"7200", 455=>x"7200",
---- 456=>x"6900", 457=>x"7000", 458=>x"6f00", 459=>x"6d00", 460=>x"7300", 461=>x"7100", 462=>x"6c00",
---- 463=>x"6b00", 464=>x"6b00", 465=>x"6c00", 466=>x"7400", 467=>x"7700", 468=>x"6f00", 469=>x"6e00",
---- 470=>x"7400", 471=>x"6c00", 472=>x"6e00", 473=>x"6d00", 474=>x"7000", 475=>x"7400", 476=>x"7000",
---- 477=>x"7100", 478=>x"7500", 479=>x"7500", 480=>x"7000", 481=>x"6c00", 482=>x"6900", 483=>x"7400",
---- 484=>x"7300", 485=>x"7400", 486=>x"7300", 487=>x"7800", 488=>x"6e00", 489=>x"6700", 490=>x"6f00",
---- 491=>x"7b00", 492=>x"6e00", 493=>x"7000", 494=>x"7400", 495=>x"7300", 496=>x"6900", 497=>x"6d00",
---- 498=>x"7200", 499=>x"8600", 500=>x"7000", 501=>x"6800", 502=>x"7900", 503=>x"7200", 504=>x"6a00",
---- 505=>x"7200", 506=>x"7400", 507=>x"6b00", 508=>x"6000", 509=>x"6f00", 510=>x"7500", 511=>x"6f00",
---- 512=>x"6d00", 513=>x"9500", 514=>x"6600", 515=>x"5e00", 516=>x"6d00", 517=>x"7700", 518=>x"7700",
---- 519=>x"7800", 520=>x"6a00", 521=>x"5e00", 522=>x"5b00", 523=>x"7300", 524=>x"7500", 525=>x"7200",
---- 526=>x"7500", 527=>x"8200", 528=>x"6300", 529=>x"6400", 530=>x"7000", 531=>x"7b00", 532=>x"7200",
---- 533=>x"7800", 534=>x"7500", 535=>x"7500", 536=>x"6a00", 537=>x"7200", 538=>x"6f00", 539=>x"6f00",
---- 540=>x"7300", 541=>x"6f00", 542=>x"6800", 543=>x"7600", 544=>x"6e00", 545=>x"8e00", 546=>x"6500",
---- 547=>x"6d00", 548=>x"6c00", 549=>x"6200", 550=>x"7200", 551=>x"7800", 552=>x"6a00", 553=>x"6400",
---- 554=>x"6700", 555=>x"6000", 556=>x"6600", 557=>x"7400", 558=>x"7700", 559=>x"7700", 560=>x"6100",
---- 561=>x"6500", 562=>x"6000", 563=>x"6800", 564=>x"6900", 565=>x"6b00", 566=>x"7200", 567=>x"6700",
---- 568=>x"6f00", 569=>x"6700", 570=>x"6600", 571=>x"6a00", 572=>x"6800", 573=>x"7000", 574=>x"6a00",
---- 575=>x"6c00", 576=>x"6b00", 577=>x"6e00", 578=>x"6900", 579=>x"6c00", 580=>x"6a00", 581=>x"6b00",
---- 582=>x"7200", 583=>x"7000", 584=>x"6a00", 585=>x"6300", 586=>x"6900", 587=>x"7000", 588=>x"6c00",
---- 589=>x"7200", 590=>x"7500", 591=>x"7000", 592=>x"6600", 593=>x"6600", 594=>x"6a00", 595=>x"6e00",
---- 596=>x"6f00", 597=>x"7200", 598=>x"7900", 599=>x"7700", 600=>x"6d00", 601=>x"6900", 602=>x"6900",
---- 603=>x"6900", 604=>x"6f00", 605=>x"7300", 606=>x"6400", 607=>x"6c00", 608=>x"6900", 609=>x"6a00",
---- 610=>x"6800", 611=>x"6d00", 612=>x"6d00", 613=>x"6600", 614=>x"6300", 615=>x"7400", 616=>x"6800",
---- 617=>x"6800", 618=>x"6a00", 619=>x"6b00", 620=>x"6800", 621=>x"7400", 622=>x"6e00", 623=>x"7200",
---- 624=>x"7300", 625=>x"7000", 626=>x"5e00", 627=>x"5a00", 628=>x"7000", 629=>x"6b00", 630=>x"6e00",
---- 631=>x"7b00", 632=>x"7800", 633=>x"6700", 634=>x"5c00", 635=>x"6300", 636=>x"6100", 637=>x"6900",
---- 638=>x"7700", 639=>x"7400", 640=>x"7000", 641=>x"6600", 642=>x"6700", 643=>x"5b00", 644=>x"5c00",
---- 645=>x"6f00", 646=>x"6f00", 647=>x"6d00", 648=>x"6a00", 649=>x"6b00", 650=>x"6200", 651=>x"6600",
---- 652=>x"6e00", 653=>x"6c00", 654=>x"6c00", 655=>x"6100", 656=>x"7400", 657=>x"7200", 658=>x"6b00",
---- 659=>x"6900", 660=>x"6b00", 661=>x"6d00", 662=>x"6400", 663=>x"7c00", 664=>x"7900", 665=>x"7b00",
---- 666=>x"7200", 667=>x"6a00", 668=>x"6700", 669=>x"5e00", 670=>x"7600", 671=>x"8600", 672=>x"8100",
---- 673=>x"7700", 674=>x"6a00", 675=>x"9600", 676=>x"a400", 677=>x"7300", 678=>x"8d00", 679=>x"8800",
---- 680=>x"8e00", 681=>x"7c00", 682=>x"7100", 683=>x"a600", 684=>x"6500", 685=>x"8600", 686=>x"8a00",
---- 687=>x"8b00", 688=>x"9200", 689=>x"8700", 690=>x"6c00", 691=>x"6200", 692=>x"7800", 693=>x"8300",
---- 694=>x"8100", 695=>x"8200", 696=>x"9d00", 697=>x"8600", 698=>x"7100", 699=>x"7a00", 700=>x"7a00",
---- 701=>x"7e00", 702=>x"7c00", 703=>x"7d00", 704=>x"9300", 705=>x"8800", 706=>x"7b00", 707=>x"7500",
---- 708=>x"7a00", 709=>x"7600", 710=>x"7400", 711=>x"7c00", 712=>x"9f00", 713=>x"9600", 714=>x"7300",
---- 715=>x"6d00", 716=>x"7300", 717=>x"7c00", 718=>x"7200", 719=>x"7a00", 720=>x"9c00", 721=>x"7800",
---- 722=>x"6900", 723=>x"6c00", 724=>x"7100", 725=>x"7c00", 726=>x"7c00", 727=>x"8000", 728=>x"7f00",
---- 729=>x"7400", 730=>x"7100", 731=>x"7000", 732=>x"6f00", 733=>x"7100", 734=>x"8400", 735=>x"7100",
---- 736=>x"8800", 737=>x"8100", 738=>x"7300", 739=>x"8800", 740=>x"7400", 741=>x"7600", 742=>x"7600",
---- 743=>x"6700", 744=>x"8f00", 745=>x"9300", 746=>x"7e00", 747=>x"7900", 748=>x"8000", 749=>x"6f00",
---- 750=>x"6100", 751=>x"6f00", 752=>x"9500", 753=>x"8200", 754=>x"8f00", 755=>x"7f00", 756=>x"7200",
---- 757=>x"6600", 758=>x"6b00", 759=>x"7200", 760=>x"9200", 761=>x"9600", 762=>x"8900", 763=>x"8400",
---- 764=>x"6400", 765=>x"6900", 766=>x"7000", 767=>x"7500", 768=>x"8c00", 769=>x"9800", 770=>x"8e00",
---- 771=>x"6c00", 772=>x"6300", 773=>x"7600", 774=>x"7700", 775=>x"8400", 776=>x"9a00", 777=>x"7d00",
---- 778=>x"7700", 779=>x"6b00", 780=>x"6d00", 781=>x"8c00", 782=>x"8400", 783=>x"8b00", 784=>x"a100",
---- 785=>x"8c00", 786=>x"6400", 787=>x"6900", 788=>x"7a00", 789=>x"7e00", 790=>x"8900", 791=>x"8500",
---- 792=>x"9100", 793=>x"8e00", 794=>x"5e00", 795=>x"7100", 796=>x"8000", 797=>x"8100", 798=>x"8b00",
---- 799=>x"8800", 800=>x"8c00", 801=>x"6000", 802=>x"6300", 803=>x"7e00", 804=>x"8300", 805=>x"7900",
---- 806=>x"7f00", 807=>x"8a00", 808=>x"9300", 809=>x"5c00", 810=>x"7100", 811=>x"8c00", 812=>x"8200",
---- 813=>x"8300", 814=>x"7c00", 815=>x"8000", 816=>x"9000", 817=>x"6e00", 818=>x"8400", 819=>x"8400",
---- 820=>x"8100", 821=>x"8400", 822=>x"8000", 823=>x"7400", 824=>x"6d00", 825=>x"8200", 826=>x"8c00",
---- 827=>x"7400", 828=>x"8200", 829=>x"8400", 830=>x"7d00", 831=>x"7400", 832=>x"6b00", 833=>x"9400",
---- 834=>x"7f00", 835=>x"7100", 836=>x"7a00", 837=>x"7d00", 838=>x"7100", 839=>x"7500", 840=>x"8800",
---- 841=>x"8c00", 842=>x"7700", 843=>x"7300", 844=>x"7600", 845=>x"7000", 846=>x"6600", 847=>x"7600",
---- 848=>x"9400", 849=>x"7800", 850=>x"8300", 851=>x"7d00", 852=>x"7200", 853=>x"6300", 854=>x"6d00",
---- 855=>x"7900", 856=>x"8600", 857=>x"7800", 858=>x"7c00", 859=>x"7e00", 860=>x"7500", 861=>x"9600",
---- 862=>x"7700", 863=>x"7c00", 864=>x"6900", 865=>x"7400", 866=>x"7e00", 867=>x"7800", 868=>x"7400",
---- 869=>x"7b00", 870=>x"7e00", 871=>x"7a00", 872=>x"6300", 873=>x"7600", 874=>x"7b00", 875=>x"7400",
---- 876=>x"7700", 877=>x"7b00", 878=>x"7d00", 879=>x"7100", 880=>x"6600", 881=>x"6e00", 882=>x"7300",
---- 883=>x"7000", 884=>x"7500", 885=>x"7800", 886=>x"7100", 887=>x"6c00", 888=>x"6c00", 889=>x"6900",
---- 890=>x"6b00", 891=>x"7400", 892=>x"7200", 893=>x"7500", 894=>x"6e00", 895=>x"7b00", 896=>x"7200",
---- 897=>x"7300", 898=>x"6e00", 899=>x"7300", 900=>x"6b00", 901=>x"6800", 902=>x"8000", 903=>x"8800",
---- 904=>x"7700", 905=>x"7a00", 906=>x"7400", 907=>x"6800", 908=>x"6400", 909=>x"7a00", 910=>x"8800",
---- 911=>x"7e00", 912=>x"7300", 913=>x"7700", 914=>x"7600", 915=>x"6900", 916=>x"7800", 917=>x"7e00",
---- 918=>x"7f00", 919=>x"7d00", 920=>x"7000", 921=>x"6b00", 922=>x"7300", 923=>x"7f00", 924=>x"8200",
---- 925=>x"7900", 926=>x"7600", 927=>x"8500", 928=>x"7300", 929=>x"6900", 930=>x"7b00", 931=>x"8300",
---- 932=>x"7900", 933=>x"8400", 934=>x"8400", 935=>x"7d00", 936=>x"6a00", 937=>x"7300", 938=>x"7800",
---- 939=>x"8500", 940=>x"8100", 941=>x"8200", 942=>x"8800", 943=>x"8300", 944=>x"7100", 945=>x"8300",
---- 946=>x"8900", 947=>x"8700", 948=>x"8a00", 949=>x"7f00", 950=>x"7e00", 951=>x"7d00", 952=>x"8100",
---- 953=>x"7f00", 954=>x"8600", 955=>x"7400", 956=>x"7d00", 957=>x"7f00", 958=>x"7c00", 959=>x"6700",
---- 960=>x"7800", 961=>x"7f00", 962=>x"7f00", 963=>x"8100", 964=>x"7d00", 965=>x"7400", 966=>x"7c00",
---- 967=>x"7100", 968=>x"7100", 969=>x"7b00", 970=>x"7f00", 971=>x"8500", 972=>x"7800", 973=>x"7600",
---- 974=>x"8100", 975=>x"5700", 976=>x"8200", 977=>x"7800", 978=>x"8100", 979=>x"7f00", 980=>x"7000",
---- 981=>x"7a00", 982=>x"7000", 983=>x"3800", 984=>x"9d00", 985=>x"ac00", 986=>x"8400", 987=>x"6e00",
---- 988=>x"6700", 989=>x"6600", 990=>x"3b00", 991=>x"3300", 992=>x"b300", 993=>x"c100", 994=>x"8800",
---- 995=>x"5800", 996=>x"4a00", 997=>x"5200", 998=>x"3600", 999=>x"3a00", 1000=>x"8c00", 1001=>x"6000",
---- 1002=>x"6a00", 1003=>x"4800", 1004=>x"4a00", 1005=>x"5400", 1006=>x"3600", 1007=>x"4800", 1008=>x"7e00",
---- 1009=>x"5500", 1010=>x"ac00", 1011=>x"5c00", 1012=>x"4600", 1013=>x"4000", 1014=>x"3c00", 1015=>x"5f00",
---- 1016=>x"9000", 1017=>x"7000", 1018=>x"4100", 1019=>x"4900", 1020=>x"2f00", 1021=>x"3600", 1022=>x"4700",
---- 1023=>x"6e00", 1024=>x"5800", 1025=>x"4100", 1026=>x"3900", 1027=>x"3800", 1028=>x"3400", 1029=>x"4d00",
---- 1030=>x"6500", 1031=>x"6e00", 1032=>x"2100", 1033=>x"2200", 1034=>x"bf00", 1035=>x"5200", 1036=>x"5000",
---- 1037=>x"5b00", 1038=>x"8400", 1039=>x"5100", 1040=>x"1f00", 1041=>x"4100", 1042=>x"7100", 1043=>x"5b00",
---- 1044=>x"4700", 1045=>x"7400", 1046=>x"6700", 1047=>x"5700", 1048=>x"4400", 1049=>x"7f00", 1050=>x"5c00",
---- 1051=>x"3100", 1052=>x"5800", 1053=>x"6100", 1054=>x"3100", 1055=>x"4f00", 1056=>x"7600", 1057=>x"5f00",
---- 1058=>x"2300", 1059=>x"4400", 1060=>x"6a00", 1061=>x"2a00", 1062=>x"2200", 1063=>x"4100", 1064=>x"4600",
---- 1065=>x"2600", 1066=>x"c700", 1067=>x"5a00", 1068=>x"4000", 1069=>x"d700", 1070=>x"2900", 1071=>x"4800",
---- 1072=>x"2500", 1073=>x"3900", 1074=>x"5000", 1075=>x"3800", 1076=>x"4700", 1077=>x"3800", 1078=>x"2b00",
---- 1079=>x"4b00", 1080=>x"3400", 1081=>x"4900", 1082=>x"4600", 1083=>x"3700", 1084=>x"4600", 1085=>x"4400",
---- 1086=>x"3c00", 1087=>x"5e00", 1088=>x"3600", 1089=>x"3f00", 1090=>x"5200", 1091=>x"4a00", 1092=>x"b000",
---- 1093=>x"5a00", 1094=>x"5000", 1095=>x"6300", 1096=>x"2100", 1097=>x"4500", 1098=>x"4700", 1099=>x"5400",
---- 1100=>x"5800", 1101=>x"4e00", 1102=>x"4b00", 1103=>x"6800", 1104=>x"2700", 1105=>x"5f00", 1106=>x"3f00",
---- 1107=>x"4f00", 1108=>x"5500", 1109=>x"4700", 1110=>x"5100", 1111=>x"6600", 1112=>x"3000", 1113=>x"5e00",
---- 1114=>x"4900", 1115=>x"4e00", 1116=>x"6500", 1117=>x"3700", 1118=>x"4000", 1119=>x"6800", 1120=>x"2700",
---- 1121=>x"4d00", 1122=>x"4e00", 1123=>x"4300", 1124=>x"6900", 1125=>x"4900", 1126=>x"3600", 1127=>x"6b00",
---- 1128=>x"2700", 1129=>x"3900", 1130=>x"5600", 1131=>x"3d00", 1132=>x"5e00", 1133=>x"6e00", 1134=>x"5100",
---- 1135=>x"5700", 1136=>x"2600", 1137=>x"3700", 1138=>x"4900", 1139=>x"4200", 1140=>x"3700", 1141=>x"7000",
---- 1142=>x"7800", 1143=>x"5600", 1144=>x"3000", 1145=>x"3400", 1146=>x"4900", 1147=>x"5a00", 1148=>x"3300",
---- 1149=>x"3400", 1150=>x"7900", 1151=>x"9700", 1152=>x"2e00", 1153=>x"3700", 1154=>x"5f00", 1155=>x"7900",
---- 1156=>x"5900", 1157=>x"3c00", 1158=>x"4900", 1159=>x"6200", 1160=>x"3000", 1161=>x"3000", 1162=>x"3a00",
---- 1163=>x"6000", 1164=>x"6b00", 1165=>x"6600", 1166=>x"6900", 1167=>x"5500", 1168=>x"2c00", 1169=>x"d300",
---- 1170=>x"2a00", 1171=>x"3d00", 1172=>x"5300", 1173=>x"5300", 1174=>x"7900", 1175=>x"8300", 1176=>x"2e00",
---- 1177=>x"2e00", 1178=>x"2e00", 1179=>x"3000", 1180=>x"4300", 1181=>x"5100", 1182=>x"4200", 1183=>x"4b00",
---- 1184=>x"d200", 1185=>x"2d00", 1186=>x"3300", 1187=>x"3300", 1188=>x"2c00", 1189=>x"4900", 1190=>x"5100",
---- 1191=>x"3100", 1192=>x"3200", 1193=>x"2e00", 1194=>x"cb00", 1195=>x"3300", 1196=>x"2e00", 1197=>x"3900",
---- 1198=>x"3c00", 1199=>x"3900", 1200=>x"3500", 1201=>x"3200", 1202=>x"3100", 1203=>x"3200", 1204=>x"3200",
---- 1205=>x"3a00", 1206=>x"2e00", 1207=>x"2b00", 1208=>x"2e00", 1209=>x"3300", 1210=>x"2e00", 1211=>x"2f00",
---- 1212=>x"2f00", 1213=>x"3000", 1214=>x"5600", 1215=>x"3b00", 1216=>x"2e00", 1217=>x"2d00", 1218=>x"2a00",
---- 1219=>x"2f00", 1220=>x"2900", 1221=>x"2f00", 1222=>x"5400", 1223=>x"3b00", 1224=>x"d800", 1225=>x"2800",
---- 1226=>x"2800", 1227=>x"2c00", 1228=>x"2b00", 1229=>x"3100", 1230=>x"4b00", 1231=>x"4900", 1232=>x"2500",
---- 1233=>x"2700", 1234=>x"2200", 1235=>x"2600", 1236=>x"3200", 1237=>x"4a00", 1238=>x"6f00", 1239=>x"5c00",
---- 1240=>x"2400", 1241=>x"2900", 1242=>x"2400", 1243=>x"3400", 1244=>x"3700", 1245=>x"4000", 1246=>x"7100",
---- 1247=>x"6d00", 1248=>x"2900", 1249=>x"2a00", 1250=>x"2800", 1251=>x"3000", 1252=>x"3e00", 1253=>x"af00",
---- 1254=>x"5000", 1255=>x"5e00", 1256=>x"3500", 1257=>x"3300", 1258=>x"2f00", 1259=>x"2a00", 1260=>x"3500",
---- 1261=>x"5d00", 1262=>x"4100", 1263=>x"4700", 1264=>x"3e00", 1265=>x"2800", 1266=>x"2200", 1267=>x"2900",
---- 1268=>x"3c00", 1269=>x"4800", 1270=>x"4f00", 1271=>x"6c00", 1272=>x"2c00", 1273=>x"3500", 1274=>x"2800",
---- 1275=>x"2800", 1276=>x"3e00", 1277=>x"4c00", 1278=>x"8200", 1279=>x"8500", 1280=>x"3000", 1281=>x"4d00",
---- 1282=>x"2c00", 1283=>x"2100", 1284=>x"2e00", 1285=>x"4400", 1286=>x"4000", 1287=>x"3000", 1288=>x"3900",
---- 1289=>x"5000", 1290=>x"2d00", 1291=>x"2200", 1292=>x"2c00", 1293=>x"3600", 1294=>x"3e00", 1295=>x"3800",
---- 1296=>x"4d00", 1297=>x"3c00", 1298=>x"2f00", 1299=>x"2200", 1300=>x"2200", 1301=>x"2100", 1302=>x"2900",
---- 1303=>x"4700", 1304=>x"3100", 1305=>x"5200", 1306=>x"7100", 1307=>x"3800", 1308=>x"2600", 1309=>x"2800",
---- 1310=>x"2200", 1311=>x"2400", 1312=>x"2600", 1313=>x"6b00", 1314=>x"a900", 1315=>x"6000", 1316=>x"3200",
---- 1317=>x"1f00", 1318=>x"2300", 1319=>x"2100", 1320=>x"2a00", 1321=>x"6000", 1322=>x"a500", 1323=>x"9c00",
---- 1324=>x"4100", 1325=>x"1900", 1326=>x"1a00", 1327=>x"4500", 1328=>x"3100", 1329=>x"4f00", 1330=>x"8900",
---- 1331=>x"7a00", 1332=>x"4400", 1333=>x"2500", 1334=>x"3200", 1335=>x"4d00", 1336=>x"4700", 1337=>x"4c00",
---- 1338=>x"6f00", 1339=>x"5e00", 1340=>x"3c00", 1341=>x"3e00", 1342=>x"4600", 1343=>x"2b00", 1344=>x"5e00",
---- 1345=>x"5800", 1346=>x"5900", 1347=>x"5a00", 1348=>x"3c00", 1349=>x"3400", 1350=>x"3d00", 1351=>x"2300",
---- 1352=>x"7000", 1353=>x"6c00", 1354=>x"4000", 1355=>x"4000", 1356=>x"3000", 1357=>x"1f00", 1358=>x"3600",
---- 1359=>x"4100", 1360=>x"9600", 1361=>x"5f00", 1362=>x"2d00", 1363=>x"2a00", 1364=>x"3700", 1365=>x"3a00",
---- 1366=>x"4500", 1367=>x"6400", 1368=>x"9400", 1369=>x"3600", 1370=>x"2700", 1371=>x"2c00", 1372=>x"2f00",
---- 1373=>x"6d00", 1374=>x"7200", 1375=>x"6200", 1376=>x"5e00", 1377=>x"1b00", 1378=>x"2200", 1379=>x"3200",
---- 1380=>x"6a00", 1381=>x"8b00", 1382=>x"9e00", 1383=>x"9800", 1384=>x"7b00", 1385=>x"3a00", 1386=>x"1b00",
---- 1387=>x"5200", 1388=>x"6f00", 1389=>x"7400", 1390=>x"a200", 1391=>x"c600", 1392=>x"7300", 1393=>x"6d00",
---- 1394=>x"5a00", 1395=>x"9000", 1396=>x"8800", 1397=>x"6c00", 1398=>x"9f00", 1399=>x"c200", 1400=>x"5900",
---- 1401=>x"4600", 1402=>x"8300", 1403=>x"9900", 1404=>x"8100", 1405=>x"8900", 1406=>x"b800", 1407=>x"bf00",
---- 1408=>x"3900", 1409=>x"4400", 1410=>x"7100", 1411=>x"8100", 1412=>x"7f00", 1413=>x"8900", 1414=>x"bb00",
---- 1415=>x"2400", 1416=>x"5500", 1417=>x"6b00", 1418=>x"9200", 1419=>x"9500", 1420=>x"8900", 1421=>x"8400",
---- 1422=>x"9800", 1423=>x"e200", 1424=>x"7400", 1425=>x"7e00", 1426=>x"9200", 1427=>x"9600", 1428=>x"8700",
---- 1429=>x"7a00", 1430=>x"7d00", 1431=>x"d100", 1432=>x"8100", 1433=>x"8200", 1434=>x"8f00", 1435=>x"9600",
---- 1436=>x"8000", 1437=>x"7800", 1438=>x"a100", 1439=>x"cd00", 1440=>x"8600", 1441=>x"9800", 1442=>x"8d00",
---- 1443=>x"9900", 1444=>x"7500", 1445=>x"8300", 1446=>x"d400", 1447=>x"ac00", 1448=>x"9100", 1449=>x"a700",
---- 1450=>x"9f00", 1451=>x"8f00", 1452=>x"7300", 1453=>x"8300", 1454=>x"c900", 1455=>x"9200", 1456=>x"6300",
---- 1457=>x"8000", 1458=>x"9300", 1459=>x"8700", 1460=>x"7e00", 1461=>x"8a00", 1462=>x"ca00", 1463=>x"a600",
---- 1464=>x"5f00", 1465=>x"6800", 1466=>x"7600", 1467=>x"7400", 1468=>x"7b00", 1469=>x"9f00", 1470=>x"c900",
---- 1471=>x"9600", 1472=>x"4500", 1473=>x"7200", 1474=>x"7f00", 1475=>x"6d00", 1476=>x"7100", 1477=>x"9b00",
---- 1478=>x"c900", 1479=>x"a300", 1480=>x"3200", 1481=>x"6400", 1482=>x"7b00", 1483=>x"7300", 1484=>x"8000",
---- 1485=>x"af00", 1486=>x"da00", 1487=>x"cc00", 1488=>x"5f00", 1489=>x"7900", 1490=>x"6100", 1491=>x"6000",
---- 1492=>x"7300", 1493=>x"a000", 1494=>x"d700", 1495=>x"c200", 1496=>x"6f00", 1497=>x"8c00", 1498=>x"5e00",
---- 1499=>x"4f00", 1500=>x"6f00", 1501=>x"7600", 1502=>x"c100", 1503=>x"7d00", 1504=>x"6100", 1505=>x"9600",
---- 1506=>x"6f00", 1507=>x"3a00", 1508=>x"6800", 1509=>x"7900", 1510=>x"b700", 1511=>x"6500", 1512=>x"7600",
---- 1513=>x"9300", 1514=>x"7d00", 1515=>x"5700", 1516=>x"5b00", 1517=>x"6200", 1518=>x"5700", 1519=>x"4700",
---- 1520=>x"8800", 1521=>x"9500", 1522=>x"6a00", 1523=>x"5f00", 1524=>x"6100", 1525=>x"6c00", 1526=>x"3700",
---- 1527=>x"3f00", 1528=>x"7e00", 1529=>x"9300", 1530=>x"9f00", 1531=>x"5600", 1532=>x"4800", 1533=>x"6200",
---- 1534=>x"5b00", 1535=>x"3e00", 1536=>x"7f00", 1537=>x"9600", 1538=>x"a800", 1539=>x"7c00", 1540=>x"7300",
---- 1541=>x"7b00", 1542=>x"7d00", 1543=>x"4b00", 1544=>x"8f00", 1545=>x"9d00", 1546=>x"9000", 1547=>x"8700",
---- 1548=>x"9800", 1549=>x"a700", 1550=>x"9b00", 1551=>x"7f00", 1552=>x"8200", 1553=>x"9e00", 1554=>x"9100",
---- 1555=>x"7200", 1556=>x"5100", 1557=>x"7600", 1558=>x"9600", 1559=>x"a600", 1560=>x"5800", 1561=>x"9400",
---- 1562=>x"a100", 1563=>x"8800", 1564=>x"5500", 1565=>x"3600", 1566=>x"4900", 1567=>x"9c00", 1568=>x"5b00",
---- 1569=>x"7c00", 1570=>x"9400", 1571=>x"7e00", 1572=>x"7a00", 1573=>x"6500", 1574=>x"3100", 1575=>x"6300",
---- 1576=>x"6000", 1577=>x"5c00", 1578=>x"7200", 1579=>x"7e00", 1580=>x"6000", 1581=>x"6600", 1582=>x"4a00",
---- 1583=>x"4900", 1584=>x"6900", 1585=>x"5f00", 1586=>x"5c00", 1587=>x"8200", 1588=>x"7800", 1589=>x"3e00",
---- 1590=>x"6400", 1591=>x"7f00", 1592=>x"5300", 1593=>x"6d00", 1594=>x"7000", 1595=>x"6900", 1596=>x"7300",
---- 1597=>x"6000", 1598=>x"6e00", 1599=>x"9800", 1600=>x"6300", 1601=>x"6400", 1602=>x"7600", 1603=>x"7600",
---- 1604=>x"6f00", 1605=>x"6f00", 1606=>x"7100", 1607=>x"7600", 1608=>x"6900", 1609=>x"6f00", 1610=>x"5300",
---- 1611=>x"8a00", 1612=>x"7e00", 1613=>x"8e00", 1614=>x"8200", 1615=>x"7c00", 1616=>x"7700", 1617=>x"7700",
---- 1618=>x"5b00", 1619=>x"7300", 1620=>x"9c00", 1621=>x"7a00", 1622=>x"8600", 1623=>x"7900", 1624=>x"7700",
---- 1625=>x"7a00", 1626=>x"7500", 1627=>x"8500", 1628=>x"9500", 1629=>x"8b00", 1630=>x"7f00", 1631=>x"8600",
---- 1632=>x"6000", 1633=>x"7900", 1634=>x"7d00", 1635=>x"8a00", 1636=>x"8900", 1637=>x"8b00", 1638=>x"8b00",
---- 1639=>x"9200", 1640=>x"5600", 1641=>x"5c00", 1642=>x"7000", 1643=>x"8100", 1644=>x"8700", 1645=>x"8100",
---- 1646=>x"9600", 1647=>x"9500", 1648=>x"6200", 1649=>x"5200", 1650=>x"5a00", 1651=>x"7e00", 1652=>x"9000",
---- 1653=>x"8100", 1654=>x"9000", 1655=>x"8200", 1656=>x"7400", 1657=>x"6000", 1658=>x"5100", 1659=>x"7400",
---- 1660=>x"8f00", 1661=>x"8700", 1662=>x"8500", 1663=>x"7600", 1664=>x"6700", 1665=>x"7200", 1666=>x"5400",
---- 1667=>x"6f00", 1668=>x"9300", 1669=>x"8200", 1670=>x"8300", 1671=>x"8500", 1672=>x"4b00", 1673=>x"6d00",
---- 1674=>x"5d00", 1675=>x"7100", 1676=>x"7c00", 1677=>x"8c00", 1678=>x"7300", 1679=>x"8e00", 1680=>x"3d00",
---- 1681=>x"5000", 1682=>x"5f00", 1683=>x"7500", 1684=>x"6300", 1685=>x"6400", 1686=>x"7a00", 1687=>x"7e00",
---- 1688=>x"5c00", 1689=>x"4300", 1690=>x"4d00", 1691=>x"7200", 1692=>x"5d00", 1693=>x"6f00", 1694=>x"8d00",
---- 1695=>x"6b00", 1696=>x"7600", 1697=>x"6500", 1698=>x"4300", 1699=>x"5e00", 1700=>x"5300", 1701=>x"6d00",
---- 1702=>x"8e00", 1703=>x"8300", 1704=>x"6a00", 1705=>x"6600", 1706=>x"4f00", 1707=>x"5500", 1708=>x"5100",
---- 1709=>x"5c00", 1710=>x"8f00", 1711=>x"9d00", 1712=>x"6500", 1713=>x"5700", 1714=>x"4e00", 1715=>x"5800",
---- 1716=>x"4f00", 1717=>x"5f00", 1718=>x"8a00", 1719=>x"6a00", 1720=>x"6f00", 1721=>x"5d00", 1722=>x"5700",
---- 1723=>x"4c00", 1724=>x"4700", 1725=>x"6500", 1726=>x"8500", 1727=>x"9000", 1728=>x"7700", 1729=>x"6500",
---- 1730=>x"5200", 1731=>x"4f00", 1732=>x"3d00", 1733=>x"5e00", 1734=>x"9500", 1735=>x"8700", 1736=>x"8100",
---- 1737=>x"7200", 1738=>x"3f00", 1739=>x"3b00", 1740=>x"3700", 1741=>x"5500", 1742=>x"9900", 1743=>x"8900",
---- 1744=>x"6b00", 1745=>x"8500", 1746=>x"4700", 1747=>x"3600", 1748=>x"4e00", 1749=>x"6600", 1750=>x"8f00",
---- 1751=>x"8900", 1752=>x"7200", 1753=>x"7600", 1754=>x"6900", 1755=>x"5800", 1756=>x"6100", 1757=>x"6d00",
---- 1758=>x"8b00", 1759=>x"8700", 1760=>x"4e00", 1761=>x"5400", 1762=>x"7000", 1763=>x"7e00", 1764=>x"7a00",
---- 1765=>x"7900", 1766=>x"8400", 1767=>x"8f00", 1768=>x"2c00", 1769=>x"3500", 1770=>x"4a00", 1771=>x"7500",
---- 1772=>x"8b00", 1773=>x"8600", 1774=>x"7900", 1775=>x"8800", 1776=>x"2200", 1777=>x"2c00", 1778=>x"3f00",
---- 1779=>x"6e00", 1780=>x"9100", 1781=>x"8800", 1782=>x"7800", 1783=>x"8400", 1784=>x"2700", 1785=>x"2d00",
---- 1786=>x"4400", 1787=>x"6700", 1788=>x"8500", 1789=>x"6300", 1790=>x"8900", 1791=>x"7500", 1792=>x"5100",
---- 1793=>x"3d00", 1794=>x"5000", 1795=>x"6100", 1796=>x"7900", 1797=>x"6800", 1798=>x"7800", 1799=>x"7c00",
---- 1800=>x"5500", 1801=>x"5b00", 1802=>x"4e00", 1803=>x"6200", 1804=>x"6100", 1805=>x"7800", 1806=>x"7300",
---- 1807=>x"6a00", 1808=>x"2a00", 1809=>x"5e00", 1810=>x"6900", 1811=>x"5000", 1812=>x"5300", 1813=>x"6600",
---- 1814=>x"7300", 1815=>x"7400", 1816=>x"2e00", 1817=>x"2800", 1818=>x"7400", 1819=>x"9a00", 1820=>x"8300",
---- 1821=>x"8100", 1822=>x"7700", 1823=>x"7c00", 1824=>x"5600", 1825=>x"2100", 1826=>x"3200", 1827=>x"6d00",
---- 1828=>x"6000", 1829=>x"7c00", 1830=>x"7900", 1831=>x"7700", 1832=>x"6100", 1833=>x"4300", 1834=>x"3100",
---- 1835=>x"2700", 1836=>x"3500", 1837=>x"3b00", 1838=>x"5b00", 1839=>x"8b00", 1840=>x"7800", 1841=>x"4d00",
---- 1842=>x"4700", 1843=>x"3800", 1844=>x"3700", 1845=>x"2800", 1846=>x"2800", 1847=>x"6600", 1848=>x"8000",
---- 1849=>x"7600", 1850=>x"3a00", 1851=>x"4400", 1852=>x"3500", 1853=>x"2500", 1854=>x"2e00", 1855=>x"4100",
---- 1856=>x"7c00", 1857=>x"9100", 1858=>x"5a00", 1859=>x"2a00", 1860=>x"4300", 1861=>x"4700", 1862=>x"2d00",
---- 1863=>x"3b00", 1864=>x"8a00", 1865=>x"8000", 1866=>x"9600", 1867=>x"5400", 1868=>x"3300", 1869=>x"4900",
---- 1870=>x"4000", 1871=>x"4000", 1872=>x"6600", 1873=>x"7600", 1874=>x"8900", 1875=>x"9600", 1876=>x"6700",
---- 1877=>x"3400", 1878=>x"3d00", 1879=>x"5b00", 1880=>x"9c00", 1881=>x"7400", 1882=>x"7900", 1883=>x"8500",
---- 1884=>x"9300", 1885=>x"6b00", 1886=>x"6500", 1887=>x"6b00", 1888=>x"5e00", 1889=>x"6c00", 1890=>x"8600",
---- 1891=>x"8f00", 1892=>x"7100", 1893=>x"8500", 1894=>x"7b00", 1895=>x"6600", 1896=>x"3000", 1897=>x"5200",
---- 1898=>x"7000", 1899=>x"9d00", 1900=>x"8b00", 1901=>x"7a00", 1902=>x"8200", 1903=>x"5400", 1904=>x"2c00",
---- 1905=>x"2700", 1906=>x"4d00", 1907=>x"7d00", 1908=>x"8900", 1909=>x"8d00", 1910=>x"8600", 1911=>x"6400",
---- 1912=>x"2e00", 1913=>x"2b00", 1914=>x"3900", 1915=>x"5200", 1916=>x"7500", 1917=>x"7200", 1918=>x"a700",
---- 1919=>x"8b00", 1920=>x"3600", 1921=>x"4100", 1922=>x"3c00", 1923=>x"4300", 1924=>x"4a00", 1925=>x"5400",
---- 1926=>x"7600", 1927=>x"8a00", 1928=>x"3000", 1929=>x"4c00", 1930=>x"5600", 1931=>x"3500", 1932=>x"4e00",
---- 1933=>x"4b00", 1934=>x"5c00", 1935=>x"5000", 1936=>x"3200", 1937=>x"4000", 1938=>x"6700", 1939=>x"3f00",
---- 1940=>x"4700", 1941=>x"7800", 1942=>x"8100", 1943=>x"4200", 1944=>x"3300", 1945=>x"4300", 1946=>x"3e00",
---- 1947=>x"5200", 1948=>x"4800", 1949=>x"6400", 1950=>x"9700", 1951=>x"6600", 1952=>x"4800", 1953=>x"3800",
---- 1954=>x"3b00", 1955=>x"4b00", 1956=>x"5000", 1957=>x"4a00", 1958=>x"8a00", 1959=>x"8200", 1960=>x"7b00",
---- 1961=>x"3500", 1962=>x"3700", 1963=>x"3a00", 1964=>x"5400", 1965=>x"6600", 1966=>x"7400", 1967=>x"9d00",
---- 1968=>x"6e00", 1969=>x"5d00", 1970=>x"4000", 1971=>x"3800", 1972=>x"4d00", 1973=>x"7300", 1974=>x"6e00",
---- 1975=>x"8500", 1976=>x"4600", 1977=>x"6a00", 1978=>x"4c00", 1979=>x"4200", 1980=>x"3d00", 1981=>x"7100",
---- 1982=>x"7800", 1983=>x"6300", 1984=>x"4800", 1985=>x"5200", 1986=>x"6600", 1987=>x"3c00", 1988=>x"4400",
---- 1989=>x"5f00", 1990=>x"7100", 1991=>x"7500", 1992=>x"d200", 1993=>x"5200", 1994=>x"7200", 1995=>x"4a00",
---- 1996=>x"2a00", 1997=>x"4c00", 1998=>x"6c00", 1999=>x"7800", 2000=>x"2000", 2001=>x"4400", 2002=>x"5b00",
---- 2003=>x"7c00", 2004=>x"3300", 2005=>x"2900", 2006=>x"4c00", 2007=>x"5d00", 2008=>x"1e00", 2009=>x"3800",
---- 2010=>x"4900", 2011=>x"6900", 2012=>x"6b00", 2013=>x"2400", 2014=>x"3c00", 2015=>x"4a00", 2016=>x"3d00",
---- 2017=>x"2a00", 2018=>x"4e00", 2019=>x"4600", 2020=>x"6800", 2021=>x"4200", 2022=>x"3800", 2023=>x"4c00",
---- 2024=>x"4000", 2025=>x"3a00", 2026=>x"4500", 2027=>x"5600", 2028=>x"4400", 2029=>x"4a00", 2030=>x"2e00",
---- 2031=>x"4300", 2032=>x"2500", 2033=>x"3000", 2034=>x"3f00", 2035=>x"5800", 2036=>x"4900", 2037=>x"3d00",
---- 2038=>x"3300", 2039=>x"2e00", 2040=>x"2d00", 2041=>x"2e00", 2042=>x"3000", 2043=>x"4200", 2044=>x"4e00",
---- 2045=>x"4700", 2046=>x"3f00", 2047=>x"2c00"),
---- 10 => (0=>x"8100", 1=>x"8600", 2=>x"8500", 3=>x"8600", 4=>x"8600", 5=>x"8500", 6=>x"8600", 7=>x"8600",
---- 8=>x"8200", 9=>x"8400", 10=>x"8500", 11=>x"8600", 12=>x"8500", 13=>x"8600", 14=>x"8600",
---- 15=>x"8400", 16=>x"8300", 17=>x"7900", 18=>x"8600", 19=>x"8700", 20=>x"8600", 21=>x"8400",
---- 22=>x"8600", 23=>x"8500", 24=>x"8300", 25=>x"8500", 26=>x"8700", 27=>x"8700", 28=>x"8500",
---- 29=>x"8400", 30=>x"8500", 31=>x"7800", 32=>x"8400", 33=>x"8300", 34=>x"8300", 35=>x"8500",
---- 36=>x"8500", 37=>x"8500", 38=>x"8600", 39=>x"8500", 40=>x"8200", 41=>x"8300", 42=>x"7b00",
---- 43=>x"8600", 44=>x"8400", 45=>x"8400", 46=>x"8500", 47=>x"8500", 48=>x"8000", 49=>x"8300",
---- 50=>x"8500", 51=>x"8400", 52=>x"8400", 53=>x"8300", 54=>x"8400", 55=>x"8400", 56=>x"8100",
---- 57=>x"8300", 58=>x"8000", 59=>x"8200", 60=>x"8100", 61=>x"8500", 62=>x"8600", 63=>x"8500",
---- 64=>x"8400", 65=>x"8600", 66=>x"8700", 67=>x"8400", 68=>x"8300", 69=>x"8700", 70=>x"8400",
---- 71=>x"8600", 72=>x"8300", 73=>x"8300", 74=>x"8600", 75=>x"8200", 76=>x"8300", 77=>x"8400",
---- 78=>x"8600", 79=>x"8500", 80=>x"8200", 81=>x"8000", 82=>x"8300", 83=>x"8300", 84=>x"8300",
---- 85=>x"8100", 86=>x"8400", 87=>x"8400", 88=>x"8100", 89=>x"8300", 90=>x"8400", 91=>x"8400",
---- 92=>x"8100", 93=>x"8300", 94=>x"8300", 95=>x"8400", 96=>x"8100", 97=>x"8100", 98=>x"8300",
---- 99=>x"8200", 100=>x"8000", 101=>x"8300", 102=>x"8600", 103=>x"8500", 104=>x"8100", 105=>x"8300",
---- 106=>x"8100", 107=>x"8000", 108=>x"7e00", 109=>x"8100", 110=>x"8000", 111=>x"8200", 112=>x"8200",
---- 113=>x"8200", 114=>x"8100", 115=>x"8400", 116=>x"8100", 117=>x"8100", 118=>x"8000", 119=>x"8400",
---- 120=>x"8000", 121=>x"8300", 122=>x"8200", 123=>x"8100", 124=>x"8200", 125=>x"8200", 126=>x"8000",
---- 127=>x"8300", 128=>x"8400", 129=>x"8200", 130=>x"8300", 131=>x"8300", 132=>x"8300", 133=>x"7d00",
---- 134=>x"8300", 135=>x"8200", 136=>x"8400", 137=>x"8200", 138=>x"8100", 139=>x"7f00", 140=>x"8100",
---- 141=>x"8300", 142=>x"8400", 143=>x"7f00", 144=>x"8000", 145=>x"7d00", 146=>x"8100", 147=>x"7f00",
---- 148=>x"8000", 149=>x"7f00", 150=>x"7e00", 151=>x"8000", 152=>x"8200", 153=>x"7f00", 154=>x"8200",
---- 155=>x"7f00", 156=>x"7c00", 157=>x"7d00", 158=>x"8000", 159=>x"8000", 160=>x"8300", 161=>x"8100",
---- 162=>x"8100", 163=>x"8000", 164=>x"7e00", 165=>x"8100", 166=>x"8200", 167=>x"8000", 168=>x"8000",
---- 169=>x"7d00", 170=>x"7f00", 171=>x"8000", 172=>x"7c00", 173=>x"8100", 174=>x"8000", 175=>x"7f00",
---- 176=>x"8000", 177=>x"7f00", 178=>x"7d00", 179=>x"7a00", 180=>x"7e00", 181=>x"8100", 182=>x"8100",
---- 183=>x"8000", 184=>x"8200", 185=>x"8000", 186=>x"7d00", 187=>x"7d00", 188=>x"7f00", 189=>x"8900",
---- 190=>x"8500", 191=>x"8000", 192=>x"8100", 193=>x"7f00", 194=>x"7e00", 195=>x"8000", 196=>x"7f00",
---- 197=>x"7f00", 198=>x"8000", 199=>x"8200", 200=>x"8200", 201=>x"7f00", 202=>x"7f00", 203=>x"7f00",
---- 204=>x"7f00", 205=>x"7f00", 206=>x"8100", 207=>x"8200", 208=>x"8200", 209=>x"8300", 210=>x"8000",
---- 211=>x"7f00", 212=>x"8000", 213=>x"8100", 214=>x"7f00", 215=>x"8000", 216=>x"8000", 217=>x"7e00",
---- 218=>x"7f00", 219=>x"7c00", 220=>x"7e00", 221=>x"7f00", 222=>x"7f00", 223=>x"7f00", 224=>x"8000",
---- 225=>x"7e00", 226=>x"7c00", 227=>x"7d00", 228=>x"7c00", 229=>x"7d00", 230=>x"8000", 231=>x"8200",
---- 232=>x"7d00", 233=>x"7a00", 234=>x"7b00", 235=>x"7a00", 236=>x"7e00", 237=>x"9100", 238=>x"9100",
---- 239=>x"9400", 240=>x"7900", 241=>x"7d00", 242=>x"a300", 243=>x"9900", 244=>x"9300", 245=>x"9f00",
---- 246=>x"9400", 247=>x"8e00", 248=>x"8600", 249=>x"8000", 250=>x"8d00", 251=>x"8d00", 252=>x"8d00",
---- 253=>x"8500", 254=>x"8200", 255=>x"7b00", 256=>x"9000", 257=>x"6f00", 258=>x"7b00", 259=>x"7b00",
---- 260=>x"7e00", 261=>x"7c00", 262=>x"7900", 263=>x"7700", 264=>x"5b00", 265=>x"6700", 266=>x"7b00",
---- 267=>x"7900", 268=>x"7800", 269=>x"7700", 270=>x"7b00", 271=>x"7600", 272=>x"6000", 273=>x"6e00",
---- 274=>x"7600", 275=>x"7600", 276=>x"7d00", 277=>x"7700", 278=>x"7900", 279=>x"7900", 280=>x"7300",
---- 281=>x"7000", 282=>x"7400", 283=>x"7700", 284=>x"7a00", 285=>x"7500", 286=>x"7700", 287=>x"7b00",
---- 288=>x"7200", 289=>x"7500", 290=>x"7600", 291=>x"7400", 292=>x"6e00", 293=>x"7000", 294=>x"7900",
---- 295=>x"7600", 296=>x"7500", 297=>x"7000", 298=>x"6f00", 299=>x"6d00", 300=>x"6e00", 301=>x"7200",
---- 302=>x"7400", 303=>x"7600", 304=>x"6c00", 305=>x"6e00", 306=>x"6900", 307=>x"6c00", 308=>x"7100",
---- 309=>x"7700", 310=>x"7800", 311=>x"7600", 312=>x"6a00", 313=>x"9400", 314=>x"6c00", 315=>x"7000",
---- 316=>x"7600", 317=>x"7800", 318=>x"7400", 319=>x"7400", 320=>x"6a00", 321=>x"6d00", 322=>x"6f00",
---- 323=>x"7100", 324=>x"7900", 325=>x"7500", 326=>x"7200", 327=>x"7400", 328=>x"7100", 329=>x"7100",
---- 330=>x"7500", 331=>x"7700", 332=>x"7a00", 333=>x"7500", 334=>x"7200", 335=>x"7c00", 336=>x"6f00",
---- 337=>x"8900", 338=>x"7800", 339=>x"7600", 340=>x"7400", 341=>x"7600", 342=>x"7d00", 343=>x"7800",
---- 344=>x"7300", 345=>x"7700", 346=>x"7200", 347=>x"7400", 348=>x"7a00", 349=>x"7b00", 350=>x"7a00",
---- 351=>x"7700", 352=>x"7300", 353=>x"7100", 354=>x"6f00", 355=>x"7a00", 356=>x"7b00", 357=>x"7500",
---- 358=>x"7200", 359=>x"7b00", 360=>x"6f00", 361=>x"7300", 362=>x"7d00", 363=>x"7500", 364=>x"7500",
---- 365=>x"7200", 366=>x"7200", 367=>x"7a00", 368=>x"7200", 369=>x"7900", 370=>x"7800", 371=>x"7600",
---- 372=>x"7700", 373=>x"7600", 374=>x"7600", 375=>x"7500", 376=>x"7700", 377=>x"7500", 378=>x"7300",
---- 379=>x"8700", 380=>x"7100", 381=>x"6f00", 382=>x"6e00", 383=>x"6a00", 384=>x"7800", 385=>x"7500",
---- 386=>x"7700", 387=>x"7000", 388=>x"6e00", 389=>x"7100", 390=>x"6e00", 391=>x"7300", 392=>x"7400",
---- 393=>x"7600", 394=>x"6f00", 395=>x"7400", 396=>x"7500", 397=>x"7900", 398=>x"7800", 399=>x"7b00",
---- 400=>x"7600", 401=>x"7700", 402=>x"7100", 403=>x"7800", 404=>x"7900", 405=>x"7a00", 406=>x"7600",
---- 407=>x"7600", 408=>x"7100", 409=>x"7000", 410=>x"7200", 411=>x"7400", 412=>x"7100", 413=>x"7600",
---- 414=>x"7700", 415=>x"7700", 416=>x"7400", 417=>x"7200", 418=>x"8d00", 419=>x"7100", 420=>x"7500",
---- 421=>x"7500", 422=>x"7400", 423=>x"7b00", 424=>x"7200", 425=>x"7200", 426=>x"6f00", 427=>x"6f00",
---- 428=>x"7300", 429=>x"8500", 430=>x"7b00", 431=>x"7b00", 432=>x"6f00", 433=>x"7100", 434=>x"7200",
---- 435=>x"7500", 436=>x"7800", 437=>x"7c00", 438=>x"8000", 439=>x"7600", 440=>x"7400", 441=>x"7900",
---- 442=>x"7700", 443=>x"7a00", 444=>x"7a00", 445=>x"7a00", 446=>x"7d00", 447=>x"7f00", 448=>x"7600",
---- 449=>x"7800", 450=>x"7b00", 451=>x"7600", 452=>x"7700", 453=>x"7d00", 454=>x"7f00", 455=>x"7b00",
---- 456=>x"6d00", 457=>x"7800", 458=>x"7700", 459=>x"7800", 460=>x"7d00", 461=>x"7c00", 462=>x"8200",
---- 463=>x"8000", 464=>x"7100", 465=>x"7700", 466=>x"7500", 467=>x"7500", 468=>x"7d00", 469=>x"8200",
---- 470=>x"8100", 471=>x"8400", 472=>x"7300", 473=>x"7c00", 474=>x"8900", 475=>x"7500", 476=>x"7d00",
---- 477=>x"8000", 478=>x"8400", 479=>x"7f00", 480=>x"7600", 481=>x"7800", 482=>x"7700", 483=>x"7900",
---- 484=>x"8200", 485=>x"7c00", 486=>x"8600", 487=>x"8300", 488=>x"7800", 489=>x"7000", 490=>x"7600",
---- 491=>x"7e00", 492=>x"8400", 493=>x"8500", 494=>x"8100", 495=>x"7600", 496=>x"7000", 497=>x"7700",
---- 498=>x"8000", 499=>x"8500", 500=>x"8400", 501=>x"7d00", 502=>x"7900", 503=>x"7a00", 504=>x"7d00",
---- 505=>x"8200", 506=>x"7e00", 507=>x"8200", 508=>x"7e00", 509=>x"7800", 510=>x"7800", 511=>x"7400",
---- 512=>x"7b00", 513=>x"7f00", 514=>x"7800", 515=>x"7900", 516=>x"7d00", 517=>x"7100", 518=>x"7100",
---- 519=>x"7b00", 520=>x"7900", 521=>x"7900", 522=>x"7c00", 523=>x"7a00", 524=>x"7600", 525=>x"7700",
---- 526=>x"7900", 527=>x"8600", 528=>x"7d00", 529=>x"7d00", 530=>x"6d00", 531=>x"7200", 532=>x"7b00",
---- 533=>x"8300", 534=>x"7800", 535=>x"7e00", 536=>x"7a00", 537=>x"6a00", 538=>x"7400", 539=>x"8000",
---- 540=>x"7a00", 541=>x"7b00", 542=>x"8100", 543=>x"7d00", 544=>x"7200", 545=>x"7500", 546=>x"7a00",
---- 547=>x"7a00", 548=>x"8100", 549=>x"8100", 550=>x"8200", 551=>x"7f00", 552=>x"7100", 553=>x"7100",
---- 554=>x"7c00", 555=>x"7d00", 556=>x"8100", 557=>x"8000", 558=>x"7300", 559=>x"7000", 560=>x"6800",
---- 561=>x"7600", 562=>x"7800", 563=>x"7c00", 564=>x"7d00", 565=>x"7000", 566=>x"6d00", 567=>x"7a00",
---- 568=>x"7700", 569=>x"7a00", 570=>x"7c00", 571=>x"7300", 572=>x"6e00", 573=>x"7400", 574=>x"7d00",
---- 575=>x"7e00", 576=>x"7300", 577=>x"7b00", 578=>x"7100", 579=>x"6d00", 580=>x"7900", 581=>x"8100",
---- 582=>x"8200", 583=>x"7a00", 584=>x"7800", 585=>x"7400", 586=>x"6f00", 587=>x"7c00", 588=>x"8000",
---- 589=>x"7d00", 590=>x"7800", 591=>x"6b00", 592=>x"7600", 593=>x"7e00", 594=>x"7a00", 595=>x"7c00",
---- 596=>x"8200", 597=>x"7800", 598=>x"6500", 599=>x"7300", 600=>x"7900", 601=>x"7700", 602=>x"7a00",
---- 603=>x"7d00", 604=>x"7b00", 605=>x"7000", 606=>x"7000", 607=>x"8a00", 608=>x"7900", 609=>x"7400",
---- 610=>x"7900", 611=>x"7400", 612=>x"6c00", 613=>x"7400", 614=>x"8e00", 615=>x"8900", 616=>x"8100",
---- 617=>x"7100", 618=>x"6300", 619=>x"6600", 620=>x"7800", 621=>x"9000", 622=>x"8c00", 623=>x"8e00",
---- 624=>x"7800", 625=>x"6c00", 626=>x"6100", 627=>x"7200", 628=>x"9000", 629=>x"9400", 630=>x"8a00",
---- 631=>x"8800", 632=>x"7400", 633=>x"6700", 634=>x"7400", 635=>x"8b00", 636=>x"8e00", 637=>x"8d00",
---- 638=>x"8e00", 639=>x"8300", 640=>x"6000", 641=>x"7800", 642=>x"9200", 643=>x"8b00", 644=>x"8600",
---- 645=>x"8a00", 646=>x"8700", 647=>x"8700", 648=>x"6f00", 649=>x"9100", 650=>x"9000", 651=>x"8b00",
---- 652=>x"8a00", 653=>x"8000", 654=>x"8400", 655=>x"8e00", 656=>x"8f00", 657=>x"9000", 658=>x"8c00",
---- 659=>x"8700", 660=>x"8600", 661=>x"7e00", 662=>x"8600", 663=>x"8f00", 664=>x"8a00", 665=>x"8e00",
---- 666=>x"8800", 667=>x"8600", 668=>x"7c00", 669=>x"8d00", 670=>x"8400", 671=>x"8f00", 672=>x"7900",
---- 673=>x"8700", 674=>x"8700", 675=>x"7f00", 676=>x"8e00", 677=>x"8b00", 678=>x"7000", 679=>x"7700",
---- 680=>x"8300", 681=>x"7b00", 682=>x"8400", 683=>x"8900", 684=>x"8800", 685=>x"6e00", 686=>x"7e00",
---- 687=>x"7b00", 688=>x"8500", 689=>x"7c00", 690=>x"8800", 691=>x"8d00", 692=>x"6c00", 693=>x"7500",
---- 694=>x"7d00", 695=>x"8100", 696=>x"7d00", 697=>x"8800", 698=>x"8700", 699=>x"7200", 700=>x"6c00",
---- 701=>x"7e00", 702=>x"7f00", 703=>x"8f00", 704=>x"7f00", 705=>x"8900", 706=>x"7000", 707=>x"6f00",
---- 708=>x"7600", 709=>x"8200", 710=>x"9000", 711=>x"8c00", 712=>x"8600", 713=>x"6e00", 714=>x"6800",
---- 715=>x"7800", 716=>x"7e00", 717=>x"8c00", 718=>x"8d00", 719=>x"8900", 720=>x"6d00", 721=>x"6200",
---- 722=>x"7700", 723=>x"8500", 724=>x"8d00", 725=>x"8a00", 726=>x"8600", 727=>x"8500", 728=>x"6300",
---- 729=>x"7100", 730=>x"7700", 731=>x"8800", 732=>x"8b00", 733=>x"8700", 734=>x"8600", 735=>x"8600",
---- 736=>x"7300", 737=>x"7700", 738=>x"8300", 739=>x"8c00", 740=>x"8600", 741=>x"8700", 742=>x"8600",
---- 743=>x"8a00", 744=>x"7400", 745=>x"8000", 746=>x"8800", 747=>x"8b00", 748=>x"7500", 749=>x"8800",
---- 750=>x"8600", 751=>x"7b00", 752=>x"7e00", 753=>x"8600", 754=>x"8900", 755=>x"8500", 756=>x"8a00",
---- 757=>x"8900", 758=>x"7800", 759=>x"7300", 760=>x"8900", 761=>x"8400", 762=>x"8500", 763=>x"8900",
---- 764=>x"8400", 765=>x"7f00", 766=>x"7000", 767=>x"7f00", 768=>x"8700", 769=>x"8800", 770=>x"8500",
---- 771=>x"8900", 772=>x"7700", 773=>x"6d00", 774=>x"7b00", 775=>x"8100", 776=>x"8700", 777=>x"8600",
---- 778=>x"8500", 779=>x"7900", 780=>x"6a00", 781=>x"7700", 782=>x"7f00", 783=>x"7d00", 784=>x"8800",
---- 785=>x"8700", 786=>x"7200", 787=>x"6000", 788=>x"7000", 789=>x"7d00", 790=>x"7f00", 791=>x"7f00",
---- 792=>x"8600", 793=>x"8300", 794=>x"6b00", 795=>x"7400", 796=>x"7b00", 797=>x"7d00", 798=>x"8000",
---- 799=>x"7f00", 800=>x"7c00", 801=>x"6900", 802=>x"7300", 803=>x"8200", 804=>x"7d00", 805=>x"8000",
---- 806=>x"7b00", 807=>x"7800", 808=>x"7200", 809=>x"6900", 810=>x"7c00", 811=>x"7f00", 812=>x"8000",
---- 813=>x"7c00", 814=>x"7a00", 815=>x"7800", 816=>x"6d00", 817=>x"7900", 818=>x"7f00", 819=>x"8500",
---- 820=>x"8200", 821=>x"7d00", 822=>x"7a00", 823=>x"7a00", 824=>x"7500", 825=>x"7c00", 826=>x"8200",
---- 827=>x"8000", 828=>x"8500", 829=>x"8700", 830=>x"7e00", 831=>x"8100", 832=>x"8100", 833=>x"7e00",
---- 834=>x"8500", 835=>x"7e00", 836=>x"7d00", 837=>x"8100", 838=>x"7500", 839=>x"7d00", 840=>x"7f00",
---- 841=>x"8100", 842=>x"8300", 843=>x"7600", 844=>x"7300", 845=>x"6a00", 846=>x"7100", 847=>x"7d00",
---- 848=>x"8000", 849=>x"8100", 850=>x"7800", 851=>x"7000", 852=>x"6b00", 853=>x"7a00", 854=>x"8600",
---- 855=>x"8700", 856=>x"7b00", 857=>x"7500", 858=>x"7000", 859=>x"7c00", 860=>x"8200", 861=>x"8d00",
---- 862=>x"8500", 863=>x"7f00", 864=>x"6a00", 865=>x"6b00", 866=>x"7b00", 867=>x"8600", 868=>x"8b00",
---- 869=>x"8600", 870=>x"8600", 871=>x"8300", 872=>x"6700", 873=>x"7400", 874=>x"8800", 875=>x"8900",
---- 876=>x"8500", 877=>x"8300", 878=>x"7d00", 879=>x"7900", 880=>x"7800", 881=>x"8100", 882=>x"7e00",
---- 883=>x"8500", 884=>x"8100", 885=>x"8200", 886=>x"7500", 887=>x"7b00", 888=>x"8000", 889=>x"8200",
---- 890=>x"8300", 891=>x"6d00", 892=>x"7000", 893=>x"7900", 894=>x"7100", 895=>x"7200", 896=>x"7800",
---- 897=>x"7900", 898=>x"7d00", 899=>x"6500", 900=>x"5000", 901=>x"5f00", 902=>x"5a00", 903=>x"4b00",
---- 904=>x"8300", 905=>x"7900", 906=>x"5c00", 907=>x"5d00", 908=>x"4600", 909=>x"4500", 910=>x"5500",
---- 911=>x"3c00", 912=>x"8500", 913=>x"8900", 914=>x"7900", 915=>x"7000", 916=>x"6900", 917=>x"5900",
---- 918=>x"4700", 919=>x"2e00", 920=>x"8300", 921=>x"8000", 922=>x"6d00", 923=>x"6700", 924=>x"5700",
---- 925=>x"4000", 926=>x"3400", 927=>x"3700", 928=>x"8100", 929=>x"6900", 930=>x"6200", 931=>x"5a00",
---- 932=>x"3a00", 933=>x"3000", 934=>x"3800", 935=>x"5300", 936=>x"7900", 937=>x"6200", 938=>x"4400",
---- 939=>x"3100", 940=>x"3400", 941=>x"3400", 942=>x"6000", 943=>x"5d00", 944=>x"6300", 945=>x"4600",
---- 946=>x"2e00", 947=>x"4300", 948=>x"3400", 949=>x"2200", 950=>x"4d00", 951=>x"5200", 952=>x"5500",
---- 953=>x"3100", 954=>x"3800", 955=>x"5200", 956=>x"2700", 957=>x"1e00", 958=>x"5100", 959=>x"5300",
---- 960=>x"5000", 961=>x"2c00", 962=>x"5700", 963=>x"5300", 964=>x"2200", 965=>x"1f00", 966=>x"5700",
---- 967=>x"6300", 968=>x"2d00", 969=>x"3800", 970=>x"6400", 971=>x"4900", 972=>x"1f00", 973=>x"2100",
---- 974=>x"5300", 975=>x"7200", 976=>x"3700", 977=>x"5200", 978=>x"6400", 979=>x"3100", 980=>x"2200",
---- 981=>x"2c00", 982=>x"6200", 983=>x"6b00", 984=>x"5000", 985=>x"5b00", 986=>x"5700", 987=>x"2400",
---- 988=>x"2700", 989=>x"3b00", 990=>x"8000", 991=>x"6100", 992=>x"5200", 993=>x"7000", 994=>x"4100",
---- 995=>x"2500", 996=>x"2e00", 997=>x"4f00", 998=>x"7e00", 999=>x"6800", 1000=>x"5e00", 1001=>x"5300",
---- 1002=>x"d600", 1003=>x"2b00", 1004=>x"4800", 1005=>x"5c00", 1006=>x"5900", 1007=>x"7000", 1008=>x"5800",
---- 1009=>x"3000", 1010=>x"2b00", 1011=>x"3e00", 1012=>x"6c00", 1013=>x"4500", 1014=>x"3800", 1015=>x"7f00",
---- 1016=>x"5f00", 1017=>x"3d00", 1018=>x"3f00", 1019=>x"6200", 1020=>x"6500", 1021=>x"2200", 1022=>x"2800",
---- 1023=>x"6e00", 1024=>x"3700", 1025=>x"4f00", 1026=>x"4d00", 1027=>x"6400", 1028=>x"5800", 1029=>x"1c00",
---- 1030=>x"2400", 1031=>x"4e00", 1032=>x"3100", 1033=>x"5700", 1034=>x"5200", 1035=>x"6800", 1036=>x"5100",
---- 1037=>x"2200", 1038=>x"2c00", 1039=>x"4b00", 1040=>x"4800", 1041=>x"5b00", 1042=>x"4f00", 1043=>x"7b00",
---- 1044=>x"5300", 1045=>x"2100", 1046=>x"2d00", 1047=>x"4b00", 1048=>x"5800", 1049=>x"4f00", 1050=>x"5b00",
---- 1051=>x"8f00", 1052=>x"4700", 1053=>x"2000", 1054=>x"2e00", 1055=>x"4900", 1056=>x"6b00", 1057=>x"6100",
---- 1058=>x"6800", 1059=>x"7400", 1060=>x"3200", 1061=>x"d900", 1062=>x"2e00", 1063=>x"3a00", 1064=>x"7700",
---- 1065=>x"5b00", 1066=>x"6300", 1067=>x"6600", 1068=>x"3100", 1069=>x"2f00", 1070=>x"3000", 1071=>x"2b00",
---- 1072=>x"7700", 1073=>x"4f00", 1074=>x"7300", 1075=>x"7000", 1076=>x"2e00", 1077=>x"3000", 1078=>x"2d00",
---- 1079=>x"2e00", 1080=>x"8300", 1081=>x"5b00", 1082=>x"7c00", 1083=>x"7600", 1084=>x"2b00", 1085=>x"2900",
---- 1086=>x"3300", 1087=>x"2f00", 1088=>x"7700", 1089=>x"4d00", 1090=>x"7300", 1091=>x"8000", 1092=>x"3300",
---- 1093=>x"2e00", 1094=>x"3500", 1095=>x"2a00", 1096=>x"8200", 1097=>x"4200", 1098=>x"7700", 1099=>x"8a00",
---- 1100=>x"5700", 1101=>x"3f00", 1102=>x"3300", 1103=>x"2c00", 1104=>x"8c00", 1105=>x"5900", 1106=>x"8500",
---- 1107=>x"8400", 1108=>x"6000", 1109=>x"3b00", 1110=>x"5300", 1111=>x"3300", 1112=>x"7a00", 1113=>x"6b00",
---- 1114=>x"8200", 1115=>x"6a00", 1116=>x"5600", 1117=>x"7b00", 1118=>x"5000", 1119=>x"2100", 1120=>x"6500",
---- 1121=>x"7900", 1122=>x"7f00", 1123=>x"7600", 1124=>x"8700", 1125=>x"6900", 1126=>x"2100", 1127=>x"2b00",
---- 1128=>x"4700", 1129=>x"6d00", 1130=>x"7700", 1131=>x"8900", 1132=>x"8000", 1133=>x"4e00", 1134=>x"3c00",
---- 1135=>x"3c00", 1136=>x"5d00", 1137=>x"6400", 1138=>x"5800", 1139=>x"7700", 1140=>x"4500", 1141=>x"5e00",
---- 1142=>x"4a00", 1143=>x"3e00", 1144=>x"8300", 1145=>x"5200", 1146=>x"4800", 1147=>x"5400", 1148=>x"7400",
---- 1149=>x"7400", 1150=>x"2100", 1151=>x"2a00", 1152=>x"7a00", 1153=>x"5400", 1154=>x"5800", 1155=>x"8500",
---- 1156=>x"9e00", 1157=>x"4300", 1158=>x"3200", 1159=>x"3600", 1160=>x"a600", 1161=>x"8100", 1162=>x"a000",
---- 1163=>x"9200", 1164=>x"4e00", 1165=>x"5900", 1166=>x"5f00", 1167=>x"4e00", 1168=>x"7900", 1169=>x"6000",
---- 1170=>x"4d00", 1171=>x"3500", 1172=>x"3600", 1173=>x"8300", 1174=>x"8300", 1175=>x"6700", 1176=>x"6d00",
---- 1177=>x"3800", 1178=>x"1a00", 1179=>x"2500", 1180=>x"4700", 1181=>x"7c00", 1182=>x"8c00", 1183=>x"7300",
---- 1184=>x"4e00", 1185=>x"3300", 1186=>x"2300", 1187=>x"2400", 1188=>x"5100", 1189=>x"7500", 1190=>x"8e00",
---- 1191=>x"6b00", 1192=>x"4c00", 1193=>x"c200", 1194=>x"2100", 1195=>x"2200", 1196=>x"4d00", 1197=>x"7700",
---- 1198=>x"8800", 1199=>x"8700", 1200=>x"4400", 1201=>x"4100", 1202=>x"1d00", 1203=>x"3200", 1204=>x"5600",
---- 1205=>x"7500", 1206=>x"6f00", 1207=>x"7000", 1208=>x"2700", 1209=>x"3e00", 1210=>x"2a00", 1211=>x"2a00",
---- 1212=>x"5000", 1213=>x"7600", 1214=>x"5d00", 1215=>x"6600", 1216=>x"2d00", 1217=>x"3b00", 1218=>x"2d00",
---- 1219=>x"2f00", 1220=>x"5600", 1221=>x"7b00", 1222=>x"7e00", 1223=>x"4e00", 1224=>x"4d00", 1225=>x"3900",
---- 1226=>x"3900", 1227=>x"4f00", 1228=>x"5f00", 1229=>x"9300", 1230=>x"9e00", 1231=>x"6100", 1232=>x"4e00",
---- 1233=>x"3100", 1234=>x"4900", 1235=>x"5c00", 1236=>x"7900", 1237=>x"aa00", 1238=>x"b600", 1239=>x"8400",
---- 1240=>x"3d00", 1241=>x"3a00", 1242=>x"5000", 1243=>x"7400", 1244=>x"7400", 1245=>x"a400", 1246=>x"c900",
---- 1247=>x"9c00", 1248=>x"3e00", 1249=>x"6c00", 1250=>x"8500", 1251=>x"7400", 1252=>x"5800", 1253=>x"5300",
---- 1254=>x"9300", 1255=>x"8200", 1256=>x"5400", 1257=>x"8b00", 1258=>x"7b00", 1259=>x"5b00", 1260=>x"4500",
---- 1261=>x"4900", 1262=>x"5b00", 1263=>x"3a00", 1264=>x"5600", 1265=>x"9200", 1266=>x"9200", 1267=>x"7300",
---- 1268=>x"5800", 1269=>x"6600", 1270=>x"5e00", 1271=>x"3100", 1272=>x"3e00", 1273=>x"3f00", 1274=>x"6700",
---- 1275=>x"7e00", 1276=>x"5000", 1277=>x"2b00", 1278=>x"2700", 1279=>x"2300", 1280=>x"2800", 1281=>x"2800",
---- 1282=>x"4200", 1283=>x"7400", 1284=>x"5800", 1285=>x"2b00", 1286=>x"2300", 1287=>x"2200", 1288=>x"2800",
---- 1289=>x"5400", 1290=>x"8800", 1291=>x"4c00", 1292=>x"2700", 1293=>x"2800", 1294=>x"d600", 1295=>x"2b00",
---- 1296=>x"4300", 1297=>x"7200", 1298=>x"a700", 1299=>x"3d00", 1300=>x"2500", 1301=>x"2c00", 1302=>x"2e00",
---- 1303=>x"2e00", 1304=>x"5200", 1305=>x"7e00", 1306=>x"5500", 1307=>x"2b00", 1308=>x"3200", 1309=>x"3800",
---- 1310=>x"3400", 1311=>x"2d00", 1312=>x"6700", 1313=>x"6c00", 1314=>x"3600", 1315=>x"1d00", 1316=>x"3f00",
---- 1317=>x"4f00", 1318=>x"5900", 1319=>x"5f00", 1320=>x"5d00", 1321=>x"3d00", 1322=>x"4600", 1323=>x"3600",
---- 1324=>x"5500", 1325=>x"6700", 1326=>x"6e00", 1327=>x"8200", 1328=>x"2e00", 1329=>x"3b00", 1330=>x"5e00",
---- 1331=>x"6b00", 1332=>x"6d00", 1333=>x"6f00", 1334=>x"8700", 1335=>x"aa00", 1336=>x"2500", 1337=>x"3c00",
---- 1338=>x"7e00", 1339=>x"8400", 1340=>x"8400", 1341=>x"9c00", 1342=>x"a700", 1343=>x"bc00", 1344=>x"2e00",
---- 1345=>x"7900", 1346=>x"a200", 1347=>x"8e00", 1348=>x"a200", 1349=>x"a800", 1350=>x"b500", 1351=>x"ae00",
---- 1352=>x"5600", 1353=>x"9200", 1354=>x"9d00", 1355=>x"9600", 1356=>x"ab00", 1357=>x"b800", 1358=>x"c500",
---- 1359=>x"8400", 1360=>x"9500", 1361=>x"7400", 1362=>x"8e00", 1363=>x"6100", 1364=>x"ac00", 1365=>x"c600",
---- 1366=>x"a200", 1367=>x"5b00", 1368=>x"6100", 1369=>x"7c00", 1370=>x"9700", 1371=>x"a000", 1372=>x"bf00",
---- 1373=>x"b800", 1374=>x"6400", 1375=>x"5e00", 1376=>x"8400", 1377=>x"8f00", 1378=>x"b400", 1379=>x"b900",
---- 1380=>x"c400", 1381=>x"7300", 1382=>x"5f00", 1383=>x"6200", 1384=>x"c200", 1385=>x"c100", 1386=>x"cb00",
---- 1387=>x"c500", 1388=>x"8100", 1389=>x"5a00", 1390=>x"6100", 1391=>x"5b00", 1392=>x"2e00", 1393=>x"cf00",
---- 1394=>x"cc00", 1395=>x"9200", 1396=>x"5900", 1397=>x"6a00", 1398=>x"5a00", 1399=>x"7000", 1400=>x"ce00",
---- 1401=>x"d100", 1402=>x"ac00", 1403=>x"5900", 1404=>x"6900", 1405=>x"6200", 1406=>x"6200", 1407=>x"ae00",
---- 1408=>x"d600", 1409=>x"cc00", 1410=>x"8000", 1411=>x"5a00", 1412=>x"5f00", 1413=>x"5e00", 1414=>x"9b00",
---- 1415=>x"b800", 1416=>x"d600", 1417=>x"a200", 1418=>x"6300", 1419=>x"6600", 1420=>x"5e00", 1421=>x"8d00",
---- 1422=>x"c500", 1423=>x"6700", 1424=>x"bb00", 1425=>x"6d00", 1426=>x"6300", 1427=>x"6f00", 1428=>x"8f00",
---- 1429=>x"c400", 1430=>x"8d00", 1431=>x"2e00", 1432=>x"7600", 1433=>x"6000", 1434=>x"7800", 1435=>x"9800",
---- 1436=>x"b300", 1437=>x"9d00", 1438=>x"3c00", 1439=>x"2e00", 1440=>x"5900", 1441=>x"8100", 1442=>x"9b00",
---- 1443=>x"bf00", 1444=>x"a000", 1445=>x"4400", 1446=>x"2d00", 1447=>x"3600", 1448=>x"7900", 1449=>x"9e00",
---- 1450=>x"b900", 1451=>x"ba00", 1452=>x"6100", 1453=>x"d200", 1454=>x"3a00", 1455=>x"3400", 1456=>x"a000",
---- 1457=>x"b000", 1458=>x"cf00", 1459=>x"6a00", 1460=>x"3000", 1461=>x"3600", 1462=>x"3400", 1463=>x"3600",
---- 1464=>x"a300", 1465=>x"c500", 1466=>x"8900", 1467=>x"2c00", 1468=>x"3100", 1469=>x"3300", 1470=>x"3100",
---- 1471=>x"3200", 1472=>x"c800", 1473=>x"a100", 1474=>x"3200", 1475=>x"3200", 1476=>x"3300", 1477=>x"3400",
---- 1478=>x"3500", 1479=>x"3300", 1480=>x"be00", 1481=>x"5100", 1482=>x"2c00", 1483=>x"2d00", 1484=>x"3000",
---- 1485=>x"3400", 1486=>x"3000", 1487=>x"3000", 1488=>x"5d00", 1489=>x"2e00", 1490=>x"3200", 1491=>x"3200",
---- 1492=>x"3300", 1493=>x"3800", 1494=>x"3500", 1495=>x"3200", 1496=>x"2600", 1497=>x"3b00", 1498=>x"3000",
---- 1499=>x"3000", 1500=>x"3400", 1501=>x"3200", 1502=>x"3300", 1503=>x"3300", 1504=>x"3900", 1505=>x"4500",
---- 1506=>x"2c00", 1507=>x"3200", 1508=>x"3200", 1509=>x"3400", 1510=>x"3300", 1511=>x"3300", 1512=>x"5200",
---- 1513=>x"3900", 1514=>x"3200", 1515=>x"3500", 1516=>x"3b00", 1517=>x"3500", 1518=>x"3100", 1519=>x"3500",
---- 1520=>x"3f00", 1521=>x"3500", 1522=>x"3100", 1523=>x"3200", 1524=>x"c600", 1525=>x"3500", 1526=>x"3000",
---- 1527=>x"3000", 1528=>x"3400", 1529=>x"3800", 1530=>x"3300", 1531=>x"3200", 1532=>x"3500", 1533=>x"cb00",
---- 1534=>x"3400", 1535=>x"3200", 1536=>x"2e00", 1537=>x"2e00", 1538=>x"2f00", 1539=>x"3400", 1540=>x"3100",
---- 1541=>x"3400", 1542=>x"3600", 1543=>x"3300", 1544=>x"3600", 1545=>x"2e00", 1546=>x"2f00", 1547=>x"3200",
---- 1548=>x"3400", 1549=>x"3400", 1550=>x"3700", 1551=>x"3300", 1552=>x"6e00", 1553=>x"4100", 1554=>x"2d00",
---- 1555=>x"2c00", 1556=>x"2d00", 1557=>x"3000", 1558=>x"3200", 1559=>x"3000", 1560=>x"ae00", 1561=>x"9000",
---- 1562=>x"4400", 1563=>x"2300", 1564=>x"2b00", 1565=>x"2c00", 1566=>x"3000", 1567=>x"3100", 1568=>x"ae00",
---- 1569=>x"ae00", 1570=>x"9100", 1571=>x"4300", 1572=>x"2b00", 1573=>x"3300", 1574=>x"3000", 1575=>x"3400",
---- 1576=>x"8b00", 1577=>x"8800", 1578=>x"9b00", 1579=>x"9600", 1580=>x"3800", 1581=>x"2b00", 1582=>x"3000",
---- 1583=>x"3500", 1584=>x"9700", 1585=>x"7a00", 1586=>x"5b00", 1587=>x"9b00", 1588=>x"8700", 1589=>x"2e00",
---- 1590=>x"2e00", 1591=>x"3500", 1592=>x"b300", 1593=>x"7e00", 1594=>x"5300", 1595=>x"4e00", 1596=>x"a800",
---- 1597=>x"5f00", 1598=>x"2200", 1599=>x"3300", 1600=>x"a700", 1601=>x"5f00", 1602=>x"5100", 1603=>x"4600",
---- 1604=>x"5900", 1605=>x"8400", 1606=>x"3e00", 1607=>x"3200", 1608=>x"8600", 1609=>x"9700", 1610=>x"5600",
---- 1611=>x"3000", 1612=>x"5800", 1613=>x"8500", 1614=>x"7f00", 1615=>x"2e00", 1616=>x"5d00", 1617=>x"8700",
---- 1618=>x"8e00", 1619=>x"3500", 1620=>x"3900", 1621=>x"6400", 1622=>x"9400", 1623=>x"4f00", 1624=>x"5100",
---- 1625=>x"3c00", 1626=>x"7700", 1627=>x"7800", 1628=>x"2400", 1629=>x"3b00", 1630=>x"8100", 1631=>x"8900",
---- 1632=>x"6c00", 1633=>x"1d00", 1634=>x"3e00", 1635=>x"ab00", 1636=>x"6200", 1637=>x"2800", 1638=>x"5300",
---- 1639=>x"9d00", 1640=>x"9600", 1641=>x"3600", 1642=>x"2000", 1643=>x"8500", 1644=>x"b600", 1645=>x"4700",
---- 1646=>x"4800", 1647=>x"8100", 1648=>x"8400", 1649=>x"7000", 1650=>x"3500", 1651=>x"5300", 1652=>x"b600",
---- 1653=>x"9400", 1654=>x"5900", 1655=>x"5600", 1656=>x"6d00", 1657=>x"8d00", 1658=>x"6e00", 1659=>x"6400",
---- 1660=>x"7800", 1661=>x"9600", 1662=>x"6100", 1663=>x"2800", 1664=>x"7a00", 1665=>x"9300", 1666=>x"6600",
---- 1667=>x"6a00", 1668=>x"5200", 1669=>x"6d00", 1670=>x"a700", 1671=>x"2400", 1672=>x"8500", 1673=>x"a200",
---- 1674=>x"8e00", 1675=>x"7d00", 1676=>x"4200", 1677=>x"3500", 1678=>x"b400", 1679=>x"6200", 1680=>x"7f00",
---- 1681=>x"a900", 1682=>x"a500", 1683=>x"7700", 1684=>x"2f00", 1685=>x"1c00", 1686=>x"6000", 1687=>x"8100",
---- 1688=>x"7c00", 1689=>x"9f00", 1690=>x"a700", 1691=>x"7700", 1692=>x"4000", 1693=>x"2000", 1694=>x"2f00",
---- 1695=>x"7600", 1696=>x"8a00", 1697=>x"9400", 1698=>x"8e00", 1699=>x"4500", 1700=>x"4700", 1701=>x"2b00",
---- 1702=>x"3300", 1703=>x"8500", 1704=>x"8d00", 1705=>x"9400", 1706=>x"9300", 1707=>x"4300", 1708=>x"2500",
---- 1709=>x"4d00", 1710=>x"3400", 1711=>x"7500", 1712=>x"9000", 1713=>x"8900", 1714=>x"a600", 1715=>x"6400",
---- 1716=>x"2200", 1717=>x"4100", 1718=>x"2c00", 1719=>x"6c00", 1720=>x"7300", 1721=>x"8b00", 1722=>x"9b00",
---- 1723=>x"6f00", 1724=>x"3d00", 1725=>x"2400", 1726=>x"2500", 1727=>x"6300", 1728=>x"7100", 1729=>x"9800",
---- 1730=>x"8c00", 1731=>x"8000", 1732=>x"7900", 1733=>x"3d00", 1734=>x"2900", 1735=>x"6f00", 1736=>x"8a00",
---- 1737=>x"9d00", 1738=>x"6900", 1739=>x"5300", 1740=>x"9b00", 1741=>x"6a00", 1742=>x"6400", 1743=>x"a200",
---- 1744=>x"9200", 1745=>x"a400", 1746=>x"8f00", 1747=>x"5300", 1748=>x"7d00", 1749=>x"5100", 1750=>x"7500",
---- 1751=>x"af00", 1752=>x"9200", 1753=>x"7a00", 1754=>x"8600", 1755=>x"8a00", 1756=>x"8700", 1757=>x"8a00",
---- 1758=>x"b000", 1759=>x"a000", 1760=>x"8c00", 1761=>x"4b00", 1762=>x"5700", 1763=>x"8a00", 1764=>x"8d00",
---- 1765=>x"a300", 1766=>x"b500", 1767=>x"9300", 1768=>x"8400", 1769=>x"6e00", 1770=>x"5a00", 1771=>x"5a00",
---- 1772=>x"6a00", 1773=>x"8a00", 1774=>x"7c00", 1775=>x"9e00", 1776=>x"8300", 1777=>x"6900", 1778=>x"6100",
---- 1779=>x"2c00", 1780=>x"2100", 1781=>x"4400", 1782=>x"5500", 1783=>x"4200", 1784=>x"6c00", 1785=>x"8000",
---- 1786=>x"6700", 1787=>x"4e00", 1788=>x"1d00", 1789=>x"3000", 1790=>x"5c00", 1791=>x"2300", 1792=>x"6500",
---- 1793=>x"7b00", 1794=>x"8400", 1795=>x"7c00", 1796=>x"3300", 1797=>x"2b00", 1798=>x"6300", 1799=>x"3100",
---- 1800=>x"6900", 1801=>x"6c00", 1802=>x"8700", 1803=>x"9500", 1804=>x"6500", 1805=>x"2500", 1806=>x"6200",
---- 1807=>x"3e00", 1808=>x"5900", 1809=>x"4300", 1810=>x"5e00", 1811=>x"7f00", 1812=>x"8f00", 1813=>x"5100",
---- 1814=>x"5300", 1815=>x"4300", 1816=>x"6600", 1817=>x"4c00", 1818=>x"3a00", 1819=>x"6900", 1820=>x"8000",
---- 1821=>x"8000", 1822=>x"6800", 1823=>x"4e00", 1824=>x"5200", 1825=>x"3f00", 1826=>x"3500", 1827=>x"5a00",
---- 1828=>x"7900", 1829=>x"9100", 1830=>x"8800", 1831=>x"8500", 1832=>x"6d00", 1833=>x"3800", 1834=>x"2f00",
---- 1835=>x"3f00", 1836=>x"ab00", 1837=>x"8300", 1838=>x"a900", 1839=>x"4f00", 1840=>x"9400", 1841=>x"3d00",
---- 1842=>x"3300", 1843=>x"5700", 1844=>x"5400", 1845=>x"4d00", 1846=>x"8100", 1847=>x"8c00", 1848=>x"6200",
---- 1849=>x"4600", 1850=>x"2b00", 1851=>x"5c00", 1852=>x"7c00", 1853=>x"5800", 1854=>x"6200", 1855=>x"7200",
---- 1856=>x"3500", 1857=>x"3300", 1858=>x"d100", 1859=>x"5f00", 1860=>x"6100", 1861=>x"5600", 1862=>x"7a00",
---- 1863=>x"5600", 1864=>x"4900", 1865=>x"4300", 1866=>x"4800", 1867=>x"8f00", 1868=>x"4d00", 1869=>x"3600",
---- 1870=>x"a300", 1871=>x"3e00", 1872=>x"6a00", 1873=>x"7700", 1874=>x"b500", 1875=>x"5300", 1876=>x"3300",
---- 1877=>x"2d00", 1878=>x"2b00", 1879=>x"3400", 1880=>x"5e00", 1881=>x"7300", 1882=>x"5c00", 1883=>x"2f00",
---- 1884=>x"2600", 1885=>x"2e00", 1886=>x"2d00", 1887=>x"3300", 1888=>x"5800", 1889=>x"4700", 1890=>x"6300",
---- 1891=>x"5600", 1892=>x"2e00", 1893=>x"2600", 1894=>x"2e00", 1895=>x"3600", 1896=>x"5b00", 1897=>x"6e00",
---- 1898=>x"8800", 1899=>x"5c00", 1900=>x"2d00", 1901=>x"2600", 1902=>x"3300", 1903=>x"3500", 1904=>x"6800",
---- 1905=>x"6700", 1906=>x"6600", 1907=>x"7c00", 1908=>x"3900", 1909=>x"2600", 1910=>x"3400", 1911=>x"3100",
---- 1912=>x"6200", 1913=>x"5700", 1914=>x"7000", 1915=>x"8300", 1916=>x"3f00", 1917=>x"2d00", 1918=>x"3200",
---- 1919=>x"2c00", 1920=>x"7a00", 1921=>x"6300", 1922=>x"6100", 1923=>x"4500", 1924=>x"2f00", 1925=>x"3100",
---- 1926=>x"2e00", 1927=>x"d500", 1928=>x"7c00", 1929=>x"9400", 1930=>x"5e00", 1931=>x"2600", 1932=>x"3000",
---- 1933=>x"2f00", 1934=>x"2e00", 1935=>x"2e00", 1936=>x"4b00", 1937=>x"6300", 1938=>x"6c00", 1939=>x"3a00",
---- 1940=>x"2f00", 1941=>x"2e00", 1942=>x"2d00", 1943=>x"2d00", 1944=>x"4800", 1945=>x"2800", 1946=>x"5000",
---- 1947=>x"4d00", 1948=>x"2a00", 1949=>x"2c00", 1950=>x"2b00", 1951=>x"d400", 1952=>x"4a00", 1953=>x"3700",
---- 1954=>x"4500", 1955=>x"4a00", 1956=>x"2d00", 1957=>x"2500", 1958=>x"2900", 1959=>x"3000", 1960=>x"7700",
---- 1961=>x"3800", 1962=>x"3600", 1963=>x"c400", 1964=>x"3700", 1965=>x"2300", 1966=>x"2b00", 1967=>x"3100",
---- 1968=>x"6400", 1969=>x"5f00", 1970=>x"3300", 1971=>x"3500", 1972=>x"3400", 1973=>x"2500", 1974=>x"2c00",
---- 1975=>x"2c00", 1976=>x"5f00", 1977=>x"7900", 1978=>x"5a00", 1979=>x"3300", 1980=>x"3100", 1981=>x"2d00",
---- 1982=>x"3000", 1983=>x"2e00", 1984=>x"4500", 1985=>x"6200", 1986=>x"6800", 1987=>x"3e00", 1988=>x"2c00",
---- 1989=>x"2b00", 1990=>x"3400", 1991=>x"3600", 1992=>x"6f00", 1993=>x"5100", 1994=>x"4b00", 1995=>x"4100",
---- 1996=>x"2600", 1997=>x"2700", 1998=>x"2d00", 1999=>x"3100", 2000=>x"7200", 2001=>x"5200", 2002=>x"2a00",
---- 2003=>x"3700", 2004=>x"2f00", 2005=>x"2b00", 2006=>x"2c00", 2007=>x"3000", 2008=>x"6b00", 2009=>x"6900",
---- 2010=>x"4000", 2011=>x"3c00", 2012=>x"3800", 2013=>x"2600", 2014=>x"2900", 2015=>x"2b00", 2016=>x"5d00",
---- 2017=>x"6500", 2018=>x"5f00", 2019=>x"7100", 2020=>x"3b00", 2021=>x"2000", 2022=>x"2100", 2023=>x"2400",
---- 2024=>x"5900", 2025=>x"6c00", 2026=>x"4f00", 2027=>x"7800", 2028=>x"7500", 2029=>x"3600", 2030=>x"2100",
---- 2031=>x"2700", 2032=>x"3b00", 2033=>x"5700", 2034=>x"4a00", 2035=>x"5300", 2036=>x"7f00", 2037=>x"7400",
---- 2038=>x"3c00", 2039=>x"3000", 2040=>x"2f00", 2041=>x"5400", 2042=>x"5a00", 2043=>x"2e00", 2044=>x"5b00",
---- 2045=>x"5b00", 2046=>x"6600", 2047=>x"3d00"),
---- 11 => (0=>x"8600", 1=>x"8600", 2=>x"8500", 3=>x"8300", 4=>x"8500", 5=>x"8800", 6=>x"8400", 7=>x"7b00",
---- 8=>x"8600", 9=>x"8500", 10=>x"8600", 11=>x"8300", 12=>x"8500", 13=>x"8800", 14=>x"8500",
---- 15=>x"8400", 16=>x"8700", 17=>x"8600", 18=>x"8500", 19=>x"7c00", 20=>x"8500", 21=>x"8600",
---- 22=>x"8500", 23=>x"8400", 24=>x"8400", 25=>x"8500", 26=>x"8500", 27=>x"8300", 28=>x"8200",
---- 29=>x"8200", 30=>x"8200", 31=>x"8300", 32=>x"8200", 33=>x"8400", 34=>x"8700", 35=>x"8600",
---- 36=>x"8100", 37=>x"8600", 38=>x"8500", 39=>x"8400", 40=>x"7b00", 41=>x"8600", 42=>x"8600",
---- 43=>x"8100", 44=>x"8200", 45=>x"8500", 46=>x"8400", 47=>x"8300", 48=>x"8500", 49=>x"8400",
---- 50=>x"8200", 51=>x"8300", 52=>x"8500", 53=>x"8300", 54=>x"8300", 55=>x"8400", 56=>x"8300",
---- 57=>x"8200", 58=>x"8200", 59=>x"8500", 60=>x"8500", 61=>x"8400", 62=>x"8700", 63=>x"8200",
---- 64=>x"8700", 65=>x"8600", 66=>x"8500", 67=>x"8400", 68=>x"8400", 69=>x"8500", 70=>x"8600",
---- 71=>x"8400", 72=>x"8600", 73=>x"8700", 74=>x"8500", 75=>x"8300", 76=>x"8300", 77=>x"8300",
---- 78=>x"8500", 79=>x"8400", 80=>x"8400", 81=>x"8200", 82=>x"8100", 83=>x"8500", 84=>x"8200",
---- 85=>x"8200", 86=>x"8400", 87=>x"8200", 88=>x"8300", 89=>x"8200", 90=>x"8200", 91=>x"8200",
---- 92=>x"8100", 93=>x"8000", 94=>x"8500", 95=>x"8200", 96=>x"8400", 97=>x"8100", 98=>x"8200",
---- 99=>x"8100", 100=>x"8200", 101=>x"8000", 102=>x"8300", 103=>x"8300", 104=>x"8300", 105=>x"8300",
---- 106=>x"8100", 107=>x"8000", 108=>x"8100", 109=>x"8300", 110=>x"8400", 111=>x"8500", 112=>x"8300",
---- 113=>x"8200", 114=>x"8000", 115=>x"7d00", 116=>x"8100", 117=>x"8200", 118=>x"8100", 119=>x"8400",
---- 120=>x"8100", 121=>x"8200", 122=>x"8000", 123=>x"8000", 124=>x"8200", 125=>x"7c00", 126=>x"8100",
---- 127=>x"8400", 128=>x"7f00", 129=>x"8100", 130=>x"8400", 131=>x"8400", 132=>x"8100", 133=>x"7f00",
---- 134=>x"8300", 135=>x"8200", 136=>x"8000", 137=>x"8100", 138=>x"8100", 139=>x"8100", 140=>x"8000",
---- 141=>x"8100", 142=>x"8000", 143=>x"8100", 144=>x"8100", 145=>x"8200", 146=>x"8300", 147=>x"8200",
---- 148=>x"8100", 149=>x"8100", 150=>x"7f00", 151=>x"8100", 152=>x"8100", 153=>x"8100", 154=>x"8600",
---- 155=>x"8400", 156=>x"8300", 157=>x"8000", 158=>x"8000", 159=>x"7f00", 160=>x"8000", 161=>x"8000",
---- 162=>x"8200", 163=>x"7f00", 164=>x"8000", 165=>x"8100", 166=>x"7f00", 167=>x"8000", 168=>x"8300",
---- 169=>x"8100", 170=>x"8000", 171=>x"8000", 172=>x"8200", 173=>x"8000", 174=>x"7f00", 175=>x"8100",
---- 176=>x"8000", 177=>x"8100", 178=>x"8100", 179=>x"8200", 180=>x"8000", 181=>x"8100", 182=>x"7e00",
---- 183=>x"7e00", 184=>x"8200", 185=>x"8600", 186=>x"8200", 187=>x"7e00", 188=>x"8000", 189=>x"7f00",
---- 190=>x"8100", 191=>x"7f00", 192=>x"8200", 193=>x"8400", 194=>x"8100", 195=>x"8000", 196=>x"8000",
---- 197=>x"8000", 198=>x"8000", 199=>x"7e00", 200=>x"8700", 201=>x"7f00", 202=>x"8000", 203=>x"8100",
---- 204=>x"7f00", 205=>x"7f00", 206=>x"7c00", 207=>x"7a00", 208=>x"8200", 209=>x"8000", 210=>x"7f00",
---- 211=>x"7e00", 212=>x"7e00", 213=>x"7d00", 214=>x"8100", 215=>x"8800", 216=>x"7d00", 217=>x"7c00",
---- 218=>x"7d00", 219=>x"7f00", 220=>x"8000", 221=>x"8000", 222=>x"8a00", 223=>x"9500", 224=>x"8800",
---- 225=>x"8900", 226=>x"8800", 227=>x"8100", 228=>x"7f00", 229=>x"8600", 230=>x"9500", 231=>x"9100",
---- 232=>x"9400", 233=>x"8900", 234=>x"7d00", 235=>x"7500", 236=>x"7e00", 237=>x"8600", 238=>x"8b00",
---- 239=>x"8a00", 240=>x"8100", 241=>x"7e00", 242=>x"7900", 243=>x"7a00", 244=>x"7b00", 245=>x"7d00",
---- 246=>x"8400", 247=>x"8700", 248=>x"7f00", 249=>x"7d00", 250=>x"7900", 251=>x"7a00", 252=>x"7900",
---- 253=>x"7e00", 254=>x"8a00", 255=>x"8700", 256=>x"7c00", 257=>x"7a00", 258=>x"7d00", 259=>x"7c00",
---- 260=>x"7e00", 261=>x"8200", 262=>x"8800", 263=>x"8300", 264=>x"7a00", 265=>x"7900", 266=>x"7a00",
---- 267=>x"7600", 268=>x"7900", 269=>x"8500", 270=>x"8500", 271=>x"8400", 272=>x"8000", 273=>x"7a00",
---- 274=>x"7600", 275=>x"7700", 276=>x"7b00", 277=>x"7e00", 278=>x"8100", 279=>x"8500", 280=>x"7b00",
---- 281=>x"7c00", 282=>x"7600", 283=>x"7b00", 284=>x"8000", 285=>x"8400", 286=>x"8800", 287=>x"8600",
---- 288=>x"7900", 289=>x"7c00", 290=>x"8000", 291=>x"7e00", 292=>x"7900", 293=>x"8700", 294=>x"8100",
---- 295=>x"8200", 296=>x"7c00", 297=>x"8300", 298=>x"7d00", 299=>x"7700", 300=>x"8500", 301=>x"8100",
---- 302=>x"7500", 303=>x"8100", 304=>x"7b00", 305=>x"7a00", 306=>x"7a00", 307=>x"8000", 308=>x"7e00",
---- 309=>x"7a00", 310=>x"7f00", 311=>x"8300", 312=>x"7100", 313=>x"7b00", 314=>x"7e00", 315=>x"8100",
---- 316=>x"7900", 317=>x"7c00", 318=>x"8300", 319=>x"8300", 320=>x"7700", 321=>x"7e00", 322=>x"7c00",
---- 323=>x"7d00", 324=>x"7900", 325=>x"7f00", 326=>x"8000", 327=>x"8100", 328=>x"7c00", 329=>x"7600",
---- 330=>x"7d00", 331=>x"7800", 332=>x"7600", 333=>x"7d00", 334=>x"7800", 335=>x"7c00", 336=>x"7600",
---- 337=>x"7900", 338=>x"7a00", 339=>x"7500", 340=>x"7800", 341=>x"7800", 342=>x"7800", 343=>x"7a00",
---- 344=>x"7a00", 345=>x"7700", 346=>x"7800", 347=>x"7800", 348=>x"7400", 349=>x"7700", 350=>x"8000",
---- 351=>x"7d00", 352=>x"7800", 353=>x"7400", 354=>x"7300", 355=>x"7100", 356=>x"7400", 357=>x"7d00",
---- 358=>x"7d00", 359=>x"8400", 360=>x"6f00", 361=>x"7100", 362=>x"7400", 363=>x"7a00", 364=>x"7700",
---- 365=>x"7f00", 366=>x"8300", 367=>x"7900", 368=>x"6b00", 369=>x"6e00", 370=>x"7900", 371=>x"8000",
---- 372=>x"8000", 373=>x"8000", 374=>x"7d00", 375=>x"7f00", 376=>x"7100", 377=>x"7600", 378=>x"7800",
---- 379=>x"8000", 380=>x"8400", 381=>x"7e00", 382=>x"8100", 383=>x"8200", 384=>x"7700", 385=>x"7800",
---- 386=>x"7900", 387=>x"7c00", 388=>x"8100", 389=>x"8100", 390=>x"7f00", 391=>x"8500", 392=>x"7500",
---- 393=>x"7c00", 394=>x"7e00", 395=>x"8400", 396=>x"7f00", 397=>x"7a00", 398=>x"8100", 399=>x"8000",
---- 400=>x"7700", 401=>x"7c00", 402=>x"8200", 403=>x"8200", 404=>x"8000", 405=>x"7f00", 406=>x"7d00",
---- 407=>x"8600", 408=>x"8000", 409=>x"8900", 410=>x"8400", 411=>x"8100", 412=>x"7f00", 413=>x"8800",
---- 414=>x"8900", 415=>x"8b00", 416=>x"8400", 417=>x"8200", 418=>x"7f00", 419=>x"8600", 420=>x"8900",
---- 421=>x"8c00", 422=>x"9100", 423=>x"9000", 424=>x"7b00", 425=>x"8200", 426=>x"8900", 427=>x"8500",
---- 428=>x"8700", 429=>x"9000", 430=>x"9000", 431=>x"8c00", 432=>x"7d00", 433=>x"8300", 434=>x"8700",
---- 435=>x"8300", 436=>x"8c00", 437=>x"9400", 438=>x"8d00", 439=>x"8200", 440=>x"7e00", 441=>x"7e00",
---- 442=>x"8700", 443=>x"8d00", 444=>x"9200", 445=>x"8900", 446=>x"7f00", 447=>x"8200", 448=>x"8400",
---- 449=>x"8600", 450=>x"8f00", 451=>x"8b00", 452=>x"8500", 453=>x"8200", 454=>x"8800", 455=>x"8200",
---- 456=>x"8600", 457=>x"8700", 458=>x"8300", 459=>x"8600", 460=>x"8b00", 461=>x"8d00", 462=>x"8800",
---- 463=>x"8800", 464=>x"8b00", 465=>x"8a00", 466=>x"8400", 467=>x"8500", 468=>x"8f00", 469=>x"8d00",
---- 470=>x"8000", 471=>x"7f00", 472=>x"8a00", 473=>x"8d00", 474=>x"8300", 475=>x"8500", 476=>x"8500",
---- 477=>x"7d00", 478=>x"8100", 479=>x"8700", 480=>x"8000", 481=>x"7d00", 482=>x"8700", 483=>x"7800",
---- 484=>x"7300", 485=>x"8300", 486=>x"8900", 487=>x"8800", 488=>x"7c00", 489=>x"7e00", 490=>x"6c00",
---- 491=>x"7100", 492=>x"8700", 493=>x"8d00", 494=>x"8800", 495=>x"7b00", 496=>x"7700", 497=>x"7100",
---- 498=>x"8700", 499=>x"8700", 500=>x"8b00", 501=>x"8300", 502=>x"7b00", 503=>x"7f00", 504=>x"7400",
---- 505=>x"8300", 506=>x"8d00", 507=>x"8600", 508=>x"7900", 509=>x"7700", 510=>x"8200", 511=>x"8100",
---- 512=>x"8000", 513=>x"8600", 514=>x"8800", 515=>x"7a00", 516=>x"7900", 517=>x"8600", 518=>x"8300",
---- 519=>x"7600", 520=>x"8400", 521=>x"8400", 522=>x"8600", 523=>x"8b00", 524=>x"8600", 525=>x"8400",
---- 526=>x"7700", 527=>x"6700", 528=>x"8600", 529=>x"8500", 530=>x"8300", 531=>x"8100", 532=>x"8000",
---- 533=>x"7800", 534=>x"5f00", 535=>x"6a00", 536=>x"8300", 537=>x"7700", 538=>x"7200", 539=>x"7d00",
---- 540=>x"7900", 541=>x"6100", 542=>x"6d00", 543=>x"8d00", 544=>x"7400", 545=>x"7600", 546=>x"7800",
---- 547=>x"7400", 548=>x"6600", 549=>x"7400", 550=>x"9300", 551=>x"a000", 552=>x"7800", 553=>x"7b00",
---- 554=>x"7500", 555=>x"6900", 556=>x"7600", 557=>x"8c00", 558=>x"9700", 559=>x"9d00", 560=>x"7600",
---- 561=>x"7200", 562=>x"7100", 563=>x"7f00", 564=>x"9500", 565=>x"9000", 566=>x"9400", 567=>x"9a00",
---- 568=>x"7a00", 569=>x"6f00", 570=>x"7e00", 571=>x"9c00", 572=>x"9300", 573=>x"9700", 574=>x"9300",
---- 575=>x"9200", 576=>x"6b00", 577=>x"7900", 578=>x"9400", 579=>x"9600", 580=>x"9400", 581=>x"9c00",
---- 582=>x"9600", 583=>x"8600", 584=>x"7800", 585=>x"9500", 586=>x"9000", 587=>x"9400", 588=>x"9900",
---- 589=>x"9700", 590=>x"8e00", 591=>x"8700", 592=>x"9300", 593=>x"9700", 594=>x"9300", 595=>x"9100",
---- 596=>x"9100", 597=>x"8d00", 598=>x"8e00", 599=>x"9800", 600=>x"9200", 601=>x"9400", 602=>x"9700",
---- 603=>x"8c00", 604=>x"8200", 605=>x"8b00", 606=>x"9f00", 607=>x"8e00", 608=>x"9000", 609=>x"9700",
---- 610=>x"8e00", 611=>x"8b00", 612=>x"8900", 613=>x"9a00", 614=>x"8b00", 615=>x"7200", 616=>x"9300",
---- 617=>x"8f00", 618=>x"8b00", 619=>x"8a00", 620=>x"9c00", 621=>x"8400", 622=>x"6e00", 623=>x"8100",
---- 624=>x"8d00", 625=>x"8900", 626=>x"9200", 627=>x"9900", 628=>x"7800", 629=>x"7100", 630=>x"8200",
---- 631=>x"9300", 632=>x"8400", 633=>x"8d00", 634=>x"9b00", 635=>x"7e00", 636=>x"6b00", 637=>x"7e00",
---- 638=>x"8f00", 639=>x"9400", 640=>x"8a00", 641=>x"9400", 642=>x"7a00", 643=>x"7200", 644=>x"7e00",
---- 645=>x"8c00", 646=>x"8a00", 647=>x"9200", 648=>x"8c00", 649=>x"7500", 650=>x"7100", 651=>x"7900",
---- 652=>x"8b00", 653=>x"9300", 654=>x"8c00", 655=>x"8e00", 656=>x"6d00", 657=>x"7c00", 658=>x"7f00",
---- 659=>x"8a00", 660=>x"8e00", 661=>x"8f00", 662=>x"9600", 663=>x"8d00", 664=>x"7300", 665=>x"8600",
---- 666=>x"8800", 667=>x"9700", 668=>x"8f00", 669=>x"8e00", 670=>x"9600", 671=>x"8d00", 672=>x"7800",
---- 673=>x"8800", 674=>x"8e00", 675=>x"8a00", 676=>x"9000", 677=>x"9700", 678=>x"8b00", 679=>x"8c00",
---- 680=>x"8600", 681=>x"9400", 682=>x"8b00", 683=>x"8700", 684=>x"8e00", 685=>x"8c00", 686=>x"8800",
---- 687=>x"8d00", 688=>x"6b00", 689=>x"9000", 690=>x"8a00", 691=>x"8c00", 692=>x"8b00", 693=>x"8f00",
---- 694=>x"8c00", 695=>x"7300", 696=>x"7400", 697=>x"8f00", 698=>x"8b00", 699=>x"8400", 700=>x"8e00",
---- 701=>x"8700", 702=>x"7800", 703=>x"8000", 704=>x"8800", 705=>x"8500", 706=>x"8900", 707=>x"8800",
---- 708=>x"8000", 709=>x"7500", 710=>x"7800", 711=>x"8500", 712=>x"8900", 713=>x"8800", 714=>x"8900",
---- 715=>x"7e00", 716=>x"7000", 717=>x"8100", 718=>x"8300", 719=>x"8100", 720=>x"8900", 721=>x"8f00",
---- 722=>x"7b00", 723=>x"7800", 724=>x"8000", 725=>x"8200", 726=>x"8100", 727=>x"8800", 728=>x"8900",
---- 729=>x"7d00", 730=>x"7500", 731=>x"8500", 732=>x"8300", 733=>x"8600", 734=>x"8300", 735=>x"8400",
---- 736=>x"7c00", 737=>x"6f00", 738=>x"7b00", 739=>x"8200", 740=>x"8600", 741=>x"8800", 742=>x"8800",
---- 743=>x"8300", 744=>x"7400", 745=>x"7f00", 746=>x"8000", 747=>x"8300", 748=>x"8700", 749=>x"8600",
---- 750=>x"8400", 751=>x"8300", 752=>x"8200", 753=>x"7c00", 754=>x"8200", 755=>x"8500", 756=>x"8300",
---- 757=>x"8500", 758=>x"8000", 759=>x"7700", 760=>x"7f00", 761=>x"7d00", 762=>x"8000", 763=>x"8700",
---- 764=>x"8400", 765=>x"7d00", 766=>x"7800", 767=>x"8200", 768=>x"8100", 769=>x"8000", 770=>x"8000",
---- 771=>x"8500", 772=>x"8100", 773=>x"7900", 774=>x"7800", 775=>x"8a00", 776=>x"8400", 777=>x"8300",
---- 778=>x"7900", 779=>x"7e00", 780=>x"7d00", 781=>x"7300", 782=>x"8700", 783=>x"8d00", 784=>x"7d00",
---- 785=>x"8100", 786=>x"7f00", 787=>x"7800", 788=>x"7300", 789=>x"7b00", 790=>x"7f00", 791=>x"6e00",
---- 792=>x"7500", 793=>x"7d00", 794=>x"8000", 795=>x"7500", 796=>x"7e00", 797=>x"8f00", 798=>x"8900",
---- 799=>x"8400", 800=>x"7400", 801=>x"8300", 802=>x"7800", 803=>x"7b00", 804=>x"8800", 805=>x"8d00",
---- 806=>x"8f00", 807=>x"8c00", 808=>x"7900", 809=>x"7d00", 810=>x"8600", 811=>x"7500", 812=>x"8700",
---- 813=>x"8400", 814=>x"8100", 815=>x"7700", 816=>x"7800", 817=>x"7900", 818=>x"8600", 819=>x"8900",
---- 820=>x"7800", 821=>x"6c00", 822=>x"6a00", 823=>x"6f00", 824=>x"7700", 825=>x"7600", 826=>x"8600",
---- 827=>x"8100", 828=>x"8000", 829=>x"8000", 830=>x"7f00", 831=>x"7000", 832=>x"8000", 833=>x"7f00",
---- 834=>x"7000", 835=>x"6b00", 836=>x"7d00", 837=>x"7b00", 838=>x"6e00", 839=>x"5300", 840=>x"8200",
---- 841=>x"8400", 842=>x"8300", 843=>x"8300", 844=>x"7100", 845=>x"6600", 846=>x"4b00", 847=>x"4100",
---- 848=>x"8200", 849=>x"7200", 850=>x"6300", 851=>x"8a00", 852=>x"8300", 853=>x"6c00", 854=>x"4800",
---- 855=>x"4200", 856=>x"8200", 857=>x"6f00", 858=>x"6000", 859=>x"7a00", 860=>x"6f00", 861=>x"6100",
---- 862=>x"4800", 863=>x"4600", 864=>x"7700", 865=>x"6400", 866=>x"5900", 867=>x"6500", 868=>x"4a00",
---- 869=>x"3f00", 870=>x"5500", 871=>x"5000", 872=>x"7d00", 873=>x"5a00", 874=>x"3300", 875=>x"3c00",
---- 876=>x"3000", 877=>x"3700", 878=>x"5a00", 879=>x"3e00", 880=>x"7f00", 881=>x"5d00", 882=>x"2a00",
---- 883=>x"2a00", 884=>x"3300", 885=>x"4900", 886=>x"4900", 887=>x"3100", 888=>x"6f00", 889=>x"6100",
---- 890=>x"3200", 891=>x"2800", 892=>x"4000", 893=>x"5f00", 894=>x"3800", 895=>x"2800", 896=>x"4700",
---- 897=>x"4e00", 898=>x"3c00", 899=>x"2d00", 900=>x"5000", 901=>x"5d00", 902=>x"2e00", 903=>x"2900",
---- 904=>x"3f00", 905=>x"4e00", 906=>x"3800", 907=>x"2800", 908=>x"5f00", 909=>x"5200", 910=>x"2a00",
---- 911=>x"2a00", 912=>x"3000", 913=>x"2e00", 914=>x"2700", 915=>x"3000", 916=>x"6100", 917=>x"b500",
---- 918=>x"2500", 919=>x"2b00", 920=>x"3c00", 921=>x"2800", 922=>x"2900", 923=>x"d600", 924=>x"5500",
---- 925=>x"4800", 926=>x"2400", 927=>x"3100", 928=>x"3900", 929=>x"2400", 930=>x"2900", 931=>x"2600",
---- 932=>x"4a00", 933=>x"5800", 934=>x"3c00", 935=>x"4300", 936=>x"2a00", 937=>x"2700", 938=>x"2c00",
---- 939=>x"2700", 940=>x"3300", 941=>x"6200", 942=>x"4700", 943=>x"2e00", 944=>x"2500", 945=>x"3700",
---- 946=>x"3900", 947=>x"2d00", 948=>x"2800", 949=>x"3800", 950=>x"5200", 951=>x"2c00", 952=>x"2b00",
---- 953=>x"4c00", 954=>x"2e00", 955=>x"3400", 956=>x"2900", 957=>x"2600", 958=>x"3600", 959=>x"5100",
---- 960=>x"3a00", 961=>x"3100", 962=>x"2b00", 963=>x"3400", 964=>x"3d00", 965=>x"3700", 966=>x"4d00",
---- 967=>x"6600", 968=>x"3900", 969=>x"2100", 970=>x"3100", 971=>x"2700", 972=>x"3e00", 973=>x"5a00",
---- 974=>x"6800", 975=>x"5100", 976=>x"2400", 977=>x"2800", 978=>x"3300", 979=>x"3500", 980=>x"4600",
---- 981=>x"4500", 982=>x"3900", 983=>x"3a00", 984=>x"1c00", 985=>x"3000", 986=>x"3200", 987=>x"3100",
---- 988=>x"3500", 989=>x"2f00", 990=>x"3200", 991=>x"3b00", 992=>x"1c00", 993=>x"2b00", 994=>x"2800",
---- 995=>x"2e00", 996=>x"4000", 997=>x"4500", 998=>x"3200", 999=>x"4200", 1000=>x"1e00", 1001=>x"2600",
---- 1002=>x"2c00", 1003=>x"4800", 1004=>x"4600", 1005=>x"3d00", 1006=>x"4300", 1007=>x"3d00", 1008=>x"3400",
---- 1009=>x"2400", 1010=>x"3000", 1011=>x"4700", 1012=>x"3d00", 1013=>x"2f00", 1014=>x"3600", 1015=>x"4200",
---- 1016=>x"5000", 1017=>x"2600", 1018=>x"2c00", 1019=>x"4b00", 1020=>x"3900", 1021=>x"2500", 1022=>x"2500",
---- 1023=>x"3700", 1024=>x"5800", 1025=>x"2b00", 1026=>x"2c00", 1027=>x"5400", 1028=>x"3d00", 1029=>x"2700",
---- 1030=>x"2500", 1031=>x"3000", 1032=>x"4c00", 1033=>x"3a00", 1034=>x"2600", 1035=>x"5800", 1036=>x"3b00",
---- 1037=>x"2300", 1038=>x"2500", 1039=>x"2a00", 1040=>x"3100", 1041=>x"4700", 1042=>x"3000", 1043=>x"5a00",
---- 1044=>x"4300", 1045=>x"2400", 1046=>x"2700", 1047=>x"2400", 1048=>x"2e00", 1049=>x"3b00", 1050=>x"4200",
---- 1051=>x"5f00", 1052=>x"5300", 1053=>x"2600", 1054=>x"2f00", 1055=>x"2700", 1056=>x"3000", 1057=>x"2f00",
---- 1058=>x"2a00", 1059=>x"5500", 1060=>x"6500", 1061=>x"2900", 1062=>x"2f00", 1063=>x"2d00", 1064=>x"2600",
---- 1065=>x"3100", 1066=>x"2600", 1067=>x"3f00", 1068=>x"7400", 1069=>x"3800", 1070=>x"3300", 1071=>x"2600",
---- 1072=>x"2d00", 1073=>x"2f00", 1074=>x"2700", 1075=>x"3000", 1076=>x"6f00", 1077=>x"5200", 1078=>x"2e00",
---- 1079=>x"2900", 1080=>x"3500", 1081=>x"3200", 1082=>x"2800", 1083=>x"2b00", 1084=>x"5900", 1085=>x"4f00",
---- 1086=>x"2800", 1087=>x"3400", 1088=>x"3800", 1089=>x"3000", 1090=>x"2c00", 1091=>x"2c00", 1092=>x"3c00",
---- 1093=>x"3500", 1094=>x"2e00", 1095=>x"3b00", 1096=>x"3300", 1097=>x"2700", 1098=>x"2500", 1099=>x"2c00",
---- 1100=>x"3300", 1101=>x"2f00", 1102=>x"3900", 1103=>x"3a00", 1104=>x"2c00", 1105=>x"2700", 1106=>x"2800",
---- 1107=>x"2d00", 1108=>x"3100", 1109=>x"2e00", 1110=>x"3100", 1111=>x"2e00", 1112=>x"2d00", 1113=>x"2c00",
---- 1114=>x"2e00", 1115=>x"2a00", 1116=>x"2d00", 1117=>x"2f00", 1118=>x"3000", 1119=>x"2b00", 1120=>x"3500",
---- 1121=>x"2d00", 1122=>x"3100", 1123=>x"3000", 1124=>x"2d00", 1125=>x"3000", 1126=>x"2e00", 1127=>x"2d00",
---- 1128=>x"2e00", 1129=>x"2c00", 1130=>x"2f00", 1131=>x"3000", 1132=>x"2e00", 1133=>x"2e00", 1134=>x"3400",
---- 1135=>x"3000", 1136=>x"2f00", 1137=>x"2a00", 1138=>x"2c00", 1139=>x"2d00", 1140=>x"2c00", 1141=>x"2a00",
---- 1142=>x"3200", 1143=>x"3200", 1144=>x"2f00", 1145=>x"2e00", 1146=>x"3000", 1147=>x"2d00", 1148=>x"2b00",
---- 1149=>x"2b00", 1150=>x"2f00", 1151=>x"3600", 1152=>x"3400", 1153=>x"2f00", 1154=>x"3400", 1155=>x"3300",
---- 1156=>x"2b00", 1157=>x"2c00", 1158=>x"2d00", 1159=>x"3100", 1160=>x"4c00", 1161=>x"2c00", 1162=>x"2a00",
---- 1163=>x"3500", 1164=>x"2c00", 1165=>x"2c00", 1166=>x"2d00", 1167=>x"2e00", 1168=>x"5b00", 1169=>x"3400",
---- 1170=>x"2e00", 1171=>x"3200", 1172=>x"3000", 1173=>x"2e00", 1174=>x"2f00", 1175=>x"2f00", 1176=>x"4b00",
---- 1177=>x"3500", 1178=>x"2b00", 1179=>x"2e00", 1180=>x"2e00", 1181=>x"2e00", 1182=>x"2d00", 1183=>x"2d00",
---- 1184=>x"5f00", 1185=>x"3e00", 1186=>x"2b00", 1187=>x"2b00", 1188=>x"2d00", 1189=>x"2a00", 1190=>x"2e00",
---- 1191=>x"2d00", 1192=>x"7b00", 1193=>x"3200", 1194=>x"2d00", 1195=>x"2a00", 1196=>x"2800", 1197=>x"2600",
---- 1198=>x"2c00", 1199=>x"2700", 1200=>x"9700", 1201=>x"5100", 1202=>x"2000", 1203=>x"2500", 1204=>x"2700",
---- 1205=>x"2200", 1206=>x"2600", 1207=>x"2100", 1208=>x"ac00", 1209=>x"9200", 1210=>x"4500", 1211=>x"2800",
---- 1212=>x"2700", 1213=>x"2300", 1214=>x"2500", 1215=>x"2300", 1216=>x"7400", 1217=>x"9b00", 1218=>x"9a00",
---- 1219=>x"3b00", 1220=>x"2200", 1221=>x"2700", 1222=>x"2900", 1223=>x"2300", 1224=>x"3600", 1225=>x"7500",
---- 1226=>x"aa00", 1227=>x"5e00", 1228=>x"1c00", 1229=>x"2500", 1230=>x"1e00", 1231=>x"2f00", 1232=>x"2f00",
---- 1233=>x"4d00", 1234=>x"8600", 1235=>x"5400", 1236=>x"1b00", 1237=>x"1e00", 1238=>x"1900", 1239=>x"5d00",
---- 1240=>x"3500", 1241=>x"3300", 1242=>x"6400", 1243=>x"3200", 1244=>x"1c00", 1245=>x"1b00", 1246=>x"2900",
---- 1247=>x"8000", 1248=>x"3b00", 1249=>x"2500", 1250=>x"3700", 1251=>x"2600", 1252=>x"2300", 1253=>x"1a00",
---- 1254=>x"4a00", 1255=>x"9000", 1256=>x"2a00", 1257=>x"2800", 1258=>x"3300", 1259=>x"2200", 1260=>x"2400",
---- 1261=>x"4000", 1262=>x"6f00", 1263=>x"7d00", 1264=>x"2300", 1265=>x"2900", 1266=>x"2900", 1267=>x"1d00",
---- 1268=>x"5000", 1269=>x"8400", 1270=>x"7f00", 1271=>x"6d00", 1272=>x"2400", 1273=>x"2b00", 1274=>x"1c00",
---- 1275=>x"3800", 1276=>x"9f00", 1277=>x"a600", 1278=>x"9800", 1279=>x"8f00", 1280=>x"2900", 1281=>x"2400",
---- 1282=>x"1600", 1283=>x"6300", 1284=>x"ac00", 1285=>x"a500", 1286=>x"ab00", 1287=>x"ac00", 1288=>x"2700",
---- 1289=>x"1f00", 1290=>x"1d00", 1291=>x"8e00", 1292=>x"b400", 1293=>x"b200", 1294=>x"b600", 1295=>x"b500",
---- 1296=>x"2300", 1297=>x"1800", 1298=>x"3d00", 1299=>x"a100", 1300=>x"aa00", 1301=>x"b900", 1302=>x"be00",
---- 1303=>x"c000", 1304=>x"3200", 1305=>x"3400", 1306=>x"6700", 1307=>x"8f00", 1308=>x"9a00", 1309=>x"a900",
---- 1310=>x"af00", 1311=>x"b700", 1312=>x"6300", 1313=>x"7700", 1314=>x"7200", 1315=>x"7400", 1316=>x"8200",
---- 1317=>x"7d00", 1318=>x"9e00", 1319=>x"bf00", 1320=>x"9f00", 1321=>x"9c00", 1322=>x"6800", 1323=>x"6800",
---- 1324=>x"6800", 1325=>x"7f00", 1326=>x"2f00", 1327=>x"af00", 1328=>x"b700", 1329=>x"6e00", 1330=>x"6500",
---- 1331=>x"6b00", 1332=>x"7b00", 1333=>x"b100", 1334=>x"cf00", 1335=>x"4d00", 1336=>x"8800", 1337=>x"5700",
---- 1338=>x"5e00", 1339=>x"7300", 1340=>x"a300", 1341=>x"d100", 1342=>x"7500", 1343=>x"2800", 1344=>x"5d00",
---- 1345=>x"5e00", 1346=>x"5700", 1347=>x"6900", 1348=>x"c300", 1349=>x"8b00", 1350=>x"2600", 1351=>x"2a00",
---- 1352=>x"5d00", 1353=>x"a200", 1354=>x"5900", 1355=>x"9900", 1356=>x"a800", 1357=>x"3000", 1358=>x"2300",
---- 1359=>x"2d00", 1360=>x"5e00", 1361=>x"5700", 1362=>x"7a00", 1363=>x"b300", 1364=>x"4a00", 1365=>x"2300",
---- 1366=>x"2f00", 1367=>x"3100", 1368=>x"5800", 1369=>x"6500", 1370=>x"b400", 1371=>x"5e00", 1372=>x"1f00",
---- 1373=>x"2700", 1374=>x"3100", 1375=>x"4400", 1376=>x"6400", 1377=>x"5f00", 1378=>x"8e00", 1379=>x"2500",
---- 1380=>x"2c00", 1381=>x"2400", 1382=>x"4100", 1383=>x"5c00", 1384=>x"8c00", 1385=>x"ae00", 1386=>x"3500",
---- 1387=>x"2700", 1388=>x"2900", 1389=>x"2500", 1390=>x"4100", 1391=>x"6600", 1392=>x"ba00", 1393=>x"5c00",
---- 1394=>x"1c00", 1395=>x"2700", 1396=>x"2c00", 1397=>x"2900", 1398=>x"3000", 1399=>x"5200", 1400=>x"9a00",
---- 1401=>x"2300", 1402=>x"2f00", 1403=>x"3000", 1404=>x"3500", 1405=>x"d600", 1406=>x"2a00", 1407=>x"4800",
---- 1408=>x"4000", 1409=>x"2600", 1410=>x"2f00", 1411=>x"3200", 1412=>x"2f00", 1413=>x"2c00", 1414=>x"2b00",
---- 1415=>x"3b00", 1416=>x"2200", 1417=>x"3400", 1418=>x"3500", 1419=>x"3300", 1420=>x"3100", 1421=>x"2a00",
---- 1422=>x"2a00", 1423=>x"3c00", 1424=>x"3400", 1425=>x"3400", 1426=>x"3600", 1427=>x"3500", 1428=>x"3000",
---- 1429=>x"2a00", 1430=>x"2a00", 1431=>x"3600", 1432=>x"3300", 1433=>x"3300", 1434=>x"3300", 1435=>x"3500",
---- 1436=>x"3200", 1437=>x"2e00", 1438=>x"2c00", 1439=>x"2b00", 1440=>x"3000", 1441=>x"3200", 1442=>x"3700",
---- 1443=>x"3800", 1444=>x"3600", 1445=>x"2f00", 1446=>x"2c00", 1447=>x"3100", 1448=>x"3500", 1449=>x"3600",
---- 1450=>x"3b00", 1451=>x"3700", 1452=>x"c100", 1453=>x"3500", 1454=>x"3300", 1455=>x"3700", 1456=>x"3600",
---- 1457=>x"3700", 1458=>x"3a00", 1459=>x"3b00", 1460=>x"3b00", 1461=>x"3100", 1462=>x"3200", 1463=>x"3a00",
---- 1464=>x"3300", 1465=>x"3400", 1466=>x"3700", 1467=>x"3900", 1468=>x"3700", 1469=>x"d200", 1470=>x"2b00",
---- 1471=>x"3700", 1472=>x"3100", 1473=>x"3800", 1474=>x"3900", 1475=>x"3900", 1476=>x"3b00", 1477=>x"3100",
---- 1478=>x"3200", 1479=>x"3900", 1480=>x"2e00", 1481=>x"3400", 1482=>x"3900", 1483=>x"3500", 1484=>x"3a00",
---- 1485=>x"2e00", 1486=>x"2d00", 1487=>x"3a00", 1488=>x"3200", 1489=>x"3400", 1490=>x"3900", 1491=>x"3b00",
---- 1492=>x"3b00", 1493=>x"2e00", 1494=>x"2e00", 1495=>x"3b00", 1496=>x"3000", 1497=>x"3500", 1498=>x"4000",
---- 1499=>x"3800", 1500=>x"3900", 1501=>x"2d00", 1502=>x"3100", 1503=>x"3c00", 1504=>x"2f00", 1505=>x"3e00",
---- 1506=>x"4700", 1507=>x"3800", 1508=>x"3500", 1509=>x"2a00", 1510=>x"2f00", 1511=>x"3b00", 1512=>x"3200",
---- 1513=>x"3900", 1514=>x"c000", 1515=>x"3d00", 1516=>x"3800", 1517=>x"2d00", 1518=>x"3200", 1519=>x"3e00",
---- 1520=>x"3000", 1521=>x"3900", 1522=>x"3e00", 1523=>x"c000", 1524=>x"3400", 1525=>x"2d00", 1526=>x"3400",
---- 1527=>x"4300", 1528=>x"3600", 1529=>x"3d00", 1530=>x"4200", 1531=>x"4800", 1532=>x"3700", 1533=>x"2e00",
---- 1534=>x"3100", 1535=>x"4200", 1536=>x"3700", 1537=>x"3d00", 1538=>x"4800", 1539=>x"4a00", 1540=>x"3100",
---- 1541=>x"2d00", 1542=>x"3600", 1543=>x"4600", 1544=>x"3800", 1545=>x"4800", 1546=>x"b300", 1547=>x"4a00",
---- 1548=>x"2f00", 1549=>x"2800", 1550=>x"3100", 1551=>x"4b00", 1552=>x"3600", 1553=>x"4c00", 1554=>x"4d00",
---- 1555=>x"4c00", 1556=>x"2f00", 1557=>x"2900", 1558=>x"3200", 1559=>x"4200", 1560=>x"3400", 1561=>x"4500",
---- 1562=>x"4e00", 1563=>x"4700", 1564=>x"2900", 1565=>x"2600", 1566=>x"3800", 1567=>x"4800", 1568=>x"3a00",
---- 1569=>x"4600", 1570=>x"5500", 1571=>x"4300", 1572=>x"3000", 1573=>x"2a00", 1574=>x"4000", 1575=>x"5000",
---- 1576=>x"4200", 1577=>x"4600", 1578=>x"5800", 1579=>x"4000", 1580=>x"2e00", 1581=>x"2d00", 1582=>x"3a00",
---- 1583=>x"4a00", 1584=>x"c600", 1585=>x"4100", 1586=>x"5100", 1587=>x"3b00", 1588=>x"2c00", 1589=>x"2900",
---- 1590=>x"3b00", 1591=>x"5200", 1592=>x"3700", 1593=>x"4000", 1594=>x"ac00", 1595=>x"3800", 1596=>x"2c00",
---- 1597=>x"2c00", 1598=>x"3f00", 1599=>x"5300", 1600=>x"3700", 1601=>x"c000", 1602=>x"5100", 1603=>x"3600",
---- 1604=>x"2d00", 1605=>x"2700", 1606=>x"3d00", 1607=>x"5200", 1608=>x"3400", 1609=>x"4200", 1610=>x"4900",
---- 1611=>x"3400", 1612=>x"2b00", 1613=>x"2300", 1614=>x"4100", 1615=>x"4f00", 1616=>x"3100", 1617=>x"4400",
---- 1618=>x"4000", 1619=>x"3100", 1620=>x"2b00", 1621=>x"2700", 1622=>x"4200", 1623=>x"5400", 1624=>x"3000",
---- 1625=>x"3d00", 1626=>x"3e00", 1627=>x"3600", 1628=>x"3100", 1629=>x"2d00", 1630=>x"4600", 1631=>x"5200",
---- 1632=>x"5400", 1633=>x"3300", 1634=>x"3a00", 1635=>x"2f00", 1636=>x"2c00", 1637=>x"2a00", 1638=>x"bf00",
---- 1639=>x"5200", 1640=>x"8100", 1641=>x"2c00", 1642=>x"3300", 1643=>x"2c00", 1644=>x"2d00", 1645=>x"2900",
---- 1646=>x"3c00", 1647=>x"4e00", 1648=>x"9b00", 1649=>x"3f00", 1650=>x"2f00", 1651=>x"2e00", 1652=>x"3200",
---- 1653=>x"3100", 1654=>x"4200", 1655=>x"4e00", 1656=>x"9800", 1657=>x"6800", 1658=>x"d800", 1659=>x"3000",
---- 1660=>x"2f00", 1661=>x"2d00", 1662=>x"4300", 1663=>x"4f00", 1664=>x"8300", 1665=>x"9d00", 1666=>x"2200",
---- 1667=>x"2800", 1668=>x"2a00", 1669=>x"2400", 1670=>x"4400", 1671=>x"4c00", 1672=>x"6b00", 1673=>x"c000",
---- 1674=>x"2e00", 1675=>x"2200", 1676=>x"2b00", 1677=>x"2500", 1678=>x"3c00", 1679=>x"4800", 1680=>x"6600",
---- 1681=>x"c700", 1682=>x"3b00", 1683=>x"1d00", 1684=>x"2400", 1685=>x"2200", 1686=>x"3900", 1687=>x"4500",
---- 1688=>x"7700", 1689=>x"d300", 1690=>x"4f00", 1691=>x"2100", 1692=>x"2800", 1693=>x"2400", 1694=>x"3900",
---- 1695=>x"4700", 1696=>x"9d00", 1697=>x"cf00", 1698=>x"5e00", 1699=>x"1f00", 1700=>x"2900", 1701=>x"2200",
---- 1702=>x"3e00", 1703=>x"4800", 1704=>x"ba00", 1705=>x"c800", 1706=>x"4f00", 1707=>x"1d00", 1708=>x"2300",
---- 1709=>x"2100", 1710=>x"4300", 1711=>x"4000", 1712=>x"c200", 1713=>x"ba00", 1714=>x"3f00", 1715=>x"1f00",
---- 1716=>x"2a00", 1717=>x"2600", 1718=>x"4700", 1719=>x"4800", 1720=>x"c600", 1721=>x"9000", 1722=>x"2d00",
---- 1723=>x"2200", 1724=>x"2500", 1725=>x"2b00", 1726=>x"5200", 1727=>x"4800", 1728=>x"b500", 1729=>x"5700",
---- 1730=>x"5e00", 1731=>x"3900", 1732=>x"1d00", 1733=>x"2a00", 1734=>x"5300", 1735=>x"4500", 1736=>x"9800",
---- 1737=>x"6e00", 1738=>x"c100", 1739=>x"5500", 1740=>x"1b00", 1741=>x"3000", 1742=>x"4f00", 1743=>x"4000",
---- 1744=>x"9000", 1745=>x"8b00", 1746=>x"9d00", 1747=>x"3f00", 1748=>x"2100", 1749=>x"3400", 1750=>x"4900",
---- 1751=>x"3500", 1752=>x"4900", 1753=>x"2900", 1754=>x"2800", 1755=>x"2d00", 1756=>x"3f00", 1757=>x"3a00",
---- 1758=>x"4700", 1759=>x"3000", 1760=>x"5d00", 1761=>x"3000", 1762=>x"2500", 1763=>x"4f00", 1764=>x"3500",
---- 1765=>x"3900", 1766=>x"3e00", 1767=>x"3300", 1768=>x"b400", 1769=>x"8700", 1770=>x"7b00", 1771=>x"7700",
---- 1772=>x"3e00", 1773=>x"5300", 1774=>x"3f00", 1775=>x"2f00", 1776=>x"5400", 1777=>x"6000", 1778=>x"8100",
---- 1779=>x"7200", 1780=>x"8200", 1781=>x"8800", 1782=>x"7000", 1783=>x"6f00", 1784=>x"2200", 1785=>x"4000",
---- 1786=>x"2f00", 1787=>x"2000", 1788=>x"4c00", 1789=>x"5b00", 1790=>x"4e00", 1791=>x"7c00", 1792=>x"3000",
---- 1793=>x"4200", 1794=>x"1f00", 1795=>x"2800", 1796=>x"4300", 1797=>x"3a00", 1798=>x"2c00", 1799=>x"4100",
---- 1800=>x"2e00", 1801=>x"2f00", 1802=>x"2800", 1803=>x"3900", 1804=>x"4200", 1805=>x"3d00", 1806=>x"3200",
---- 1807=>x"4200", 1808=>x"2e00", 1809=>x"2400", 1810=>x"2c00", 1811=>x"4100", 1812=>x"3a00", 1813=>x"3000",
---- 1814=>x"2d00", 1815=>x"3f00", 1816=>x"7500", 1817=>x"3900", 1818=>x"2400", 1819=>x"3e00", 1820=>x"3b00",
---- 1821=>x"3400", 1822=>x"3200", 1823=>x"3c00", 1824=>x"a000", 1825=>x"3000", 1826=>x"2b00", 1827=>x"3400",
---- 1828=>x"ca00", 1829=>x"2b00", 1830=>x"3500", 1831=>x"3800", 1832=>x"6300", 1833=>x"2300", 1834=>x"3300",
---- 1835=>x"3700", 1836=>x"3100", 1837=>x"d400", 1838=>x"3b00", 1839=>x"3900", 1840=>x"2d00", 1841=>x"2900",
---- 1842=>x"3500", 1843=>x"3600", 1844=>x"2700", 1845=>x"2b00", 1846=>x"3b00", 1847=>x"3400", 1848=>x"2700",
---- 1849=>x"2f00", 1850=>x"3900", 1851=>x"3600", 1852=>x"2b00", 1853=>x"2e00", 1854=>x"2f00", 1855=>x"3100",
---- 1856=>x"2200", 1857=>x"3100", 1858=>x"3500", 1859=>x"2b00", 1860=>x"2900", 1861=>x"3400", 1862=>x"2f00",
---- 1863=>x"2f00", 1864=>x"2a00", 1865=>x"3100", 1866=>x"3100", 1867=>x"2400", 1868=>x"3000", 1869=>x"3500",
---- 1870=>x"2900", 1871=>x"2e00", 1872=>x"3900", 1873=>x"3800", 1874=>x"2c00", 1875=>x"2900", 1876=>x"3400",
---- 1877=>x"3000", 1878=>x"2800", 1879=>x"2c00", 1880=>x"3a00", 1881=>x"3400", 1882=>x"2b00", 1883=>x"2d00",
---- 1884=>x"3100", 1885=>x"2800", 1886=>x"2700", 1887=>x"2900", 1888=>x"3200", 1889=>x"2c00", 1890=>x"2f00",
---- 1891=>x"3200", 1892=>x"3200", 1893=>x"2a00", 1894=>x"2c00", 1895=>x"2a00", 1896=>x"2800", 1897=>x"2a00",
---- 1898=>x"2d00", 1899=>x"2f00", 1900=>x"2f00", 1901=>x"2b00", 1902=>x"2900", 1903=>x"2800", 1904=>x"2b00",
---- 1905=>x"2c00", 1906=>x"2b00", 1907=>x"2600", 1908=>x"2900", 1909=>x"2b00", 1910=>x"2600", 1911=>x"2a00",
---- 1912=>x"2b00", 1913=>x"2a00", 1914=>x"2c00", 1915=>x"2a00", 1916=>x"2b00", 1917=>x"2700", 1918=>x"2300",
---- 1919=>x"2a00", 1920=>x"2c00", 1921=>x"2b00", 1922=>x"2b00", 1923=>x"2e00", 1924=>x"2500", 1925=>x"2300",
---- 1926=>x"2500", 1927=>x"2f00", 1928=>x"3300", 1929=>x"2d00", 1930=>x"2a00", 1931=>x"2d00", 1932=>x"2800",
---- 1933=>x"2400", 1934=>x"2900", 1935=>x"2f00", 1936=>x"2e00", 1937=>x"2f00", 1938=>x"2900", 1939=>x"2800",
---- 1940=>x"2600", 1941=>x"2a00", 1942=>x"3100", 1943=>x"3200", 1944=>x"3300", 1945=>x"2a00", 1946=>x"2700",
---- 1947=>x"2700", 1948=>x"2300", 1949=>x"2500", 1950=>x"2a00", 1951=>x"3200", 1952=>x"2d00", 1953=>x"2700",
---- 1954=>x"2600", 1955=>x"2d00", 1956=>x"2b00", 1957=>x"2700", 1958=>x"2e00", 1959=>x"4000", 1960=>x"2a00",
---- 1961=>x"2f00", 1962=>x"2e00", 1963=>x"2a00", 1964=>x"2f00", 1965=>x"2f00", 1966=>x"3600", 1967=>x"3900",
---- 1968=>x"2900", 1969=>x"3100", 1970=>x"3100", 1971=>x"2c00", 1972=>x"2e00", 1973=>x"2d00", 1974=>x"2700",
---- 1975=>x"2900", 1976=>x"3000", 1977=>x"2c00", 1978=>x"2a00", 1979=>x"2900", 1980=>x"2800", 1981=>x"2800",
---- 1982=>x"2e00", 1983=>x"3300", 1984=>x"2b00", 1985=>x"2700", 1986=>x"2700", 1987=>x"2800", 1988=>x"3300",
---- 1989=>x"3600", 1990=>x"4000", 1991=>x"4a00", 1992=>x"2500", 1993=>x"2c00", 1994=>x"3200", 1995=>x"2f00",
---- 1996=>x"3400", 1997=>x"3a00", 1998=>x"4300", 1999=>x"5200", 2000=>x"3300", 2001=>x"2e00", 2002=>x"3100",
---- 2003=>x"3100", 2004=>x"3500", 2005=>x"4800", 2006=>x"5400", 2007=>x"5f00", 2008=>x"2f00", 2009=>x"3200",
---- 2010=>x"3400", 2011=>x"3700", 2012=>x"4700", 2013=>x"5500", 2014=>x"5d00", 2015=>x"6500", 2016=>x"2a00",
---- 2017=>x"3200", 2018=>x"3c00", 2019=>x"4b00", 2020=>x"5300", 2021=>x"5900", 2022=>x"6300", 2023=>x"9500",
---- 2024=>x"2b00", 2025=>x"3600", 2026=>x"4300", 2027=>x"4d00", 2028=>x"5700", 2029=>x"5b00", 2030=>x"6300",
---- 2031=>x"6800", 2032=>x"3900", 2033=>x"4b00", 2034=>x"5000", 2035=>x"5300", 2036=>x"5700", 2037=>x"5f00",
---- 2038=>x"6800", 2039=>x"6b00", 2040=>x"4500", 2041=>x"5400", 2042=>x"5100", 2043=>x"5a00", 2044=>x"5900",
---- 2045=>x"5f00", 2046=>x"6700", 2047=>x"6a00"),
---- 12 => (0=>x"8700", 1=>x"7900", 2=>x"8700", 3=>x"8700", 4=>x"8800", 5=>x"7a00", 6=>x"8800", 7=>x"8500",
---- 8=>x"8700", 9=>x"8600", 10=>x"8700", 11=>x"8800", 12=>x"8800", 13=>x"8600", 14=>x"8800",
---- 15=>x"8500", 16=>x"8700", 17=>x"8500", 18=>x"8700", 19=>x"8700", 20=>x"8700", 21=>x"8600",
---- 22=>x"8800", 23=>x"8500", 24=>x"8400", 25=>x"8600", 26=>x"8500", 27=>x"8400", 28=>x"8500",
---- 29=>x"8400", 30=>x"8400", 31=>x"8400", 32=>x"8500", 33=>x"8500", 34=>x"8300", 35=>x"8400",
---- 36=>x"8400", 37=>x"8200", 38=>x"8300", 39=>x"8200", 40=>x"8700", 41=>x"8400", 42=>x"8200",
---- 43=>x"8400", 44=>x"8300", 45=>x"8300", 46=>x"8400", 47=>x"8000", 48=>x"8200", 49=>x"8500",
---- 50=>x"8200", 51=>x"8300", 52=>x"8300", 53=>x"7d00", 54=>x"8400", 55=>x"8500", 56=>x"7f00",
---- 57=>x"8400", 58=>x"8400", 59=>x"8600", 60=>x"8400", 61=>x"8400", 62=>x"8400", 63=>x"8300",
---- 64=>x"8300", 65=>x"8300", 66=>x"8300", 67=>x"8600", 68=>x"8300", 69=>x"8100", 70=>x"8400",
---- 71=>x"8500", 72=>x"8500", 73=>x"8200", 74=>x"8200", 75=>x"8800", 76=>x"8600", 77=>x"8300",
---- 78=>x"8500", 79=>x"8500", 80=>x"8400", 81=>x"8100", 82=>x"8300", 83=>x"8600", 84=>x"8300",
---- 85=>x"8300", 86=>x"8100", 87=>x"8300", 88=>x"8200", 89=>x"8400", 90=>x"8100", 91=>x"8200",
---- 92=>x"8400", 93=>x"7f00", 94=>x"7f00", 95=>x"8400", 96=>x"8500", 97=>x"8400", 98=>x"8100",
---- 99=>x"8200", 100=>x"8200", 101=>x"8100", 102=>x"8000", 103=>x"8000", 104=>x"8a00", 105=>x"8600",
---- 106=>x"8500", 107=>x"8300", 108=>x"8300", 109=>x"7f00", 110=>x"7c00", 111=>x"7e00", 112=>x"8500",
---- 113=>x"8a00", 114=>x"8700", 115=>x"8300", 116=>x"8000", 117=>x"7b00", 118=>x"7c00", 119=>x"7e00",
---- 120=>x"8600", 121=>x"8400", 122=>x"7b00", 123=>x"8500", 124=>x"8200", 125=>x"8000", 126=>x"7d00",
---- 127=>x"7c00", 128=>x"8400", 129=>x"8300", 130=>x"8400", 131=>x"8100", 132=>x"8000", 133=>x"8200",
---- 134=>x"7f00", 135=>x"7c00", 136=>x"8500", 137=>x"8600", 138=>x"8400", 139=>x"8000", 140=>x"7d00",
---- 141=>x"7e00", 142=>x"7d00", 143=>x"7a00", 144=>x"7f00", 145=>x"8300", 146=>x"8100", 147=>x"7f00",
---- 148=>x"7b00", 149=>x"7f00", 150=>x"7e00", 151=>x"7c00", 152=>x"8400", 153=>x"7f00", 154=>x"7f00",
---- 155=>x"8100", 156=>x"7e00", 157=>x"7d00", 158=>x"7d00", 159=>x"7c00", 160=>x"8200", 161=>x"8100",
---- 162=>x"7d00", 163=>x"8000", 164=>x"7f00", 165=>x"7d00", 166=>x"7f00", 167=>x"7c00", 168=>x"8100",
---- 169=>x"8000", 170=>x"7e00", 171=>x"8000", 172=>x"7f00", 173=>x"7d00", 174=>x"8500", 175=>x"8100",
---- 176=>x"8200", 177=>x"8300", 178=>x"7e00", 179=>x"8000", 180=>x"7e00", 181=>x"7d00", 182=>x"7f00",
---- 183=>x"8100", 184=>x"8100", 185=>x"8800", 186=>x"8100", 187=>x"7b00", 188=>x"7d00", 189=>x"7b00",
---- 190=>x"7e00", 191=>x"7e00", 192=>x"7d00", 193=>x"7f00", 194=>x"8400", 195=>x"8600", 196=>x"8500",
---- 197=>x"8500", 198=>x"9200", 199=>x"7400", 200=>x"8100", 201=>x"8a00", 202=>x"8e00", 203=>x"9700",
---- 204=>x"9500", 205=>x"9600", 206=>x"9900", 207=>x"9b00", 208=>x"8f00", 209=>x"9500", 210=>x"9400",
---- 211=>x"9800", 212=>x"9500", 213=>x"8c00", 214=>x"9200", 215=>x"9400", 216=>x"8b00", 217=>x"8e00",
---- 218=>x"9300", 219=>x"9b00", 220=>x"8f00", 221=>x"8c00", 222=>x"8a00", 223=>x"9100", 224=>x"8a00",
---- 225=>x"9200", 226=>x"9400", 227=>x"9200", 228=>x"9100", 229=>x"9100", 230=>x"9000", 231=>x"9700",
---- 232=>x"8b00", 233=>x"9200", 234=>x"8e00", 235=>x"8e00", 236=>x"8b00", 237=>x"9300", 238=>x"9900",
---- 239=>x"9600", 240=>x"8900", 241=>x"8200", 242=>x"8400", 243=>x"8300", 244=>x"8d00", 245=>x"9500",
---- 246=>x"8d00", 247=>x"9300", 248=>x"8700", 249=>x"8100", 250=>x"7e00", 251=>x"8400", 252=>x"8f00",
---- 253=>x"8600", 254=>x"8600", 255=>x"8e00", 256=>x"8300", 257=>x"8200", 258=>x"7e00", 259=>x"8800",
---- 260=>x"7400", 261=>x"8a00", 262=>x"8900", 263=>x"8d00", 264=>x"8400", 265=>x"7e00", 266=>x"7f00",
---- 267=>x"8700", 268=>x"8700", 269=>x"8400", 270=>x"8b00", 271=>x"8700", 272=>x"7e00", 273=>x"8000",
---- 274=>x"8100", 275=>x"8200", 276=>x"8500", 277=>x"8900", 278=>x"8a00", 279=>x"8400", 280=>x"8000",
---- 281=>x"8600", 282=>x"8000", 283=>x"8600", 284=>x"8c00", 285=>x"8900", 286=>x"8100", 287=>x"8100",
---- 288=>x"8200", 289=>x"8900", 290=>x"8200", 291=>x"8b00", 292=>x"8c00", 293=>x"8200", 294=>x"7b00",
---- 295=>x"8700", 296=>x"8800", 297=>x"8700", 298=>x"8600", 299=>x"8c00", 300=>x"8100", 301=>x"8200",
---- 302=>x"8b00", 303=>x"8b00", 304=>x"8400", 305=>x"8100", 306=>x"8300", 307=>x"8800", 308=>x"8d00",
---- 309=>x"8b00", 310=>x"8d00", 311=>x"8800", 312=>x"8000", 313=>x"8000", 314=>x"7f00", 315=>x"8800",
---- 316=>x"8700", 317=>x"8400", 318=>x"8900", 319=>x"8100", 320=>x"7e00", 321=>x"7900", 322=>x"8100",
---- 323=>x"8500", 324=>x"8300", 325=>x"8600", 326=>x"8800", 327=>x"8a00", 328=>x"7f00", 329=>x"7e00",
---- 330=>x"8000", 331=>x"8700", 332=>x"8200", 333=>x"8100", 334=>x"8200", 335=>x"8400", 336=>x"8100",
---- 337=>x"8200", 338=>x"8600", 339=>x"8900", 340=>x"8a00", 341=>x"8700", 342=>x"7600", 343=>x"8700",
---- 344=>x"8500", 345=>x"8200", 346=>x"7c00", 347=>x"8e00", 348=>x"8900", 349=>x"8700", 350=>x"8c00",
---- 351=>x"8700", 352=>x"8000", 353=>x"8200", 354=>x"8700", 355=>x"8d00", 356=>x"8800", 357=>x"8200",
---- 358=>x"8900", 359=>x"8800", 360=>x"7c00", 361=>x"8700", 362=>x"8b00", 363=>x"8700", 364=>x"8100",
---- 365=>x"7400", 366=>x"8b00", 367=>x"8b00", 368=>x"8100", 369=>x"8c00", 370=>x"8d00", 371=>x"8900",
---- 372=>x"9100", 373=>x"8b00", 374=>x"8c00", 375=>x"8c00", 376=>x"8800", 377=>x"8a00", 378=>x"7200",
---- 379=>x"8a00", 380=>x"8a00", 381=>x"9000", 382=>x"9000", 383=>x"9000", 384=>x"8400", 385=>x"8700",
---- 386=>x"8200", 387=>x"8500", 388=>x"8f00", 389=>x"8c00", 390=>x"9000", 391=>x"9100", 392=>x"8d00",
---- 393=>x"8900", 394=>x"8700", 395=>x"8c00", 396=>x"8200", 397=>x"9000", 398=>x"8800", 399=>x"8e00",
---- 400=>x"8a00", 401=>x"8e00", 402=>x"8900", 403=>x"8700", 404=>x"7100", 405=>x"8f00", 406=>x"8c00",
---- 407=>x"8d00", 408=>x"8f00", 409=>x"8800", 410=>x"8d00", 411=>x"8c00", 412=>x"8600", 413=>x"8f00",
---- 414=>x"8800", 415=>x"8c00", 416=>x"8d00", 417=>x"8a00", 418=>x"8c00", 419=>x"8e00", 420=>x"8e00",
---- 421=>x"8700", 422=>x"8b00", 423=>x"8900", 424=>x"8600", 425=>x"8400", 426=>x"8c00", 427=>x"9000",
---- 428=>x"9100", 429=>x"8b00", 430=>x"9000", 431=>x"8b00", 432=>x"7b00", 433=>x"8c00", 434=>x"8700",
---- 435=>x"8c00", 436=>x"8f00", 437=>x"8900", 438=>x"8c00", 439=>x"8500", 440=>x"8a00", 441=>x"8200",
---- 442=>x"8c00", 443=>x"8c00", 444=>x"8900", 445=>x"8d00", 446=>x"8300", 447=>x"8100", 448=>x"8600",
---- 449=>x"8a00", 450=>x"8a00", 451=>x"8800", 452=>x"9000", 453=>x"8800", 454=>x"8600", 455=>x"7c00",
---- 456=>x"8400", 457=>x"8200", 458=>x"8b00", 459=>x"8e00", 460=>x"8a00", 461=>x"7700", 462=>x"7900",
---- 463=>x"7f00", 464=>x"8400", 465=>x"8b00", 466=>x"8d00", 467=>x"8200", 468=>x"7300", 469=>x"7100",
---- 470=>x"7900", 471=>x"7200", 472=>x"8b00", 473=>x"8b00", 474=>x"7f00", 475=>x"7300", 476=>x"7600",
---- 477=>x"7100", 478=>x"6400", 479=>x"7200", 480=>x"8800", 481=>x"7c00", 482=>x"8100", 483=>x"7e00",
---- 484=>x"7100", 485=>x"6500", 486=>x"7400", 487=>x"9d00", 488=>x"8000", 489=>x"7d00", 490=>x"7900",
---- 491=>x"6f00", 492=>x"6800", 493=>x"7e00", 494=>x"9f00", 495=>x"a300", 496=>x"7a00", 497=>x"7100",
---- 498=>x"6d00", 499=>x"6200", 500=>x"8100", 501=>x"a700", 502=>x"ac00", 503=>x"a800", 504=>x"7100",
---- 505=>x"6f00", 506=>x"6b00", 507=>x"8100", 508=>x"a100", 509=>x"ab00", 510=>x"ae00", 511=>x"b600",
---- 512=>x"6b00", 513=>x"6900", 514=>x"8e00", 515=>x"a300", 516=>x"9f00", 517=>x"ac00", 518=>x"b200",
---- 519=>x"ad00", 520=>x"6c00", 521=>x"8600", 522=>x"9e00", 523=>x"ab00", 524=>x"a600", 525=>x"a700",
---- 526=>x"a400", 527=>x"a000", 528=>x"9500", 529=>x"a300", 530=>x"9600", 531=>x"a400", 532=>x"b300",
---- 533=>x"9d00", 534=>x"9000", 535=>x"9900", 536=>x"9c00", 537=>x"a300", 538=>x"a400", 539=>x"9700",
---- 540=>x"9600", 541=>x"9e00", 542=>x"9200", 543=>x"9600", 544=>x"9c00", 545=>x"9d00", 546=>x"a100",
---- 547=>x"9400", 548=>x"8900", 549=>x"8d00", 550=>x"a600", 551=>x"a000", 552=>x"a400", 553=>x"9400",
---- 554=>x"9300", 555=>x"9200", 556=>x"9500", 557=>x"9a00", 558=>x"9000", 559=>x"8b00", 560=>x"9a00",
---- 561=>x"9100", 562=>x"8d00", 563=>x"9700", 564=>x"a600", 565=>x"8d00", 566=>x"7e00", 567=>x"9900",
---- 568=>x"9000", 569=>x"8c00", 570=>x"9b00", 571=>x"9700", 572=>x"8500", 573=>x"8200", 574=>x"9b00",
---- 575=>x"a000", 576=>x"8b00", 577=>x"9700", 578=>x"9a00", 579=>x"8000", 580=>x"8200", 581=>x"9900",
---- 582=>x"a000", 583=>x"9d00", 584=>x"9000", 585=>x"9700", 586=>x"7f00", 587=>x"8000", 588=>x"9800",
---- 589=>x"9500", 590=>x"9400", 591=>x"a200", 592=>x"8a00", 593=>x"7400", 594=>x"8300", 595=>x"9400",
---- 596=>x"9200", 597=>x"9600", 598=>x"9700", 599=>x"9800", 600=>x"7b00", 601=>x"8900", 602=>x"9800",
---- 603=>x"9200", 604=>x"9300", 605=>x"9200", 606=>x"5f00", 607=>x"9500", 608=>x"8500", 609=>x"9600",
---- 610=>x"9800", 611=>x"9600", 612=>x"9800", 613=>x"9b00", 614=>x"9d00", 615=>x"8900", 616=>x"9400",
---- 617=>x"9100", 618=>x"9300", 619=>x"9800", 620=>x"9a00", 621=>x"9a00", 622=>x"8e00", 623=>x"8500",
---- 624=>x"9500", 625=>x"9400", 626=>x"9100", 627=>x"9b00", 628=>x"9700", 629=>x"9500", 630=>x"9000",
---- 631=>x"8f00", 632=>x"9400", 633=>x"9a00", 634=>x"9400", 635=>x"8f00", 636=>x"8f00", 637=>x"8c00",
---- 638=>x"9a00", 639=>x"9e00", 640=>x"9a00", 641=>x"9400", 642=>x"6e00", 643=>x"8900", 644=>x"8d00",
---- 645=>x"9800", 646=>x"9500", 647=>x"9800", 648=>x"9400", 649=>x"9000", 650=>x"8600", 651=>x"9400",
---- 652=>x"8a00", 653=>x"8f00", 654=>x"8900", 655=>x"8a00", 656=>x"8600", 657=>x"8c00", 658=>x"9000",
---- 659=>x"8f00", 660=>x"8700", 661=>x"8300", 662=>x"9100", 663=>x"9200", 664=>x"8600", 665=>x"9300",
---- 666=>x"8a00", 667=>x"7c00", 668=>x"8200", 669=>x"9200", 670=>x"9800", 671=>x"9900", 672=>x"8f00",
---- 673=>x"8200", 674=>x"7400", 675=>x"8100", 676=>x"8f00", 677=>x"9600", 678=>x"9300", 679=>x"9800",
---- 680=>x"7f00", 681=>x"7d00", 682=>x"8400", 683=>x"8600", 684=>x"9600", 685=>x"9b00", 686=>x"9100",
---- 687=>x"8000", 688=>x"7b00", 689=>x"8a00", 690=>x"8b00", 691=>x"8500", 692=>x"8e00", 693=>x"9700",
---- 694=>x"8100", 695=>x"8900", 696=>x"8200", 697=>x"8500", 698=>x"8d00", 699=>x"9800", 700=>x"8600",
---- 701=>x"7d00", 702=>x"8800", 703=>x"9500", 704=>x"8300", 705=>x"8700", 706=>x"8a00", 707=>x"9100",
---- 708=>x"8200", 709=>x"8000", 710=>x"9300", 711=>x"9400", 712=>x"8700", 713=>x"8500", 714=>x"8600",
---- 715=>x"8000", 716=>x"8100", 717=>x"9300", 718=>x"8b00", 719=>x"8d00", 720=>x"8900", 721=>x"8500",
---- 722=>x"7a00", 723=>x"7f00", 724=>x"8e00", 725=>x"9600", 726=>x"8d00", 727=>x"8b00", 728=>x"8800",
---- 729=>x"8300", 730=>x"7c00", 731=>x"8b00", 732=>x"8f00", 733=>x"8c00", 734=>x"8c00", 735=>x"7100",
---- 736=>x"7c00", 737=>x"7b00", 738=>x"8700", 739=>x"8e00", 740=>x"8900", 741=>x"8900", 742=>x"8f00",
---- 743=>x"7400", 744=>x"7a00", 745=>x"8200", 746=>x"8a00", 747=>x"8b00", 748=>x"8a00", 749=>x"8300",
---- 750=>x"7700", 751=>x"6c00", 752=>x"8400", 753=>x"8f00", 754=>x"8a00", 755=>x"8c00", 756=>x"8800",
---- 757=>x"7100", 758=>x"6900", 759=>x"7c00", 760=>x"9300", 761=>x"8a00", 762=>x"8600", 763=>x"8600",
---- 764=>x"8500", 765=>x"6300", 766=>x"7200", 767=>x"8b00", 768=>x"8a00", 769=>x"8800", 770=>x"8a00",
---- 771=>x"8600", 772=>x"8900", 773=>x"6600", 774=>x"7400", 775=>x"8b00", 776=>x"8300", 777=>x"8800",
---- 778=>x"8900", 779=>x"8d00", 780=>x"9200", 781=>x"6c00", 782=>x"7200", 783=>x"8700", 784=>x"6600",
---- 785=>x"6e00", 786=>x"8100", 787=>x"9300", 788=>x"9100", 789=>x"6d00", 790=>x"9d00", 791=>x"5d00",
---- 792=>x"7500", 793=>x"6300", 794=>x"5b00", 795=>x"6d00", 796=>x"7f00", 797=>x"9000", 798=>x"4800",
---- 799=>x"3a00", 800=>x"7800", 801=>x"6100", 802=>x"6200", 803=>x"5900", 804=>x"4a00", 805=>x"5600",
---- 806=>x"4c00", 807=>x"4400", 808=>x"6500", 809=>x"3b00", 810=>x"3b00", 811=>x"4500", 812=>x"4800",
---- 813=>x"4f00", 814=>x"4a00", 815=>x"4e00", 816=>x"6d00", 817=>x"6500", 818=>x"5700", 819=>x"5000",
---- 820=>x"4b00", 821=>x"3d00", 822=>x"4300", 823=>x"5d00", 824=>x"6600", 825=>x"5f00", 826=>x"5f00",
---- 827=>x"ae00", 828=>x"4400", 829=>x"4800", 830=>x"5f00", 831=>x"5e00", 832=>x"3e00", 833=>x"5400",
---- 834=>x"4b00", 835=>x"4d00", 836=>x"5500", 837=>x"5d00", 838=>x"6500", 839=>x"5300", 840=>x"4a00",
---- 841=>x"4700", 842=>x"4b00", 843=>x"5700", 844=>x"4e00", 845=>x"6300", 846=>x"5b00", 847=>x"4400",
---- 848=>x"4800", 849=>x"3a00", 850=>x"3d00", 851=>x"4400", 852=>x"4600", 853=>x"5e00", 854=>x"5400",
---- 855=>x"4800", 856=>x"bd00", 857=>x"3900", 858=>x"3500", 859=>x"2e00", 860=>x"4200", 861=>x"5600",
---- 862=>x"4c00", 863=>x"4300", 864=>x"3800", 865=>x"3200", 866=>x"2a00", 867=>x"2c00", 868=>x"3200",
---- 869=>x"4900", 870=>x"4d00", 871=>x"4400", 872=>x"2c00", 873=>x"2f00", 874=>x"2e00", 875=>x"3000",
---- 876=>x"2d00", 877=>x"4900", 878=>x"5900", 879=>x"3f00", 880=>x"2e00", 881=>x"2c00", 882=>x"2e00",
---- 883=>x"3200", 884=>x"2e00", 885=>x"3700", 886=>x"5900", 887=>x"4b00", 888=>x"2b00", 889=>x"2f00",
---- 890=>x"2f00", 891=>x"2e00", 892=>x"3100", 893=>x"3100", 894=>x"3c00", 895=>x"5300", 896=>x"2700",
---- 897=>x"3600", 898=>x"3300", 899=>x"3700", 900=>x"3300", 901=>x"2f00", 902=>x"2e00", 903=>x"4100",
---- 904=>x"2d00", 905=>x"4300", 906=>x"3a00", 907=>x"3900", 908=>x"3000", 909=>x"2e00", 910=>x"3400",
---- 911=>x"3300", 912=>x"c100", 913=>x"4600", 914=>x"3100", 915=>x"3900", 916=>x"2e00", 917=>x"3400",
---- 918=>x"3b00", 919=>x"3000", 920=>x"3e00", 921=>x"3300", 922=>x"3a00", 923=>x"3800", 924=>x"2c00",
---- 925=>x"3600", 926=>x"3800", 927=>x"2f00", 928=>x"2d00", 929=>x"3300", 930=>x"4000", 931=>x"3000",
---- 932=>x"cd00", 933=>x"3900", 934=>x"3400", 935=>x"3200", 936=>x"2f00", 937=>x"4d00", 938=>x"4600",
---- 939=>x"2c00", 940=>x"3400", 941=>x"3700", 942=>x"2a00", 943=>x"3800", 944=>x"3d00", 945=>x"5700",
---- 946=>x"3600", 947=>x"2c00", 948=>x"3300", 949=>x"3300", 950=>x"2700", 951=>x"4300", 952=>x"6500",
---- 953=>x"4700", 954=>x"2f00", 955=>x"2600", 956=>x"3600", 957=>x"3100", 958=>x"2600", 959=>x"5000",
---- 960=>x"4900", 961=>x"3a00", 962=>x"2900", 963=>x"2800", 964=>x"3700", 965=>x"2d00", 966=>x"2800",
---- 967=>x"5a00", 968=>x"4300", 969=>x"3200", 970=>x"2a00", 971=>x"2c00", 972=>x"3800", 973=>x"3000",
---- 974=>x"3400", 975=>x"5800", 976=>x"2c00", 977=>x"2800", 978=>x"2900", 979=>x"2c00", 980=>x"3200",
---- 981=>x"3100", 982=>x"3800", 983=>x"4300", 984=>x"2d00", 985=>x"2b00", 986=>x"3300", 987=>x"3300",
---- 988=>x"2f00", 989=>x"3800", 990=>x"3e00", 991=>x"4000", 992=>x"3c00", 993=>x"2b00", 994=>x"3600",
---- 995=>x"2e00", 996=>x"2b00", 997=>x"3000", 998=>x"4600", 999=>x"6200", 1000=>x"4d00", 1001=>x"2d00",
---- 1002=>x"3600", 1003=>x"2700", 1004=>x"2800", 1005=>x"2200", 1006=>x"2700", 1007=>x"5200", 1008=>x"6000",
---- 1009=>x"4200", 1010=>x"2c00", 1011=>x"2400", 1012=>x"2900", 1013=>x"2800", 1014=>x"2700", 1015=>x"3300",
---- 1016=>x"6900", 1017=>x"5500", 1018=>x"2500", 1019=>x"2600", 1020=>x"2700", 1021=>x"2e00", 1022=>x"2b00",
---- 1023=>x"2800", 1024=>x"5800", 1025=>x"6700", 1026=>x"3200", 1027=>x"2600", 1028=>x"2a00", 1029=>x"d100",
---- 1030=>x"2e00", 1031=>x"2c00", 1032=>x"3500", 1033=>x"6e00", 1034=>x"6200", 1035=>x"3100", 1036=>x"2500",
---- 1037=>x"2c00", 1038=>x"2f00", 1039=>x"3000", 1040=>x"2200", 1041=>x"4100", 1042=>x"7a00", 1043=>x"6e00",
---- 1044=>x"4300", 1045=>x"2200", 1046=>x"2300", 1047=>x"2d00", 1048=>x"2800", 1049=>x"2500", 1050=>x"4700",
---- 1051=>x"7600", 1052=>x"6900", 1053=>x"4c00", 1054=>x"3500", 1055=>x"2700", 1056=>x"d400", 1057=>x"2b00",
---- 1058=>x"2e00", 1059=>x"3e00", 1060=>x"3500", 1061=>x"4400", 1062=>x"5800", 1063=>x"3600", 1064=>x"2900",
---- 1065=>x"2c00", 1066=>x"3200", 1067=>x"3000", 1068=>x"2700", 1069=>x"2b00", 1070=>x"3900", 1071=>x"2e00",
---- 1072=>x"2b00", 1073=>x"2b00", 1074=>x"3400", 1075=>x"3200", 1076=>x"2700", 1077=>x"2c00", 1078=>x"2a00",
---- 1079=>x"2400", 1080=>x"2e00", 1081=>x"2a00", 1082=>x"3300", 1083=>x"3100", 1084=>x"2800", 1085=>x"2500",
---- 1086=>x"2600", 1087=>x"2c00", 1088=>x"2b00", 1089=>x"2a00", 1090=>x"2f00", 1091=>x"3100", 1092=>x"2600",
---- 1093=>x"2700", 1094=>x"2200", 1095=>x"2c00", 1096=>x"2e00", 1097=>x"2f00", 1098=>x"3600", 1099=>x"cd00",
---- 1100=>x"2700", 1101=>x"2500", 1102=>x"2300", 1103=>x"2800", 1104=>x"2f00", 1105=>x"3300", 1106=>x"3200",
---- 1107=>x"2c00", 1108=>x"2300", 1109=>x"2300", 1110=>x"1b00", 1111=>x"4200", 1112=>x"3300", 1113=>x"3500",
---- 1114=>x"2c00", 1115=>x"2600", 1116=>x"2400", 1117=>x"2000", 1118=>x"2600", 1119=>x"7a00", 1120=>x"3200",
---- 1121=>x"3400", 1122=>x"2f00", 1123=>x"2400", 1124=>x"2100", 1125=>x"1c00", 1126=>x"5700", 1127=>x"9900",
---- 1128=>x"2e00", 1129=>x"2d00", 1130=>x"2900", 1131=>x"2500", 1132=>x"1f00", 1133=>x"2f00", 1134=>x"8a00",
---- 1135=>x"8700", 1136=>x"2c00", 1137=>x"2e00", 1138=>x"2900", 1139=>x"2400", 1140=>x"2200", 1141=>x"6200",
---- 1142=>x"9800", 1143=>x"6600", 1144=>x"3100", 1145=>x"3300", 1146=>x"2f00", 1147=>x"2700", 1148=>x"3c00",
---- 1149=>x"9000", 1150=>x"7700", 1151=>x"6200", 1152=>x"3400", 1153=>x"3000", 1154=>x"3000", 1155=>x"2400",
---- 1156=>x"6f00", 1157=>x"9400", 1158=>x"6200", 1159=>x"8400", 1160=>x"2e00", 1161=>x"2d00", 1162=>x"2600",
---- 1163=>x"4400", 1164=>x"9800", 1165=>x"7400", 1166=>x"6400", 1167=>x"a300", 1168=>x"2d00", 1169=>x"2a00",
---- 1170=>x"2500", 1171=>x"7200", 1172=>x"9600", 1173=>x"6400", 1174=>x"7e00", 1175=>x"b600", 1176=>x"2b00",
---- 1177=>x"2800", 1178=>x"4300", 1179=>x"9100", 1180=>x"7d00", 1181=>x"6f00", 1182=>x"9500", 1183=>x"b500",
---- 1184=>x"2400", 1185=>x"2a00", 1186=>x"7700", 1187=>x"9300", 1188=>x"6d00", 1189=>x"8200", 1190=>x"bb00",
---- 1191=>x"b700", 1192=>x"1e00", 1193=>x"4300", 1194=>x"9400", 1195=>x"7b00", 1196=>x"6f00", 1197=>x"a200",
---- 1198=>x"c600", 1199=>x"be00", 1200=>x"2100", 1201=>x"7200", 1202=>x"8f00", 1203=>x"6b00", 1204=>x"7b00",
---- 1205=>x"bc00", 1206=>x"bd00", 1207=>x"c200", 1208=>x"3e00", 1209=>x"7200", 1210=>x"7600", 1211=>x"6f00",
---- 1212=>x"9a00", 1213=>x"c200", 1214=>x"c000", 1215=>x"cb00", 1216=>x"6300", 1217=>x"8f00", 1218=>x"6600",
---- 1219=>x"7800", 1220=>x"b800", 1221=>x"c800", 1222=>x"c700", 1223=>x"da00", 1224=>x"8700", 1225=>x"8000",
---- 1226=>x"6900", 1227=>x"9200", 1228=>x"ca00", 1229=>x"ca00", 1230=>x"d000", 1231=>x"c000", 1232=>x"9600",
---- 1233=>x"6f00", 1234=>x"7200", 1235=>x"aa00", 1236=>x"cb00", 1237=>x"cb00", 1238=>x"3100", 1239=>x"5b00",
---- 1240=>x"8100", 1241=>x"7000", 1242=>x"8400", 1243=>x"c100", 1244=>x"ca00", 1245=>x"d500", 1246=>x"8200",
---- 1247=>x"1d00", 1248=>x"7300", 1249=>x"7300", 1250=>x"a600", 1251=>x"d300", 1252=>x"d400", 1253=>x"a700",
---- 1254=>x"2800", 1255=>x"2400", 1256=>x"7600", 1257=>x"8800", 1258=>x"c900", 1259=>x"bd00", 1260=>x"a700",
---- 1261=>x"5300", 1262=>x"1900", 1263=>x"2500", 1264=>x"6400", 1265=>x"8800", 1266=>x"ac00", 1267=>x"9700",
---- 1268=>x"9200", 1269=>x"4f00", 1270=>x"2700", 1271=>x"2100", 1272=>x"7e00", 1273=>x"7d00", 1274=>x"9900",
---- 1275=>x"b400", 1276=>x"8b00", 1277=>x"3500", 1278=>x"2100", 1279=>x"2700", 1280=>x"ae00", 1281=>x"b200",
---- 1282=>x"be00", 1283=>x"9600", 1284=>x"4a00", 1285=>x"2500", 1286=>x"2200", 1287=>x"2700", 1288=>x"b700",
---- 1289=>x"b400", 1290=>x"9400", 1291=>x"4400", 1292=>x"2700", 1293=>x"2100", 1294=>x"2200", 1295=>x"2700",
---- 1296=>x"c500", 1297=>x"a700", 1298=>x"3b00", 1299=>x"1f00", 1300=>x"2700", 1301=>x"2400", 1302=>x"2500",
---- 1303=>x"2b00", 1304=>x"be00", 1305=>x"6c00", 1306=>x"1d00", 1307=>x"2600", 1308=>x"2b00", 1309=>x"2b00",
---- 1310=>x"d300", 1311=>x"2c00", 1312=>x"6b00", 1313=>x"2100", 1314=>x"2500", 1315=>x"2500", 1316=>x"3a00",
---- 1317=>x"4900", 1318=>x"3f00", 1319=>x"2f00", 1320=>x"2900", 1321=>x"2500", 1322=>x"2800", 1323=>x"2a00",
---- 1324=>x"3400", 1325=>x"4100", 1326=>x"3c00", 1327=>x"3000", 1328=>x"2800", 1329=>x"3300", 1330=>x"3300",
---- 1331=>x"3100", 1332=>x"3400", 1333=>x"3700", 1334=>x"3a00", 1335=>x"3500", 1336=>x"3200", 1337=>x"3700",
---- 1338=>x"3a00", 1339=>x"3500", 1340=>x"3700", 1341=>x"3a00", 1342=>x"3e00", 1343=>x"3900", 1344=>x"2c00",
---- 1345=>x"2d00", 1346=>x"3100", 1347=>x"3400", 1348=>x"3300", 1349=>x"3800", 1350=>x"4100", 1351=>x"3f00",
---- 1352=>x"3500", 1353=>x"2e00", 1354=>x"2f00", 1355=>x"3100", 1356=>x"2d00", 1357=>x"3300", 1358=>x"4300",
---- 1359=>x"3d00", 1360=>x"3700", 1361=>x"3a00", 1362=>x"3000", 1363=>x"3300", 1364=>x"2e00", 1365=>x"3700",
---- 1366=>x"4300", 1367=>x"4400", 1368=>x"3400", 1369=>x"3400", 1370=>x"2f00", 1371=>x"3500", 1372=>x"3300",
---- 1373=>x"3400", 1374=>x"4300", 1375=>x"4a00", 1376=>x"3800", 1377=>x"3200", 1378=>x"2a00", 1379=>x"3400",
---- 1380=>x"3200", 1381=>x"3300", 1382=>x"3f00", 1383=>x"4e00", 1384=>x"3500", 1385=>x"2d00", 1386=>x"2b00",
---- 1387=>x"3300", 1388=>x"3600", 1389=>x"3700", 1390=>x"4400", 1391=>x"4b00", 1392=>x"3300", 1393=>x"2b00",
---- 1394=>x"2e00", 1395=>x"3000", 1396=>x"3400", 1397=>x"3c00", 1398=>x"ba00", 1399=>x"4500", 1400=>x"3f00",
---- 1401=>x"2700", 1402=>x"2f00", 1403=>x"2d00", 1404=>x"3200", 1405=>x"3b00", 1406=>x"3a00", 1407=>x"4400",
---- 1408=>x"4300", 1409=>x"2d00", 1410=>x"2f00", 1411=>x"3100", 1412=>x"3500", 1413=>x"3900", 1414=>x"3a00",
---- 1415=>x"3e00", 1416=>x"3e00", 1417=>x"3000", 1418=>x"2c00", 1419=>x"ca00", 1420=>x"3b00", 1421=>x"3c00",
---- 1422=>x"c200", 1423=>x"3900", 1424=>x"c600", 1425=>x"3400", 1426=>x"2b00", 1427=>x"3000", 1428=>x"3d00",
---- 1429=>x"3800", 1430=>x"3d00", 1431=>x"3900", 1432=>x"3700", 1433=>x"3700", 1434=>x"3100", 1435=>x"2d00",
---- 1436=>x"3400", 1437=>x"3900", 1438=>x"3c00", 1439=>x"3d00", 1440=>x"3500", 1441=>x"3600", 1442=>x"3400",
---- 1443=>x"3100", 1444=>x"3100", 1445=>x"4000", 1446=>x"3a00", 1447=>x"3b00", 1448=>x"3600", 1449=>x"3100",
---- 1450=>x"3500", 1451=>x"3700", 1452=>x"3500", 1453=>x"3800", 1454=>x"3f00", 1455=>x"3b00", 1456=>x"3600",
---- 1457=>x"3300", 1458=>x"3500", 1459=>x"3e00", 1460=>x"3e00", 1461=>x"3800", 1462=>x"4200", 1463=>x"3d00",
---- 1464=>x"3200", 1465=>x"3200", 1466=>x"3700", 1467=>x"c900", 1468=>x"3c00", 1469=>x"3f00", 1470=>x"3700",
---- 1471=>x"3e00", 1472=>x"3500", 1473=>x"3400", 1474=>x"3500", 1475=>x"3300", 1476=>x"3900", 1477=>x"3b00",
---- 1478=>x"3900", 1479=>x"3900", 1480=>x"3200", 1481=>x"3300", 1482=>x"3500", 1483=>x"3100", 1484=>x"3200",
---- 1485=>x"3800", 1486=>x"c300", 1487=>x"3800", 1488=>x"3200", 1489=>x"3400", 1490=>x"3900", 1491=>x"3000",
---- 1492=>x"2f00", 1493=>x"2f00", 1494=>x"3a00", 1495=>x"3800", 1496=>x"3400", 1497=>x"cf00", 1498=>x"3800",
---- 1499=>x"3100", 1500=>x"2b00", 1501=>x"2f00", 1502=>x"3300", 1503=>x"3900", 1504=>x"3500", 1505=>x"2d00",
---- 1506=>x"3500", 1507=>x"3800", 1508=>x"2e00", 1509=>x"3200", 1510=>x"3100", 1511=>x"cc00", 1512=>x"3300",
---- 1513=>x"3100", 1514=>x"3100", 1515=>x"3a00", 1516=>x"3100", 1517=>x"2d00", 1518=>x"3100", 1519=>x"3100",
---- 1520=>x"3400", 1521=>x"3200", 1522=>x"3200", 1523=>x"3a00", 1524=>x"3800", 1525=>x"2d00", 1526=>x"3000",
---- 1527=>x"2f00", 1528=>x"3400", 1529=>x"3000", 1530=>x"3700", 1531=>x"3500", 1532=>x"3700", 1533=>x"3000",
---- 1534=>x"3200", 1535=>x"3400", 1536=>x"3600", 1537=>x"3000", 1538=>x"3300", 1539=>x"3600", 1540=>x"3a00",
---- 1541=>x"3400", 1542=>x"3100", 1543=>x"3500", 1544=>x"3300", 1545=>x"3100", 1546=>x"3200", 1547=>x"3000",
---- 1548=>x"3a00", 1549=>x"3200", 1550=>x"2f00", 1551=>x"3400", 1552=>x"3300", 1553=>x"3100", 1554=>x"3300",
---- 1555=>x"2f00", 1556=>x"3600", 1557=>x"3500", 1558=>x"2e00", 1559=>x"3400", 1560=>x"3000", 1561=>x"3000",
---- 1562=>x"3000", 1563=>x"cf00", 1564=>x"3500", 1565=>x"3500", 1566=>x"2f00", 1567=>x"3200", 1568=>x"2e00",
---- 1569=>x"3000", 1570=>x"3400", 1571=>x"3000", 1572=>x"3300", 1573=>x"3900", 1574=>x"cd00", 1575=>x"2f00",
---- 1576=>x"3800", 1577=>x"3300", 1578=>x"3800", 1579=>x"3200", 1580=>x"2e00", 1581=>x"3200", 1582=>x"3600",
---- 1583=>x"3400", 1584=>x"3600", 1585=>x"3000", 1586=>x"3800", 1587=>x"3200", 1588=>x"d100", 1589=>x"2f00",
---- 1590=>x"3900", 1591=>x"3600", 1592=>x"3000", 1593=>x"3000", 1594=>x"3600", 1595=>x"2e00", 1596=>x"3000",
---- 1597=>x"2c00", 1598=>x"3600", 1599=>x"3700", 1600=>x"3000", 1601=>x"2f00", 1602=>x"3300", 1603=>x"2d00",
---- 1604=>x"3000", 1605=>x"2d00", 1606=>x"3700", 1607=>x"3900", 1608=>x"3200", 1609=>x"3100", 1610=>x"3800",
---- 1611=>x"3000", 1612=>x"3000", 1613=>x"2b00", 1614=>x"3400", 1615=>x"3b00", 1616=>x"3600", 1617=>x"3300",
---- 1618=>x"c700", 1619=>x"3600", 1620=>x"3500", 1621=>x"2f00", 1622=>x"3300", 1623=>x"3700", 1624=>x"3900",
---- 1625=>x"3700", 1626=>x"3900", 1627=>x"3400", 1628=>x"3100", 1629=>x"3000", 1630=>x"3500", 1631=>x"3800",
---- 1632=>x"3900", 1633=>x"3400", 1634=>x"3800", 1635=>x"3500", 1636=>x"3500", 1637=>x"2f00", 1638=>x"3200",
---- 1639=>x"3500", 1640=>x"3500", 1641=>x"3500", 1642=>x"3400", 1643=>x"3400", 1644=>x"3700", 1645=>x"3300",
---- 1646=>x"3500", 1647=>x"3400", 1648=>x"3900", 1649=>x"3800", 1650=>x"3900", 1651=>x"3a00", 1652=>x"3900",
---- 1653=>x"3500", 1654=>x"3700", 1655=>x"3a00", 1656=>x"3c00", 1657=>x"3f00", 1658=>x"3900", 1659=>x"3400",
---- 1660=>x"3500", 1661=>x"3000", 1662=>x"3100", 1663=>x"3900", 1664=>x"3500", 1665=>x"3b00", 1666=>x"3600",
---- 1667=>x"2e00", 1668=>x"3300", 1669=>x"2b00", 1670=>x"3200", 1671=>x"3400", 1672=>x"3900", 1673=>x"3a00",
---- 1674=>x"3800", 1675=>x"3500", 1676=>x"3400", 1677=>x"2f00", 1678=>x"3200", 1679=>x"3400", 1680=>x"3a00",
---- 1681=>x"3e00", 1682=>x"3700", 1683=>x"3200", 1684=>x"3200", 1685=>x"2b00", 1686=>x"2d00", 1687=>x"3100",
---- 1688=>x"3600", 1689=>x"4400", 1690=>x"3800", 1691=>x"3000", 1692=>x"3000", 1693=>x"2b00", 1694=>x"3200",
---- 1695=>x"cd00", 1696=>x"3800", 1697=>x"4b00", 1698=>x"3b00", 1699=>x"3100", 1700=>x"3300", 1701=>x"2e00",
---- 1702=>x"3400", 1703=>x"3200", 1704=>x"3700", 1705=>x"5800", 1706=>x"3800", 1707=>x"2f00", 1708=>x"3100",
---- 1709=>x"2b00", 1710=>x"3200", 1711=>x"3400", 1712=>x"3600", 1713=>x"6000", 1714=>x"3d00", 1715=>x"3200",
---- 1716=>x"3200", 1717=>x"3300", 1718=>x"3200", 1719=>x"2e00", 1720=>x"3600", 1721=>x"5300", 1722=>x"3800",
---- 1723=>x"3600", 1724=>x"3700", 1725=>x"3300", 1726=>x"3300", 1727=>x"3300", 1728=>x"3d00", 1729=>x"4e00",
---- 1730=>x"3600", 1731=>x"3400", 1732=>x"3300", 1733=>x"3100", 1734=>x"2f00", 1735=>x"3300", 1736=>x"3d00",
---- 1737=>x"4200", 1738=>x"3800", 1739=>x"3500", 1740=>x"3800", 1741=>x"3d00", 1742=>x"2f00", 1743=>x"3200",
---- 1744=>x"3800", 1745=>x"3a00", 1746=>x"4300", 1747=>x"3700", 1748=>x"3700", 1749=>x"4000", 1750=>x"3200",
---- 1751=>x"3700", 1752=>x"3b00", 1753=>x"3b00", 1754=>x"3f00", 1755=>x"3500", 1756=>x"3400", 1757=>x"3900",
---- 1758=>x"3200", 1759=>x"3c00", 1760=>x"4400", 1761=>x"3500", 1762=>x"3c00", 1763=>x"3900", 1764=>x"3800",
---- 1765=>x"3a00", 1766=>x"2f00", 1767=>x"3b00", 1768=>x"3700", 1769=>x"3100", 1770=>x"4400", 1771=>x"5200",
---- 1772=>x"3d00", 1773=>x"3500", 1774=>x"3600", 1775=>x"3e00", 1776=>x"6b00", 1777=>x"5c00", 1778=>x"5b00",
---- 1779=>x"4400", 1780=>x"3b00", 1781=>x"3200", 1782=>x"3000", 1783=>x"3700", 1784=>x"9300", 1785=>x"6f00",
---- 1786=>x"6700", 1787=>x"3f00", 1788=>x"3e00", 1789=>x"3400", 1790=>x"3800", 1791=>x"3800", 1792=>x"3f00",
---- 1793=>x"3900", 1794=>x"6200", 1795=>x"7200", 1796=>x"4700", 1797=>x"3400", 1798=>x"3400", 1799=>x"3400",
---- 1800=>x"3700", 1801=>x"3c00", 1802=>x"3200", 1803=>x"4e00", 1804=>x"4900", 1805=>x"3600", 1806=>x"2e00",
---- 1807=>x"2c00", 1808=>x"4000", 1809=>x"3800", 1810=>x"3200", 1811=>x"3100", 1812=>x"3900", 1813=>x"3700",
---- 1814=>x"2f00", 1815=>x"2e00", 1816=>x"4000", 1817=>x"3400", 1818=>x"3300", 1819=>x"3200", 1820=>x"3500",
---- 1821=>x"3400", 1822=>x"2a00", 1823=>x"2e00", 1824=>x"3300", 1825=>x"3100", 1826=>x"3300", 1827=>x"3300",
---- 1828=>x"2e00", 1829=>x"3000", 1830=>x"2e00", 1831=>x"2e00", 1832=>x"3400", 1833=>x"3100", 1834=>x"3300",
---- 1835=>x"2e00", 1836=>x"2c00", 1837=>x"2f00", 1838=>x"2e00", 1839=>x"3100", 1840=>x"2f00", 1841=>x"2d00",
---- 1842=>x"ce00", 1843=>x"2a00", 1844=>x"2900", 1845=>x"3100", 1846=>x"3300", 1847=>x"3300", 1848=>x"3100",
---- 1849=>x"2d00", 1850=>x"2800", 1851=>x"2800", 1852=>x"2b00", 1853=>x"3200", 1854=>x"3c00", 1855=>x"4100",
---- 1856=>x"2f00", 1857=>x"2c00", 1858=>x"2800", 1859=>x"2700", 1860=>x"2f00", 1861=>x"3200", 1862=>x"4500",
---- 1863=>x"4800", 1864=>x"2e00", 1865=>x"2c00", 1866=>x"2800", 1867=>x"2900", 1868=>x"3300", 1869=>x"3600",
---- 1870=>x"4400", 1871=>x"4f00", 1872=>x"2d00", 1873=>x"2a00", 1874=>x"2e00", 1875=>x"2b00", 1876=>x"3500",
---- 1877=>x"3b00", 1878=>x"4a00", 1879=>x"5100", 1880=>x"2800", 1881=>x"2900", 1882=>x"2a00", 1883=>x"2d00",
---- 1884=>x"3800", 1885=>x"4000", 1886=>x"5300", 1887=>x"5a00", 1888=>x"2400", 1889=>x"2a00", 1890=>x"2900",
---- 1891=>x"2c00", 1892=>x"3c00", 1893=>x"4800", 1894=>x"5600", 1895=>x"6100", 1896=>x"2600", 1897=>x"2b00",
---- 1898=>x"2d00", 1899=>x"3800", 1900=>x"4800", 1901=>x"4c00", 1902=>x"5c00", 1903=>x"6800", 1904=>x"2c00",
---- 1905=>x"2a00", 1906=>x"3100", 1907=>x"4800", 1908=>x"4e00", 1909=>x"5400", 1910=>x"6300", 1911=>x"6f00",
---- 1912=>x"2d00", 1913=>x"2b00", 1914=>x"3c00", 1915=>x"4d00", 1916=>x"4b00", 1917=>x"5800", 1918=>x"6b00",
---- 1919=>x"7300", 1920=>x"3000", 1921=>x"3400", 1922=>x"4500", 1923=>x"4f00", 1924=>x"5000", 1925=>x"6200",
---- 1926=>x"6d00", 1927=>x"7800", 1928=>x"3300", 1929=>x"4300", 1930=>x"4b00", 1931=>x"4d00", 1932=>x"5e00",
---- 1933=>x"6600", 1934=>x"6e00", 1935=>x"7900", 1936=>x"3b00", 1937=>x"4a00", 1938=>x"4c00", 1939=>x"5b00",
---- 1940=>x"6700", 1941=>x"6800", 1942=>x"7300", 1943=>x"7500", 1944=>x"4600", 1945=>x"4e00", 1946=>x"5800",
---- 1947=>x"6700", 1948=>x"6900", 1949=>x"6300", 1950=>x"5300", 1951=>x"4000", 1952=>x"4f00", 1953=>x"5600",
---- 1954=>x"5400", 1955=>x"4f00", 1956=>x"4000", 1957=>x"3800", 1958=>x"2500", 1959=>x"2500", 1960=>x"3600",
---- 1961=>x"c400", 1962=>x"2b00", 1963=>x"2500", 1964=>x"2800", 1965=>x"2d00", 1966=>x"3900", 1967=>x"4d00",
---- 1968=>x"2900", 1969=>x"2b00", 1970=>x"3500", 1971=>x"3b00", 1972=>x"4600", 1973=>x"5100", 1974=>x"5900",
---- 1975=>x"6200", 1976=>x"3f00", 1977=>x"4300", 1978=>x"5100", 1979=>x"5500", 1980=>x"5c00", 1981=>x"5a00",
---- 1982=>x"6500", 1983=>x"6a00", 1984=>x"5200", 1985=>x"5600", 1986=>x"5a00", 1987=>x"6200", 1988=>x"6500",
---- 1989=>x"6a00", 1990=>x"7200", 1991=>x"7600", 1992=>x"5900", 1993=>x"5e00", 1994=>x"6a00", 1995=>x"7100",
---- 1996=>x"7000", 1997=>x"7200", 1998=>x"7200", 1999=>x"7500", 2000=>x"6200", 2001=>x"9500", 2002=>x"7000",
---- 2003=>x"7300", 2004=>x"7400", 2005=>x"7200", 2006=>x"7300", 2007=>x"7600", 2008=>x"6900", 2009=>x"6f00",
---- 2010=>x"7100", 2011=>x"7400", 2012=>x"7600", 2013=>x"7400", 2014=>x"7400", 2015=>x"7500", 2016=>x"6a00",
---- 2017=>x"6f00", 2018=>x"6f00", 2019=>x"7000", 2020=>x"7900", 2021=>x"7700", 2022=>x"7700", 2023=>x"7600",
---- 2024=>x"6800", 2025=>x"7100", 2026=>x"7400", 2027=>x"7300", 2028=>x"7800", 2029=>x"7900", 2030=>x"7900",
---- 2031=>x"7800", 2032=>x"7000", 2033=>x"7400", 2034=>x"7600", 2035=>x"7400", 2036=>x"7700", 2037=>x"7a00",
---- 2038=>x"7800", 2039=>x"7a00", 2040=>x"6e00", 2041=>x"6f00", 2042=>x"7400", 2043=>x"7700", 2044=>x"7800",
---- 2045=>x"7b00", 2046=>x"7900", 2047=>x"7c00"),
---- 13 => (0=>x"8700", 1=>x"8600", 2=>x"8700", 3=>x"8200", 4=>x"8100", 5=>x"8200", 6=>x"7b00", 7=>x"8200",
---- 8=>x"8700", 9=>x"8600", 10=>x"8700", 11=>x"7d00", 12=>x"8300", 13=>x"8200", 14=>x"8400",
---- 15=>x"8100", 16=>x"8600", 17=>x"8600", 18=>x"8500", 19=>x"7e00", 20=>x"8100", 21=>x"8200",
---- 22=>x"8600", 23=>x"8300", 24=>x"8600", 25=>x"8500", 26=>x"8700", 27=>x"7e00", 28=>x"8200",
---- 29=>x"8100", 30=>x"8200", 31=>x"8200", 32=>x"8300", 33=>x"8200", 34=>x"8500", 35=>x"8500",
---- 36=>x"8300", 37=>x"8000", 38=>x"7f00", 39=>x"7f00", 40=>x"8100", 41=>x"8500", 42=>x"8200",
---- 43=>x"8100", 44=>x"8200", 45=>x"8200", 46=>x"8000", 47=>x"8000", 48=>x"8600", 49=>x"8500",
---- 50=>x"8400", 51=>x"8400", 52=>x"8200", 53=>x"8100", 54=>x"8200", 55=>x"8200", 56=>x"8200",
---- 57=>x"8300", 58=>x"8300", 59=>x"8300", 60=>x"8200", 61=>x"8100", 62=>x"8500", 63=>x"8200",
---- 64=>x"8600", 65=>x"8500", 66=>x"8600", 67=>x"8200", 68=>x"8600", 69=>x"8500", 70=>x"8400",
---- 71=>x"7f00", 72=>x"8300", 73=>x"8300", 74=>x"8500", 75=>x"8400", 76=>x"8900", 77=>x"8200",
---- 78=>x"8200", 79=>x"8100", 80=>x"8700", 81=>x"8200", 82=>x"8100", 83=>x"8200", 84=>x"8300",
---- 85=>x"8200", 86=>x"8700", 87=>x"8300", 88=>x"8500", 89=>x"7e00", 90=>x"8100", 91=>x"8100",
---- 92=>x"8000", 93=>x"8200", 94=>x"8100", 95=>x"8000", 96=>x"7e00", 97=>x"7f00", 98=>x"8000",
---- 99=>x"7e00", 100=>x"7f00", 101=>x"7f00", 102=>x"7e00", 103=>x"8100", 104=>x"7e00", 105=>x"7d00",
---- 106=>x"7c00", 107=>x"7e00", 108=>x"7f00", 109=>x"8000", 110=>x"7e00", 111=>x"8000", 112=>x"7c00",
---- 113=>x"7900", 114=>x"7b00", 115=>x"7b00", 116=>x"7c00", 117=>x"7e00", 118=>x"8200", 119=>x"8100",
---- 120=>x"7b00", 121=>x"7900", 122=>x"7b00", 123=>x"8500", 124=>x"7c00", 125=>x"7c00", 126=>x"7e00",
---- 127=>x"8000", 128=>x"7b00", 129=>x"7a00", 130=>x"7c00", 131=>x"7900", 132=>x"7c00", 133=>x"7900",
---- 134=>x"7900", 135=>x"8000", 136=>x"7b00", 137=>x"7d00", 138=>x"7900", 139=>x"7600", 140=>x"7a00",
---- 141=>x"7900", 142=>x"7c00", 143=>x"7d00", 144=>x"7c00", 145=>x"7d00", 146=>x"7c00", 147=>x"7900",
---- 148=>x"7d00", 149=>x"7b00", 150=>x"7d00", 151=>x"7e00", 152=>x"7c00", 153=>x"7b00", 154=>x"7800",
---- 155=>x"7a00", 156=>x"7d00", 157=>x"7900", 158=>x"7a00", 159=>x"7d00", 160=>x"8100", 161=>x"7b00",
---- 162=>x"7a00", 163=>x"7c00", 164=>x"7d00", 165=>x"7b00", 166=>x"7600", 167=>x"7700", 168=>x"7e00",
---- 169=>x"7d00", 170=>x"7f00", 171=>x"7d00", 172=>x"7b00", 173=>x"7a00", 174=>x"7a00", 175=>x"7400",
---- 176=>x"7f00", 177=>x"7c00", 178=>x"7a00", 179=>x"7b00", 180=>x"7900", 181=>x"7b00", 182=>x"7e00",
---- 183=>x"8b00", 184=>x"8700", 185=>x"8a00", 186=>x"8800", 187=>x"8700", 188=>x"8500", 189=>x"9000",
---- 190=>x"9e00", 191=>x"ac00", 192=>x"9700", 193=>x"9100", 194=>x"9100", 195=>x"6900", 196=>x"a000",
---- 197=>x"a400", 198=>x"5500", 199=>x"aa00", 200=>x"9300", 201=>x"9100", 202=>x"9a00", 203=>x"a800",
---- 204=>x"5500", 205=>x"a300", 206=>x"a700", 207=>x"ab00", 208=>x"9200", 209=>x"9900", 210=>x"a400",
---- 211=>x"ac00", 212=>x"aa00", 213=>x"a700", 214=>x"a800", 215=>x"ac00", 216=>x"9600", 217=>x"9800",
---- 218=>x"9d00", 219=>x"a800", 220=>x"a000", 221=>x"a300", 222=>x"aa00", 223=>x"ab00", 224=>x"9600",
---- 225=>x"9300", 226=>x"9800", 227=>x"9900", 228=>x"a000", 229=>x"9f00", 230=>x"a000", 231=>x"a500",
---- 232=>x"9500", 233=>x"9300", 234=>x"9700", 235=>x"9c00", 236=>x"9c00", 237=>x"9f00", 238=>x"a600",
---- 239=>x"a500", 240=>x"9700", 241=>x"9500", 242=>x"9900", 243=>x"9900", 244=>x"9800", 245=>x"a100",
---- 246=>x"aa00", 247=>x"a500", 248=>x"9500", 249=>x"9b00", 250=>x"9800", 251=>x"9600", 252=>x"9c00",
---- 253=>x"a800", 254=>x"a000", 255=>x"a000", 256=>x"9300", 257=>x"9500", 258=>x"9000", 259=>x"9900",
---- 260=>x"9e00", 261=>x"a000", 262=>x"9e00", 263=>x"9800", 264=>x"8c00", 265=>x"9000", 266=>x"8f00",
---- 267=>x"9400", 268=>x"9900", 269=>x"9800", 270=>x"9800", 271=>x"9b00", 272=>x"8c00", 273=>x"8c00",
---- 274=>x"9200", 275=>x"8e00", 276=>x"9200", 277=>x"9a00", 278=>x"9c00", 279=>x"a200", 280=>x"8900",
---- 281=>x"8600", 282=>x"8200", 283=>x"8f00", 284=>x"9100", 285=>x"9900", 286=>x"9d00", 287=>x"a200",
---- 288=>x"8d00", 289=>x"8d00", 290=>x"8c00", 291=>x"9100", 292=>x"9300", 293=>x"9000", 294=>x"9900",
---- 295=>x"a000", 296=>x"8600", 297=>x"8e00", 298=>x"8a00", 299=>x"8e00", 300=>x"8c00", 301=>x"9700",
---- 302=>x"9500", 303=>x"9900", 304=>x"8500", 305=>x"8800", 306=>x"8500", 307=>x"8900", 308=>x"9800",
---- 309=>x"6800", 310=>x"9300", 311=>x"9700", 312=>x"7400", 313=>x"8f00", 314=>x"8400", 315=>x"8f00",
---- 316=>x"9400", 317=>x"9100", 318=>x"9200", 319=>x"9600", 320=>x"8100", 321=>x"7900", 322=>x"8700",
---- 323=>x"9500", 324=>x"8d00", 325=>x"9000", 326=>x"9700", 327=>x"9800", 328=>x"8700", 329=>x"8200",
---- 330=>x"8d00", 331=>x"8f00", 332=>x"8800", 333=>x"8800", 334=>x"9300", 335=>x"9800", 336=>x"8200",
---- 337=>x"8a00", 338=>x"8600", 339=>x"8c00", 340=>x"8600", 341=>x"8b00", 342=>x"9300", 343=>x"8c00",
---- 344=>x"8800", 345=>x"8400", 346=>x"8f00", 347=>x"8c00", 348=>x"8c00", 349=>x"8d00", 350=>x"9000",
---- 351=>x"9f00", 352=>x"8500", 353=>x"9100", 354=>x"8b00", 355=>x"8d00", 356=>x"8e00", 357=>x"8d00",
---- 358=>x"9500", 359=>x"9400", 360=>x"8d00", 361=>x"8f00", 362=>x"8d00", 363=>x"8e00", 364=>x"9300",
---- 365=>x"9800", 366=>x"9100", 367=>x"9100", 368=>x"8b00", 369=>x"9300", 370=>x"9300", 371=>x"9100",
---- 372=>x"8f00", 373=>x"8d00", 374=>x"9000", 375=>x"9000", 376=>x"9400", 377=>x"9300", 378=>x"8f00",
---- 379=>x"8100", 380=>x"8e00", 381=>x"8900", 382=>x"8d00", 383=>x"9400", 384=>x"9500", 385=>x"9000",
---- 386=>x"8600", 387=>x"8a00", 388=>x"9000", 389=>x"8800", 390=>x"9100", 391=>x"6e00", 392=>x"9200",
---- 393=>x"8700", 394=>x"8e00", 395=>x"8b00", 396=>x"8c00", 397=>x"8e00", 398=>x"9100", 399=>x"9200",
---- 400=>x"8800", 401=>x"8c00", 402=>x"8400", 403=>x"8400", 404=>x"8800", 405=>x"8800", 406=>x"8f00",
---- 407=>x"8d00", 408=>x"8700", 409=>x"8500", 410=>x"8700", 411=>x"8100", 412=>x"8900", 413=>x"8d00",
---- 414=>x"8b00", 415=>x"9100", 416=>x"8500", 417=>x"8a00", 418=>x"8900", 419=>x"8500", 420=>x"8700",
---- 421=>x"8d00", 422=>x"8d00", 423=>x"8200", 424=>x"8400", 425=>x"8500", 426=>x"8200", 427=>x"7d00",
---- 428=>x"8500", 429=>x"8200", 430=>x"7e00", 431=>x"7a00", 432=>x"8500", 433=>x"8200", 434=>x"7800",
---- 435=>x"8200", 436=>x"8200", 437=>x"7600", 438=>x"7e00", 439=>x"9c00", 440=>x"8300", 441=>x"8000",
---- 442=>x"7900", 443=>x"6f00", 444=>x"6d00", 445=>x"8100", 446=>x"a400", 447=>x"ad00", 448=>x"7e00",
---- 449=>x"7b00", 450=>x"6900", 451=>x"6e00", 452=>x"9000", 453=>x"b100", 454=>x"b800", 455=>x"b000",
---- 456=>x"7900", 457=>x"6a00", 458=>x"7500", 459=>x"9700", 460=>x"a700", 461=>x"b600", 462=>x"ba00",
---- 463=>x"c100", 464=>x"6e00", 465=>x"7f00", 466=>x"a600", 467=>x"b300", 468=>x"a500", 469=>x"b300",
---- 470=>x"c700", 471=>x"c000", 472=>x"9000", 473=>x"a500", 474=>x"a500", 475=>x"b400", 476=>x"b900",
---- 477=>x"b200", 478=>x"c300", 479=>x"b300", 480=>x"ad00", 481=>x"ab00", 482=>x"ae00", 483=>x"bd00",
---- 484=>x"b400", 485=>x"a600", 486=>x"b100", 487=>x"b400", 488=>x"af00", 489=>x"b700", 490=>x"b500",
---- 491=>x"b400", 492=>x"a800", 493=>x"a000", 494=>x"a100", 495=>x"a900", 496=>x"b500", 497=>x"b800",
---- 498=>x"a900", 499=>x"a900", 500=>x"a700", 501=>x"a300", 502=>x"a300", 503=>x"b300", 504=>x"af00",
---- 505=>x"a800", 506=>x"a400", 507=>x"a200", 508=>x"a400", 509=>x"b000", 510=>x"b100", 511=>x"a700",
---- 512=>x"a900", 513=>x"a100", 514=>x"9800", 515=>x"a700", 516=>x"4900", 517=>x"ab00", 518=>x"a200",
---- 519=>x"ad00", 520=>x"9e00", 521=>x"a600", 522=>x"ac00", 523=>x"a700", 524=>x"a300", 525=>x"a000",
---- 526=>x"b500", 527=>x"b700", 528=>x"a300", 529=>x"b300", 530=>x"aa00", 531=>x"9500", 532=>x"a100",
---- 533=>x"5000", 534=>x"af00", 535=>x"b900", 536=>x"ae00", 537=>x"9e00", 538=>x"9500", 539=>x"ac00",
---- 540=>x"b300", 541=>x"ac00", 542=>x"aa00", 543=>x"ab00", 544=>x"8600", 545=>x"9500", 546=>x"ad00",
---- 547=>x"b100", 548=>x"af00", 549=>x"ab00", 550=>x"b000", 551=>x"b200", 552=>x"9600", 553=>x"9f00",
---- 554=>x"a900", 555=>x"ae00", 556=>x"aa00", 557=>x"b200", 558=>x"b300", 559=>x"b300", 560=>x"a700",
---- 561=>x"a700", 562=>x"9800", 563=>x"a400", 564=>x"b400", 565=>x"b300", 566=>x"4c00", 567=>x"a600",
---- 568=>x"a000", 569=>x"a200", 570=>x"a400", 571=>x"a700", 572=>x"ae00", 573=>x"b000", 574=>x"aa00",
---- 575=>x"a900", 576=>x"9800", 577=>x"a300", 578=>x"ae00", 579=>x"a200", 580=>x"9500", 581=>x"a400",
---- 582=>x"a900", 583=>x"a700", 584=>x"a600", 585=>x"a300", 586=>x"a100", 587=>x"a000", 588=>x"a000",
---- 589=>x"9c00", 590=>x"a100", 591=>x"ae00", 592=>x"ae00", 593=>x"9900", 594=>x"9400", 595=>x"9e00",
---- 596=>x"9f00", 597=>x"a500", 598=>x"aa00", 599=>x"aa00", 600=>x"8800", 601=>x"9d00", 602=>x"9400",
---- 603=>x"9a00", 604=>x"ac00", 605=>x"ad00", 606=>x"af00", 607=>x"ad00", 608=>x"8900", 609=>x"8d00",
---- 610=>x"9a00", 611=>x"a100", 612=>x"a500", 613=>x"b700", 614=>x"ae00", 615=>x"a900", 616=>x"8e00",
---- 617=>x"9300", 618=>x"9400", 619=>x"a200", 620=>x"9f00", 621=>x"9e00", 622=>x"b100", 623=>x"a200",
---- 624=>x"9d00", 625=>x"a200", 626=>x"9200", 627=>x"8800", 628=>x"a300", 629=>x"9c00", 630=>x"9600",
---- 631=>x"9400", 632=>x"9600", 633=>x"9100", 634=>x"9100", 635=>x"8e00", 636=>x"9800", 637=>x"9f00",
---- 638=>x"8900", 639=>x"9800", 640=>x"8a00", 641=>x"9900", 642=>x"9d00", 643=>x"9b00", 644=>x"8b00",
---- 645=>x"8e00", 646=>x"a700", 647=>x"9d00", 648=>x"9e00", 649=>x"9d00", 650=>x"a000", 651=>x"9100",
---- 652=>x"8b00", 653=>x"9300", 654=>x"a400", 655=>x"a800", 656=>x"9900", 657=>x"9500", 658=>x"8a00",
---- 659=>x"8e00", 660=>x"5f00", 661=>x"a300", 662=>x"9900", 663=>x"9c00", 664=>x"9100", 665=>x"8600",
---- 666=>x"8900", 667=>x"9900", 668=>x"9e00", 669=>x"9f00", 670=>x"a000", 671=>x"6500", 672=>x"8700",
---- 673=>x"7200", 674=>x"9e00", 675=>x"a000", 676=>x"9a00", 677=>x"9b00", 678=>x"9e00", 679=>x"9d00",
---- 680=>x"8200", 681=>x"9400", 682=>x"9c00", 683=>x"a400", 684=>x"a200", 685=>x"9c00", 686=>x"9700",
---- 687=>x"8800", 688=>x"9500", 689=>x"9100", 690=>x"9700", 691=>x"9a00", 692=>x"9300", 693=>x"7400",
---- 694=>x"6900", 695=>x"6b00", 696=>x"9d00", 697=>x"9a00", 698=>x"9300", 699=>x"8400", 700=>x"6100",
---- 701=>x"6200", 702=>x"8800", 703=>x"8c00", 704=>x"9200", 705=>x"9900", 706=>x"9200", 707=>x"6c00",
---- 708=>x"7300", 709=>x"8b00", 710=>x"9100", 711=>x"8900", 712=>x"9800", 713=>x"8d00", 714=>x"7400",
---- 715=>x"8300", 716=>x"9800", 717=>x"8e00", 718=>x"8700", 719=>x"6b00", 720=>x"8b00", 721=>x"7300",
---- 722=>x"8e00", 723=>x"8b00", 724=>x"9400", 725=>x"8300", 726=>x"6600", 727=>x"5f00", 728=>x"6d00",
---- 729=>x"6800", 730=>x"8b00", 731=>x"8f00", 732=>x"8500", 733=>x"7200", 734=>x"6800", 735=>x"8000",
---- 736=>x"6d00", 737=>x"8400", 738=>x"8300", 739=>x"8300", 740=>x"7400", 741=>x"6700", 742=>x"8000",
---- 743=>x"7f00", 744=>x"8400", 745=>x"8700", 746=>x"8500", 747=>x"7a00", 748=>x"6700", 749=>x"7c00",
---- 750=>x"8400", 751=>x"7400", 752=>x"8300", 753=>x"8900", 754=>x"8500", 755=>x"7800", 756=>x"6700",
---- 757=>x"7000", 758=>x"5700", 759=>x"4c00", 760=>x"8500", 761=>x"8200", 762=>x"7500", 763=>x"6100",
---- 764=>x"5000", 765=>x"4300", 766=>x"3e00", 767=>x"5200", 768=>x"7e00", 769=>x"6600", 770=>x"5000",
---- 771=>x"4000", 772=>x"3100", 773=>x"4f00", 774=>x"6b00", 775=>x"5800", 776=>x"5700", 777=>x"4700",
---- 778=>x"3800", 779=>x"3a00", 780=>x"5d00", 781=>x"6300", 782=>x"4300", 783=>x"2f00", 784=>x"4000",
---- 785=>x"3c00", 786=>x"4200", 787=>x"5f00", 788=>x"5200", 789=>x"3500", 790=>x"2f00", 791=>x"2b00",
---- 792=>x"4200", 793=>x"4f00", 794=>x"5300", 795=>x"4900", 796=>x"3800", 797=>x"3d00", 798=>x"3500",
---- 799=>x"3000", 800=>x"4500", 801=>x"5800", 802=>x"4f00", 803=>x"4600", 804=>x"3e00", 805=>x"3500",
---- 806=>x"3300", 807=>x"5a00", 808=>x"5600", 809=>x"5700", 810=>x"4200", 811=>x"3f00", 812=>x"3000",
---- 813=>x"2500", 814=>x"5300", 815=>x"6d00", 816=>x"4900", 817=>x"3600", 818=>x"3100", 819=>x"2d00",
---- 820=>x"2b00", 821=>x"3e00", 822=>x"7400", 823=>x"6500", 824=>x"3e00", 825=>x"2e00", 826=>x"2700",
---- 827=>x"2500", 828=>x"2e00", 829=>x"4a00", 830=>x"7a00", 831=>x"5500", 832=>x"3700", 833=>x"3300",
---- 834=>x"2f00", 835=>x"2900", 836=>x"2b00", 837=>x"5500", 838=>x"7800", 839=>x"4100", 840=>x"3b00",
---- 841=>x"3a00", 842=>x"3600", 843=>x"2a00", 844=>x"3600", 845=>x"5100", 846=>x"5e00", 847=>x"4600",
---- 848=>x"3d00", 849=>x"3100", 850=>x"2f00", 851=>x"3100", 852=>x"4100", 853=>x"4400", 854=>x"b400",
---- 855=>x"5800", 856=>x"4900", 857=>x"4200", 858=>x"3800", 859=>x"3300", 860=>x"4b00", 861=>x"3b00",
---- 862=>x"3c00", 863=>x"6e00", 864=>x"4d00", 865=>x"5800", 866=>x"4000", 867=>x"2b00", 868=>x"4a00",
---- 869=>x"3800", 870=>x"3300", 871=>x"6600", 872=>x"4900", 873=>x"5d00", 874=>x"4300", 875=>x"2800",
---- 876=>x"4a00", 877=>x"4200", 878=>x"2300", 879=>x"4c00", 880=>x"3e00", 881=>x"5200", 882=>x"4f00",
---- 883=>x"2a00", 884=>x"4300", 885=>x"4e00", 886=>x"2100", 887=>x"3200", 888=>x"4400", 889=>x"4200",
---- 890=>x"4d00", 891=>x"3900", 892=>x"4600", 893=>x"5200", 894=>x"2800", 895=>x"3800", 896=>x"4d00",
---- 897=>x"4200", 898=>x"3d00", 899=>x"3e00", 900=>x"5100", 901=>x"4600", 902=>x"3300", 903=>x"3f00",
---- 904=>x"3600", 905=>x"4100", 906=>x"3900", 907=>x"3400", 908=>x"5800", 909=>x"5800", 910=>x"5100",
---- 911=>x"4600", 912=>x"2d00", 913=>x"4000", 914=>x"3800", 915=>x"3100", 916=>x"4200", 917=>x"6a00",
---- 918=>x"7900", 919=>x"5800", 920=>x"3500", 921=>x"3f00", 922=>x"2c00", 923=>x"3a00", 924=>x"4f00",
---- 925=>x"5900", 926=>x"5900", 927=>x"6200", 928=>x"4600", 929=>x"3e00", 930=>x"2800", 931=>x"2a00",
---- 932=>x"6000", 933=>x"5100", 934=>x"4900", 935=>x"4b00", 936=>x"4a00", 937=>x"3700", 938=>x"3100",
---- 939=>x"2d00", 940=>x"4c00", 941=>x"3700", 942=>x"4a00", 943=>x"3f00", 944=>x"4300", 945=>x"4000",
---- 946=>x"3d00", 947=>x"2d00", 948=>x"2a00", 949=>x"3600", 950=>x"5000", 951=>x"4600", 952=>x"3b00",
---- 953=>x"3100", 954=>x"4700", 955=>x"3500", 956=>x"3200", 957=>x"2c00", 958=>x"6500", 959=>x"5e00",
---- 960=>x"3100", 961=>x"2b00", 962=>x"5a00", 963=>x"4900", 964=>x"3100", 965=>x"3a00", 966=>x"6300",
---- 967=>x"2f00", 968=>x"2600", 969=>x"2800", 970=>x"6100", 971=>x"4a00", 972=>x"1f00", 973=>x"5700",
---- 974=>x"3a00", 975=>x"2d00", 976=>x"1f00", 977=>x"3100", 978=>x"6700", 979=>x"3e00", 980=>x"2d00",
---- 981=>x"5b00", 982=>x"3c00", 983=>x"c700", 984=>x"2a00", 985=>x"3d00", 986=>x"5b00", 987=>x"4300",
---- 988=>x"3a00", 989=>x"4900", 990=>x"2600", 991=>x"1d00", 992=>x"3a00", 993=>x"4000", 994=>x"4a00",
---- 995=>x"4600", 996=>x"3600", 997=>x"3900", 998=>x"1f00", 999=>x"2900", 1000=>x"5200", 1001=>x"5a00",
---- 1002=>x"3900", 1003=>x"4b00", 1004=>x"3b00", 1005=>x"2b00", 1006=>x"1f00", 1007=>x"5600", 1008=>x"5300",
---- 1009=>x"7300", 1010=>x"3300", 1011=>x"4300", 1012=>x"3500", 1013=>x"1800", 1014=>x"3200", 1015=>x"8f00",
---- 1016=>x"2a00", 1017=>x"4000", 1018=>x"5200", 1019=>x"2a00", 1020=>x"1e00", 1021=>x"2200", 1022=>x"7200",
---- 1023=>x"9100", 1024=>x"2b00", 1025=>x"2400", 1026=>x"3000", 1027=>x"3900", 1028=>x"1800", 1029=>x"4900",
---- 1030=>x"9d00", 1031=>x"6e00", 1032=>x"2b00", 1033=>x"2600", 1034=>x"2500", 1035=>x"2300", 1036=>x"2b00",
---- 1037=>x"8900", 1038=>x"8c00", 1039=>x"6a00", 1040=>x"2e00", 1041=>x"2500", 1042=>x"2800", 1043=>x"1800",
---- 1044=>x"5e00", 1045=>x"9f00", 1046=>x"6a00", 1047=>x"9d00", 1048=>x"2900", 1049=>x"2500", 1050=>x"1e00",
---- 1051=>x"3800", 1052=>x"9600", 1053=>x"7800", 1054=>x"7900", 1055=>x"c400", 1056=>x"2600", 1057=>x"2000",
---- 1058=>x"1d00", 1059=>x"7100", 1060=>x"9500", 1061=>x"6000", 1062=>x"ac00", 1063=>x"b900", 1064=>x"3200",
---- 1065=>x"3d00", 1066=>x"4700", 1067=>x"9600", 1068=>x"6b00", 1069=>x"8c00", 1070=>x"c800", 1071=>x"a900",
---- 1072=>x"2500", 1073=>x"3400", 1074=>x"7000", 1075=>x"7300", 1076=>x"6700", 1077=>x"b400", 1078=>x"ac00",
---- 1079=>x"9700", 1080=>x"2400", 1081=>x"4c00", 1082=>x"7e00", 1083=>x"5100", 1084=>x"8e00", 1085=>x"a500",
---- 1086=>x"9700", 1087=>x"a500", 1088=>x"3f00", 1089=>x"8900", 1090=>x"6c00", 1091=>x"6d00", 1092=>x"bb00",
---- 1093=>x"9c00", 1094=>x"a900", 1095=>x"b600", 1096=>x"6d00", 1097=>x"8b00", 1098=>x"5e00", 1099=>x"af00",
---- 1100=>x"be00", 1101=>x"9d00", 1102=>x"af00", 1103=>x"b800", 1104=>x"9500", 1105=>x"6300", 1106=>x"8100",
---- 1107=>x"c800", 1108=>x"a900", 1109=>x"ab00", 1110=>x"b700", 1111=>x"be00", 1112=>x"8400", 1113=>x"5e00",
---- 1114=>x"5200", 1115=>x"b100", 1116=>x"a400", 1117=>x"b300", 1118=>x"ba00", 1119=>x"c500", 1120=>x"6500",
---- 1121=>x"7c00", 1122=>x"b300", 1123=>x"a300", 1124=>x"af00", 1125=>x"b200", 1126=>x"be00", 1127=>x"c800",
---- 1128=>x"6600", 1129=>x"a800", 1130=>x"ad00", 1131=>x"a600", 1132=>x"b500", 1133=>x"b900", 1134=>x"c600",
---- 1135=>x"d200", 1136=>x"7f00", 1137=>x"4800", 1138=>x"af00", 1139=>x"b300", 1140=>x"bb00", 1141=>x"c400",
---- 1142=>x"d200", 1143=>x"b000", 1144=>x"9c00", 1145=>x"b000", 1146=>x"b700", 1147=>x"bd00", 1148=>x"c200",
---- 1149=>x"d200", 1150=>x"be00", 1151=>x"5000", 1152=>x"b400", 1153=>x"ae00", 1154=>x"be00", 1155=>x"4000",
---- 1156=>x"c600", 1157=>x"ca00", 1158=>x"6000", 1159=>x"3900", 1160=>x"b400", 1161=>x"b800", 1162=>x"bd00",
---- 1163=>x"c400", 1164=>x"d100", 1165=>x"7900", 1166=>x"2d00", 1167=>x"4800", 1168=>x"b400", 1169=>x"c000",
---- 1170=>x"c300", 1171=>x"d600", 1172=>x"9800", 1173=>x"2700", 1174=>x"3400", 1175=>x"4c00", 1176=>x"bc00",
---- 1177=>x"c000", 1178=>x"cf00", 1179=>x"bd00", 1180=>x"3800", 1181=>x"2300", 1182=>x"3900", 1183=>x"5200",
---- 1184=>x"bc00", 1185=>x"3e00", 1186=>x"cf00", 1187=>x"5700", 1188=>x"2000", 1189=>x"3400", 1190=>x"3b00",
---- 1191=>x"5400", 1192=>x"bb00", 1193=>x"d000", 1194=>x"8600", 1195=>x"2000", 1196=>x"2c00", 1197=>x"3100",
---- 1198=>x"4200", 1199=>x"5800", 1200=>x"cc00", 1201=>x"4d00", 1202=>x"3600", 1203=>x"2a00", 1204=>x"3600",
---- 1205=>x"3200", 1206=>x"3f00", 1207=>x"5800", 1208=>x"d200", 1209=>x"5b00", 1210=>x"1d00", 1211=>x"2d00",
---- 1212=>x"3900", 1213=>x"3200", 1214=>x"3f00", 1215=>x"5400", 1216=>x"9500", 1217=>x"2000", 1218=>x"2500",
---- 1219=>x"2e00", 1220=>x"4200", 1221=>x"3400", 1222=>x"4300", 1223=>x"5500", 1224=>x"3f00", 1225=>x"1e00",
---- 1226=>x"2500", 1227=>x"2f00", 1228=>x"4a00", 1229=>x"3400", 1230=>x"3d00", 1231=>x"5400", 1232=>x"1b00",
---- 1233=>x"2600", 1234=>x"2100", 1235=>x"3000", 1236=>x"4f00", 1237=>x"3800", 1238=>x"3d00", 1239=>x"5100",
---- 1240=>x"2600", 1241=>x"2400", 1242=>x"2300", 1243=>x"3000", 1244=>x"5600", 1245=>x"3b00", 1246=>x"4300",
---- 1247=>x"4e00", 1248=>x"2900", 1249=>x"2800", 1250=>x"2200", 1251=>x"3100", 1252=>x"5f00", 1253=>x"4500",
---- 1254=>x"4400", 1255=>x"5100", 1256=>x"2700", 1257=>x"2600", 1258=>x"2300", 1259=>x"3500", 1260=>x"6700",
---- 1261=>x"4400", 1262=>x"4200", 1263=>x"5200", 1264=>x"2700", 1265=>x"2800", 1266=>x"2700", 1267=>x"3500",
---- 1268=>x"6900", 1269=>x"4800", 1270=>x"4500", 1271=>x"5000", 1272=>x"2b00", 1273=>x"2800", 1274=>x"2900",
---- 1275=>x"3600", 1276=>x"6b00", 1277=>x"5600", 1278=>x"4200", 1279=>x"4e00", 1280=>x"2d00", 1281=>x"2d00",
---- 1282=>x"2400", 1283=>x"3900", 1284=>x"6900", 1285=>x"5500", 1286=>x"4000", 1287=>x"5000", 1288=>x"3000",
---- 1289=>x"2900", 1290=>x"2500", 1291=>x"3800", 1292=>x"6a00", 1293=>x"5700", 1294=>x"4b00", 1295=>x"5700",
---- 1296=>x"3200", 1297=>x"3000", 1298=>x"2700", 1299=>x"3400", 1300=>x"6c00", 1301=>x"6000", 1302=>x"4b00",
---- 1303=>x"5d00", 1304=>x"2d00", 1305=>x"2e00", 1306=>x"2a00", 1307=>x"3900", 1308=>x"7100", 1309=>x"6300",
---- 1310=>x"4a00", 1311=>x"5e00", 1312=>x"2b00", 1313=>x"2b00", 1314=>x"3000", 1315=>x"3a00", 1316=>x"7400",
---- 1317=>x"6a00", 1318=>x"5000", 1319=>x"5900", 1320=>x"3000", 1321=>x"2a00", 1322=>x"2500", 1323=>x"3b00",
---- 1324=>x"7900", 1325=>x"6700", 1326=>x"5200", 1327=>x"5a00", 1328=>x"3500", 1329=>x"3000", 1330=>x"2a00",
---- 1331=>x"3c00", 1332=>x"7500", 1333=>x"6900", 1334=>x"5400", 1335=>x"5b00", 1336=>x"3300", 1337=>x"3000",
---- 1338=>x"2c00", 1339=>x"3d00", 1340=>x"6e00", 1341=>x"6b00", 1342=>x"5d00", 1343=>x"5f00", 1344=>x"3800",
---- 1345=>x"3100", 1346=>x"2e00", 1347=>x"3500", 1348=>x"6a00", 1349=>x"6f00", 1350=>x"5f00", 1351=>x"5e00",
---- 1352=>x"3300", 1353=>x"3100", 1354=>x"2800", 1355=>x"3000", 1356=>x"6700", 1357=>x"6900", 1358=>x"6500",
---- 1359=>x"5b00", 1360=>x"3300", 1361=>x"3200", 1362=>x"2900", 1363=>x"2d00", 1364=>x"5e00", 1365=>x"6500",
---- 1366=>x"6a00", 1367=>x"5700", 1368=>x"3b00", 1369=>x"3000", 1370=>x"2a00", 1371=>x"2b00", 1372=>x"5e00",
---- 1373=>x"6400", 1374=>x"6900", 1375=>x"5600", 1376=>x"4400", 1377=>x"2d00", 1378=>x"2a00", 1379=>x"2a00",
---- 1380=>x"5700", 1381=>x"6000", 1382=>x"6600", 1383=>x"5900", 1384=>x"4200", 1385=>x"2e00", 1386=>x"2c00",
---- 1387=>x"2b00", 1388=>x"5800", 1389=>x"5b00", 1390=>x"6200", 1391=>x"5700", 1392=>x"4900", 1393=>x"2f00",
---- 1394=>x"2c00", 1395=>x"2c00", 1396=>x"5c00", 1397=>x"5c00", 1398=>x"5c00", 1399=>x"5300", 1400=>x"5100",
---- 1401=>x"3300", 1402=>x"2600", 1403=>x"2900", 1404=>x"5600", 1405=>x"5200", 1406=>x"5700", 1407=>x"5a00",
---- 1408=>x"5100", 1409=>x"3a00", 1410=>x"2900", 1411=>x"2a00", 1412=>x"5200", 1413=>x"5200", 1414=>x"5500",
---- 1415=>x"5800", 1416=>x"4b00", 1417=>x"4000", 1418=>x"2c00", 1419=>x"2b00", 1420=>x"5200", 1421=>x"4e00",
---- 1422=>x"4f00", 1423=>x"5300", 1424=>x"4500", 1425=>x"4200", 1426=>x"2d00", 1427=>x"3000", 1428=>x"5000",
---- 1429=>x"4a00", 1430=>x"4b00", 1431=>x"5400", 1432=>x"4500", 1433=>x"4700", 1434=>x"3100", 1435=>x"2c00",
---- 1436=>x"bb00", 1437=>x"4500", 1438=>x"4b00", 1439=>x"5400", 1440=>x"4300", 1441=>x"4500", 1442=>x"3300",
---- 1443=>x"2e00", 1444=>x"4700", 1445=>x"4d00", 1446=>x"4c00", 1447=>x"5100", 1448=>x"b900", 1449=>x"4600",
---- 1450=>x"3900", 1451=>x"3100", 1452=>x"4400", 1453=>x"4f00", 1454=>x"4900", 1455=>x"4e00", 1456=>x"3e00",
---- 1457=>x"4700", 1458=>x"3d00", 1459=>x"3200", 1460=>x"3b00", 1461=>x"4c00", 1462=>x"4600", 1463=>x"5500",
---- 1464=>x"3b00", 1465=>x"3e00", 1466=>x"3a00", 1467=>x"3300", 1468=>x"3600", 1469=>x"4900", 1470=>x"4100",
---- 1471=>x"5200", 1472=>x"3b00", 1473=>x"3c00", 1474=>x"4200", 1475=>x"3900", 1476=>x"3100", 1477=>x"3f00",
---- 1478=>x"3b00", 1479=>x"4b00", 1480=>x"3900", 1481=>x"3d00", 1482=>x"4000", 1483=>x"3800", 1484=>x"2c00",
---- 1485=>x"3a00", 1486=>x"3d00", 1487=>x"3e00", 1488=>x"3700", 1489=>x"3d00", 1490=>x"4300", 1491=>x"3600",
---- 1492=>x"2f00", 1493=>x"3500", 1494=>x"4000", 1495=>x"3a00", 1496=>x"3700", 1497=>x"3800", 1498=>x"3e00",
---- 1499=>x"3800", 1500=>x"3200", 1501=>x"3200", 1502=>x"3e00", 1503=>x"3b00", 1504=>x"3700", 1505=>x"3900",
---- 1506=>x"3700", 1507=>x"3b00", 1508=>x"3600", 1509=>x"3500", 1510=>x"3b00", 1511=>x"3900", 1512=>x"3800",
---- 1513=>x"3a00", 1514=>x"3900", 1515=>x"3400", 1516=>x"3800", 1517=>x"3900", 1518=>x"3b00", 1519=>x"3a00",
---- 1520=>x"3200", 1521=>x"3800", 1522=>x"3c00", 1523=>x"3400", 1524=>x"3b00", 1525=>x"3300", 1526=>x"3900",
---- 1527=>x"3d00", 1528=>x"3200", 1529=>x"3400", 1530=>x"3d00", 1531=>x"3800", 1532=>x"3c00", 1533=>x"3d00",
---- 1534=>x"3400", 1535=>x"3a00", 1536=>x"2f00", 1537=>x"3000", 1538=>x"3500", 1539=>x"3700", 1540=>x"3e00",
---- 1541=>x"3d00", 1542=>x"3700", 1543=>x"3b00", 1544=>x"2f00", 1545=>x"3000", 1546=>x"3400", 1547=>x"3400",
---- 1548=>x"3a00", 1549=>x"3f00", 1550=>x"3d00", 1551=>x"3f00", 1552=>x"3400", 1553=>x"2e00", 1554=>x"3500",
---- 1555=>x"3200", 1556=>x"3800", 1557=>x"3d00", 1558=>x"3e00", 1559=>x"3800", 1560=>x"3100", 1561=>x"2f00",
---- 1562=>x"3200", 1563=>x"3200", 1564=>x"3400", 1565=>x"3b00", 1566=>x"3b00", 1567=>x"3600", 1568=>x"3100",
---- 1569=>x"2f00", 1570=>x"3100", 1571=>x"3200", 1572=>x"3600", 1573=>x"3900", 1574=>x"3d00", 1575=>x"3900",
---- 1576=>x"3100", 1577=>x"3300", 1578=>x"3400", 1579=>x"3900", 1580=>x"3300", 1581=>x"3400", 1582=>x"3d00",
---- 1583=>x"3f00", 1584=>x"3000", 1585=>x"3400", 1586=>x"3400", 1587=>x"3200", 1588=>x"3600", 1589=>x"2f00",
---- 1590=>x"3a00", 1591=>x"3c00", 1592=>x"3200", 1593=>x"3000", 1594=>x"3100", 1595=>x"3000", 1596=>x"3200",
---- 1597=>x"3300", 1598=>x"3b00", 1599=>x"4000", 1600=>x"3500", 1601=>x"3400", 1602=>x"3200", 1603=>x"2d00",
---- 1604=>x"3100", 1605=>x"3a00", 1606=>x"3900", 1607=>x"3c00", 1608=>x"3900", 1609=>x"3900", 1610=>x"3200",
---- 1611=>x"ce00", 1612=>x"3300", 1613=>x"3600", 1614=>x"3600", 1615=>x"3900", 1616=>x"3c00", 1617=>x"4600",
---- 1618=>x"3300", 1619=>x"3400", 1620=>x"3100", 1621=>x"3500", 1622=>x"3600", 1623=>x"3800", 1624=>x"3900",
---- 1625=>x"4000", 1626=>x"3a00", 1627=>x"3600", 1628=>x"3300", 1629=>x"3200", 1630=>x"3e00", 1631=>x"3e00",
---- 1632=>x"4000", 1633=>x"3d00", 1634=>x"3900", 1635=>x"3500", 1636=>x"3400", 1637=>x"3000", 1638=>x"3b00",
---- 1639=>x"3e00", 1640=>x"3e00", 1641=>x"4300", 1642=>x"3500", 1643=>x"3000", 1644=>x"3600", 1645=>x"3400",
---- 1646=>x"3e00", 1647=>x"4500", 1648=>x"3e00", 1649=>x"4500", 1650=>x"3c00", 1651=>x"3600", 1652=>x"3800",
---- 1653=>x"3700", 1654=>x"4600", 1655=>x"4e00", 1656=>x"3c00", 1657=>x"4600", 1658=>x"3a00", 1659=>x"3a00",
---- 1660=>x"3800", 1661=>x"3400", 1662=>x"3f00", 1663=>x"4a00", 1664=>x"3c00", 1665=>x"4800", 1666=>x"3700",
---- 1667=>x"3100", 1668=>x"2e00", 1669=>x"2c00", 1670=>x"3700", 1671=>x"4700", 1672=>x"3b00", 1673=>x"4200",
---- 1674=>x"3600", 1675=>x"3800", 1676=>x"3100", 1677=>x"2a00", 1678=>x"3800", 1679=>x"4800", 1680=>x"4300",
---- 1681=>x"4500", 1682=>x"3700", 1683=>x"3600", 1684=>x"3a00", 1685=>x"3000", 1686=>x"3300", 1687=>x"3e00",
---- 1688=>x"3f00", 1689=>x"5000", 1690=>x"3300", 1691=>x"3700", 1692=>x"3900", 1693=>x"2d00", 1694=>x"3700",
---- 1695=>x"3a00", 1696=>x"3e00", 1697=>x"4500", 1698=>x"3100", 1699=>x"3200", 1700=>x"3100", 1701=>x"2d00",
---- 1702=>x"3400", 1703=>x"3600", 1704=>x"3c00", 1705=>x"4000", 1706=>x"3000", 1707=>x"2e00", 1708=>x"3800",
---- 1709=>x"3900", 1710=>x"3500", 1711=>x"3a00", 1712=>x"4000", 1713=>x"3f00", 1714=>x"2d00", 1715=>x"2c00",
---- 1716=>x"3300", 1717=>x"3100", 1718=>x"3900", 1719=>x"4300", 1720=>x"3f00", 1721=>x"4100", 1722=>x"3400",
---- 1723=>x"2a00", 1724=>x"2d00", 1725=>x"3700", 1726=>x"3600", 1727=>x"4d00", 1728=>x"3900", 1729=>x"3800",
---- 1730=>x"3a00", 1731=>x"3200", 1732=>x"3100", 1733=>x"3b00", 1734=>x"3b00", 1735=>x"4e00", 1736=>x"3500",
---- 1737=>x"3300", 1738=>x"3500", 1739=>x"3a00", 1740=>x"3500", 1741=>x"3900", 1742=>x"ba00", 1743=>x"5c00",
---- 1744=>x"3500", 1745=>x"2f00", 1746=>x"3100", 1747=>x"3500", 1748=>x"3b00", 1749=>x"3e00", 1750=>x"5200",
---- 1751=>x"6e00", 1752=>x"3500", 1753=>x"3100", 1754=>x"3300", 1755=>x"3500", 1756=>x"4300", 1757=>x"4600",
---- 1758=>x"5a00", 1759=>x"7600", 1760=>x"3400", 1761=>x"3100", 1762=>x"3200", 1763=>x"3b00", 1764=>x"4600",
---- 1765=>x"4c00", 1766=>x"6200", 1767=>x"7800", 1768=>x"3400", 1769=>x"2f00", 1770=>x"3000", 1771=>x"4100",
---- 1772=>x"4800", 1773=>x"5000", 1774=>x"6600", 1775=>x"7900", 1776=>x"3000", 1777=>x"3000", 1778=>x"3200",
---- 1779=>x"4500", 1780=>x"4e00", 1781=>x"5800", 1782=>x"6d00", 1783=>x"7d00", 1784=>x"2f00", 1785=>x"3400",
---- 1786=>x"3c00", 1787=>x"4700", 1788=>x"5300", 1789=>x"6000", 1790=>x"7400", 1791=>x"7c00", 1792=>x"2d00",
---- 1793=>x"3400", 1794=>x"4300", 1795=>x"4e00", 1796=>x"5900", 1797=>x"6400", 1798=>x"7600", 1799=>x"7b00",
---- 1800=>x"2c00", 1801=>x"3a00", 1802=>x"4b00", 1803=>x"5400", 1804=>x"5e00", 1805=>x"6b00", 1806=>x"7800",
---- 1807=>x"7e00", 1808=>x"3100", 1809=>x"3c00", 1810=>x"4f00", 1811=>x"5600", 1812=>x"6600", 1813=>x"6b00",
---- 1814=>x"7700", 1815=>x"7a00", 1816=>x"3600", 1817=>x"4800", 1818=>x"5200", 1819=>x"5700", 1820=>x"6a00",
---- 1821=>x"7000", 1822=>x"7600", 1823=>x"7c00", 1824=>x"3900", 1825=>x"4a00", 1826=>x"5900", 1827=>x"6100",
---- 1828=>x"6f00", 1829=>x"7700", 1830=>x"7800", 1831=>x"7c00", 1832=>x"4000", 1833=>x"4b00", 1834=>x"5900",
---- 1835=>x"6d00", 1836=>x"7100", 1837=>x"7400", 1838=>x"7900", 1839=>x"7f00", 1840=>x"4600", 1841=>x"4f00",
---- 1842=>x"5f00", 1843=>x"6e00", 1844=>x"7200", 1845=>x"7500", 1846=>x"7800", 1847=>x"7e00", 1848=>x"4800",
---- 1849=>x"5600", 1850=>x"6900", 1851=>x"7000", 1852=>x"7500", 1853=>x"7400", 1854=>x"7a00", 1855=>x"7e00",
---- 1856=>x"4e00", 1857=>x"5f00", 1858=>x"7200", 1859=>x"7300", 1860=>x"7300", 1861=>x"7400", 1862=>x"7800",
---- 1863=>x"7c00", 1864=>x"5600", 1865=>x"6a00", 1866=>x"7300", 1867=>x"7800", 1868=>x"7600", 1869=>x"7400",
---- 1870=>x"7500", 1871=>x"7700", 1872=>x"5f00", 1873=>x"7100", 1874=>x"7800", 1875=>x"7800", 1876=>x"7700",
---- 1877=>x"7700", 1878=>x"7700", 1879=>x"7700", 1880=>x"6700", 1881=>x"7300", 1882=>x"7400", 1883=>x"7500",
---- 1884=>x"7600", 1885=>x"7800", 1886=>x"7800", 1887=>x"6a00", 1888=>x"6d00", 1889=>x"7200", 1890=>x"7300",
---- 1891=>x"7400", 1892=>x"8900", 1893=>x"7700", 1894=>x"7200", 1895=>x"4a00", 1896=>x"7100", 1897=>x"7400",
---- 1898=>x"7500", 1899=>x"7500", 1900=>x"7900", 1901=>x"7900", 1902=>x"5200", 1903=>x"2c00", 1904=>x"7500",
---- 1905=>x"7300", 1906=>x"7500", 1907=>x"7700", 1908=>x"7800", 1909=>x"6000", 1910=>x"3400", 1911=>x"2500",
---- 1912=>x"7600", 1913=>x"7500", 1914=>x"7600", 1915=>x"7a00", 1916=>x"6200", 1917=>x"2f00", 1918=>x"2a00",
---- 1919=>x"3400", 1920=>x"7400", 1921=>x"7300", 1922=>x"7800", 1923=>x"5f00", 1924=>x"2d00", 1925=>x"2000",
---- 1926=>x"2d00", 1927=>x"b200", 1928=>x"7800", 1929=>x"7500", 1930=>x"5400", 1931=>x"2c00", 1932=>x"2300",
---- 1933=>x"3000", 1934=>x"4a00", 1935=>x"6200", 1936=>x"5e00", 1937=>x"3e00", 1938=>x"2300", 1939=>x"2100",
---- 1940=>x"3700", 1941=>x"5500", 1942=>x"6100", 1943=>x"6c00", 1944=>x"2400", 1945=>x"2000", 1946=>x"3200",
---- 1947=>x"4900", 1948=>x"5f00", 1949=>x"6a00", 1950=>x"6f00", 1951=>x"7500", 1952=>x"3200", 1953=>x"4500",
---- 1954=>x"5a00", 1955=>x"6400", 1956=>x"6a00", 1957=>x"7100", 1958=>x"8700", 1959=>x"7800", 1960=>x"5a00",
---- 1961=>x"6200", 1962=>x"6700", 1963=>x"6b00", 1964=>x"7200", 1965=>x"7600", 1966=>x"8100", 1967=>x"7b00",
---- 1968=>x"6500", 1969=>x"7000", 1970=>x"7300", 1971=>x"7900", 1972=>x"7e00", 1973=>x"7d00", 1974=>x"7e00",
---- 1975=>x"7d00", 1976=>x"7000", 1977=>x"7600", 1978=>x"7a00", 1979=>x"7800", 1980=>x"7c00", 1981=>x"7900",
---- 1982=>x"7d00", 1983=>x"7f00", 1984=>x"8800", 1985=>x"7a00", 1986=>x"7a00", 1987=>x"7700", 1988=>x"7d00",
---- 1989=>x"7c00", 1990=>x"7d00", 1991=>x"8000", 1992=>x"7900", 1993=>x"7b00", 1994=>x"7d00", 1995=>x"7f00",
---- 1996=>x"7e00", 1997=>x"7f00", 1998=>x"7f00", 1999=>x"8100", 2000=>x"7a00", 2001=>x"7d00", 2002=>x"7d00",
---- 2003=>x"7d00", 2004=>x"7f00", 2005=>x"8000", 2006=>x"8200", 2007=>x"7f00", 2008=>x"7a00", 2009=>x"7d00",
---- 2010=>x"7d00", 2011=>x"7e00", 2012=>x"8300", 2013=>x"8000", 2014=>x"7f00", 2015=>x"7c00", 2016=>x"7900",
---- 2017=>x"7c00", 2018=>x"8100", 2019=>x"8000", 2020=>x"7c00", 2021=>x"7e00", 2022=>x"7d00", 2023=>x"7c00",
---- 2024=>x"7900", 2025=>x"7a00", 2026=>x"7e00", 2027=>x"8100", 2028=>x"7f00", 2029=>x"7d00", 2030=>x"7f00",
---- 2031=>x"8000", 2032=>x"7d00", 2033=>x"7d00", 2034=>x"7d00", 2035=>x"7d00", 2036=>x"7e00", 2037=>x"7e00",
---- 2038=>x"8100", 2039=>x"8100", 2040=>x"7b00", 2041=>x"7d00", 2042=>x"7f00", 2043=>x"8000", 2044=>x"7e00",
---- 2045=>x"7f00", 2046=>x"8000", 2047=>x"8000"),
---- 14 => (0=>x"8200", 1=>x"8500", 2=>x"8700", 3=>x"8400", 4=>x"8400", 5=>x"8400", 6=>x"8300", 7=>x"8400",
---- 8=>x"8200", 9=>x"8500", 10=>x"8600", 11=>x"8400", 12=>x"8400", 13=>x"8400", 14=>x"8300",
---- 15=>x"8400", 16=>x"8200", 17=>x"8100", 18=>x"8600", 19=>x"8400", 20=>x"8200", 21=>x"8300",
---- 22=>x"8200", 23=>x"8300", 24=>x"8100", 25=>x"8300", 26=>x"8700", 27=>x"8200", 28=>x"8100",
---- 29=>x"8000", 30=>x"7e00", 31=>x"8400", 32=>x"8200", 33=>x"8700", 34=>x"8500", 35=>x"8400",
---- 36=>x"8200", 37=>x"8000", 38=>x"8100", 39=>x"8400", 40=>x"8200", 41=>x"8100", 42=>x"8100",
---- 43=>x"8200", 44=>x"8000", 45=>x"8100", 46=>x"8200", 47=>x"8100", 48=>x"8200", 49=>x"8100",
---- 50=>x"8300", 51=>x"8400", 52=>x"8100", 53=>x"8000", 54=>x"8200", 55=>x"8300", 56=>x"8100",
---- 57=>x"8400", 58=>x"8200", 59=>x"8200", 60=>x"8000", 61=>x"7f00", 62=>x"8300", 63=>x"8200",
---- 64=>x"7e00", 65=>x"8400", 66=>x"8400", 67=>x"8400", 68=>x"8100", 69=>x"8100", 70=>x"8200",
---- 71=>x"8300", 72=>x"7f00", 73=>x"8400", 74=>x"8500", 75=>x"8300", 76=>x"8100", 77=>x"7f00",
---- 78=>x"8100", 79=>x"8400", 80=>x"8300", 81=>x"8300", 82=>x"8200", 83=>x"8300", 84=>x"8000",
---- 85=>x"7f00", 86=>x"8000", 87=>x"8200", 88=>x"8400", 89=>x"8200", 90=>x"8000", 91=>x"8100",
---- 92=>x"8000", 93=>x"7f00", 94=>x"8000", 95=>x"8000", 96=>x"7f00", 97=>x"8000", 98=>x"7f00",
---- 99=>x"8000", 100=>x"8000", 101=>x"7e00", 102=>x"7d00", 103=>x"8000", 104=>x"8000", 105=>x"7d00",
---- 106=>x"7e00", 107=>x"7e00", 108=>x"8000", 109=>x"7d00", 110=>x"7c00", 111=>x"7e00", 112=>x"7d00",
---- 113=>x"7d00", 114=>x"7c00", 115=>x"7c00", 116=>x"8300", 117=>x"7e00", 118=>x"7f00", 119=>x"7f00",
---- 120=>x"7f00", 121=>x"7e00", 122=>x"7d00", 123=>x"7f00", 124=>x"7c00", 125=>x"7b00", 126=>x"7e00",
---- 127=>x"7f00", 128=>x"7d00", 129=>x"7b00", 130=>x"7d00", 131=>x"7e00", 132=>x"7e00", 133=>x"7e00",
---- 134=>x"7c00", 135=>x"7c00", 136=>x"7d00", 137=>x"8100", 138=>x"7d00", 139=>x"7a00", 140=>x"7a00",
---- 141=>x"7c00", 142=>x"7a00", 143=>x"7c00", 144=>x"7c00", 145=>x"7f00", 146=>x"7b00", 147=>x"7900",
---- 148=>x"7a00", 149=>x"7700", 150=>x"7700", 151=>x"7c00", 152=>x"7d00", 153=>x"7900", 154=>x"7700",
---- 155=>x"7800", 156=>x"7800", 157=>x"7600", 158=>x"7900", 159=>x"7900", 160=>x"7900", 161=>x"7800",
---- 162=>x"7800", 163=>x"7900", 164=>x"7900", 165=>x"7700", 166=>x"7900", 167=>x"7800", 168=>x"7400",
---- 169=>x"7700", 170=>x"7500", 171=>x"7600", 172=>x"7400", 173=>x"7700", 174=>x"7500", 175=>x"7500",
---- 176=>x"8a00", 177=>x"8800", 178=>x"8900", 179=>x"8000", 180=>x"7d00", 181=>x"7b00", 182=>x"7400",
---- 183=>x"7200", 184=>x"a400", 185=>x"b100", 186=>x"ac00", 187=>x"a800", 188=>x"aa00", 189=>x"ab00",
---- 190=>x"a300", 191=>x"9f00", 192=>x"b000", 193=>x"ac00", 194=>x"ab00", 195=>x"b100", 196=>x"b700",
---- 197=>x"b800", 198=>x"bc00", 199=>x"bc00", 200=>x"b200", 201=>x"b600", 202=>x"b200", 203=>x"b100",
---- 204=>x"b000", 205=>x"b800", 206=>x"b100", 207=>x"b400", 208=>x"b400", 209=>x"b700", 210=>x"b500",
---- 211=>x"b200", 212=>x"b300", 213=>x"ae00", 214=>x"a700", 215=>x"aa00", 216=>x"b100", 217=>x"b200",
---- 218=>x"b500", 219=>x"b400", 220=>x"b000", 221=>x"ac00", 222=>x"ac00", 223=>x"ac00", 224=>x"a300",
---- 225=>x"ae00", 226=>x"b500", 227=>x"b300", 228=>x"b000", 229=>x"b300", 230=>x"b100", 231=>x"af00",
---- 232=>x"a600", 233=>x"a300", 234=>x"b000", 235=>x"af00", 236=>x"a700", 237=>x"af00", 238=>x"4b00",
---- 239=>x"b100", 240=>x"5900", 241=>x"ac00", 242=>x"a700", 243=>x"a300", 244=>x"aa00", 245=>x"b200",
---- 246=>x"b400", 247=>x"b100", 248=>x"a600", 249=>x"a700", 250=>x"a700", 251=>x"ab00", 252=>x"af00",
---- 253=>x"b500", 254=>x"b400", 255=>x"b200", 256=>x"a200", 257=>x"a000", 258=>x"ae00", 259=>x"ad00",
---- 260=>x"ac00", 261=>x"b000", 262=>x"b600", 263=>x"bd00", 264=>x"ab00", 265=>x"ae00", 266=>x"ab00",
---- 267=>x"a900", 268=>x"ae00", 269=>x"b100", 270=>x"b800", 271=>x"ba00", 272=>x"a500", 273=>x"ae00",
---- 274=>x"af00", 275=>x"b000", 276=>x"5000", 277=>x"b200", 278=>x"b400", 279=>x"b400", 280=>x"a300",
---- 281=>x"5200", 282=>x"af00", 283=>x"b200", 284=>x"ae00", 285=>x"af00", 286=>x"b500", 287=>x"ae00",
---- 288=>x"a400", 289=>x"a800", 290=>x"a700", 291=>x"ac00", 292=>x"ab00", 293=>x"ae00", 294=>x"b300",
---- 295=>x"b600", 296=>x"9f00", 297=>x"a100", 298=>x"a200", 299=>x"a500", 300=>x"a800", 301=>x"af00",
---- 302=>x"b600", 303=>x"b500", 304=>x"9b00", 305=>x"9e00", 306=>x"9f00", 307=>x"ac00", 308=>x"ac00",
---- 309=>x"b300", 310=>x"b500", 311=>x"b300", 312=>x"9b00", 313=>x"a100", 314=>x"a700", 315=>x"aa00",
---- 316=>x"ae00", 317=>x"4900", 318=>x"b600", 319=>x"b900", 320=>x"a200", 321=>x"9800", 322=>x"a400",
---- 323=>x"b000", 324=>x"b000", 325=>x"b500", 326=>x"be00", 327=>x"bc00", 328=>x"9700", 329=>x"a100",
---- 330=>x"a600", 331=>x"a600", 332=>x"b300", 333=>x"be00", 334=>x"b300", 335=>x"b400", 336=>x"9f00",
---- 337=>x"6300", 338=>x"a300", 339=>x"ab00", 340=>x"ac00", 341=>x"b600", 342=>x"ba00", 343=>x"ba00",
---- 344=>x"9b00", 345=>x"9d00", 346=>x"a800", 347=>x"a500", 348=>x"b000", 349=>x"bc00", 350=>x"af00",
---- 351=>x"b200", 352=>x"9d00", 353=>x"9800", 354=>x"a300", 355=>x"ab00", 356=>x"a700", 357=>x"ad00",
---- 358=>x"b700", 359=>x"b600", 360=>x"9600", 361=>x"9c00", 362=>x"a300", 363=>x"9c00", 364=>x"ab00",
---- 365=>x"b700", 366=>x"b100", 367=>x"b000", 368=>x"9400", 369=>x"9800", 370=>x"a200", 371=>x"ac00",
---- 372=>x"ae00", 373=>x"4f00", 374=>x"b500", 375=>x"b200", 376=>x"9100", 377=>x"9b00", 378=>x"a700",
---- 379=>x"a300", 380=>x"af00", 381=>x"af00", 382=>x"ab00", 383=>x"9a00", 384=>x"9c00", 385=>x"9b00",
---- 386=>x"a000", 387=>x"5300", 388=>x"b200", 389=>x"9b00", 390=>x"8800", 391=>x"9300", 392=>x"9000",
---- 393=>x"9900", 394=>x"ac00", 395=>x"a900", 396=>x"9100", 397=>x"7e00", 398=>x"9800", 399=>x"ba00",
---- 400=>x"9400", 401=>x"a100", 402=>x"a200", 403=>x"8e00", 404=>x"8500", 405=>x"a500", 406=>x"c700",
---- 407=>x"c100", 408=>x"8700", 409=>x"9000", 410=>x"8600", 411=>x"8c00", 412=>x"b200", 413=>x"c600",
---- 414=>x"c700", 415=>x"3a00", 416=>x"8000", 417=>x"8200", 418=>x"6600", 419=>x"b100", 420=>x"c200",
---- 421=>x"be00", 422=>x"c600", 423=>x"c600", 424=>x"8d00", 425=>x"b300", 426=>x"b900", 427=>x"b000",
---- 428=>x"b500", 429=>x"c500", 430=>x"c500", 431=>x"ca00", 432=>x"ae00", 433=>x"c300", 434=>x"ba00",
---- 435=>x"b500", 436=>x"bc00", 437=>x"c000", 438=>x"c300", 439=>x"c100", 440=>x"b500", 441=>x"b900",
---- 442=>x"c700", 443=>x"bf00", 444=>x"bf00", 445=>x"b700", 446=>x"bb00", 447=>x"b900", 448=>x"ba00",
---- 449=>x"4000", 450=>x"c200", 451=>x"3d00", 452=>x"b500", 453=>x"b900", 454=>x"b400", 455=>x"bd00",
---- 456=>x"b800", 457=>x"b900", 458=>x"b700", 459=>x"b700", 460=>x"bd00", 461=>x"bb00", 462=>x"c100",
---- 463=>x"b800", 464=>x"b900", 465=>x"ad00", 466=>x"ad00", 467=>x"ae00", 468=>x"be00", 469=>x"c400",
---- 470=>x"bf00", 471=>x"af00", 472=>x"b000", 473=>x"b200", 474=>x"ad00", 475=>x"b100", 476=>x"b700",
---- 477=>x"b100", 478=>x"ad00", 479=>x"b800", 480=>x"ab00", 481=>x"b100", 482=>x"b900", 483=>x"ae00",
---- 484=>x"a000", 485=>x"a300", 486=>x"b900", 487=>x"bd00", 488=>x"bb00", 489=>x"ba00", 490=>x"a900",
---- 491=>x"a800", 492=>x"b100", 493=>x"b700", 494=>x"b000", 495=>x"b400", 496=>x"ac00", 497=>x"a600",
---- 498=>x"ac00", 499=>x"bd00", 500=>x"bb00", 501=>x"b200", 502=>x"ae00", 503=>x"a800", 504=>x"a900",
---- 505=>x"b300", 506=>x"b200", 507=>x"4b00", 508=>x"b800", 509=>x"b200", 510=>x"af00", 511=>x"b500",
---- 512=>x"ba00", 513=>x"b900", 514=>x"b200", 515=>x"ae00", 516=>x"ae00", 517=>x"b400", 518=>x"be00",
---- 519=>x"bd00", 520=>x"b400", 521=>x"b700", 522=>x"b300", 523=>x"aa00", 524=>x"b300", 525=>x"ba00",
---- 526=>x"bd00", 527=>x"b900", 528=>x"b500", 529=>x"ac00", 530=>x"b600", 531=>x"ba00", 532=>x"b400",
---- 533=>x"b100", 534=>x"b500", 535=>x"bd00", 536=>x"b500", 537=>x"b900", 538=>x"b400", 539=>x"bf00",
---- 540=>x"b300", 541=>x"a900", 542=>x"af00", 543=>x"b200", 544=>x"af00", 545=>x"b700", 546=>x"b000",
---- 547=>x"ad00", 548=>x"b500", 549=>x"b200", 550=>x"a800", 551=>x"b400", 552=>x"ae00", 553=>x"a600",
---- 554=>x"aa00", 555=>x"ab00", 556=>x"a800", 557=>x"b900", 558=>x"bb00", 559=>x"b000", 560=>x"a700",
---- 561=>x"a800", 562=>x"a400", 563=>x"a300", 564=>x"b400", 565=>x"b700", 566=>x"bc00", 567=>x"bb00",
---- 568=>x"5900", 569=>x"a500", 570=>x"af00", 571=>x"b100", 572=>x"a500", 573=>x"b700", 574=>x"b200",
---- 575=>x"af00", 576=>x"ac00", 577=>x"ab00", 578=>x"a700", 579=>x"b800", 580=>x"ac00", 581=>x"9f00",
---- 582=>x"a400", 583=>x"9600", 584=>x"b600", 585=>x"b700", 586=>x"ac00", 587=>x"a300", 588=>x"b200",
---- 589=>x"9a00", 590=>x"6300", 591=>x"ac00", 592=>x"b100", 593=>x"b700", 594=>x"b500", 595=>x"a000",
---- 596=>x"9700", 597=>x"9b00", 598=>x"ad00", 599=>x"ba00", 600=>x"a200", 601=>x"a300", 602=>x"a600",
---- 603=>x"9900", 604=>x"a400", 605=>x"b100", 606=>x"a600", 607=>x"ae00", 608=>x"a900", 609=>x"8e00",
---- 610=>x"9300", 611=>x"ad00", 612=>x"b500", 613=>x"b300", 614=>x"ae00", 615=>x"a100", 616=>x"9700",
---- 617=>x"9600", 618=>x"a500", 619=>x"b300", 620=>x"b200", 621=>x"b000", 622=>x"ab00", 623=>x"a700",
---- 624=>x"9d00", 625=>x"b000", 626=>x"af00", 627=>x"aa00", 628=>x"a700", 629=>x"a500", 630=>x"aa00",
---- 631=>x"a900", 632=>x"aa00", 633=>x"ac00", 634=>x"b100", 635=>x"ab00", 636=>x"a500", 637=>x"a200",
---- 638=>x"a500", 639=>x"a900", 640=>x"6000", 641=>x"a800", 642=>x"a500", 643=>x"a300", 644=>x"ab00",
---- 645=>x"a800", 646=>x"a200", 647=>x"a700", 648=>x"9e00", 649=>x"9700", 650=>x"9900", 651=>x"9e00",
---- 652=>x"a200", 653=>x"b100", 654=>x"ac00", 655=>x"9e00", 656=>x"a300", 657=>x"9d00", 658=>x"9600",
---- 659=>x"9f00", 660=>x"a200", 661=>x"a200", 662=>x"a900", 663=>x"9d00", 664=>x"9200", 665=>x"9e00",
---- 666=>x"a900", 667=>x"9600", 668=>x"9900", 669=>x"9b00", 670=>x"9300", 671=>x"9100", 672=>x"9800",
---- 673=>x"9600", 674=>x"a600", 675=>x"a300", 676=>x"9c00", 677=>x"9d00", 678=>x"9400", 679=>x"8c00",
---- 680=>x"8800", 681=>x"8b00", 682=>x"8700", 683=>x"9200", 684=>x"9a00", 685=>x"9900", 686=>x"9300",
---- 687=>x"8500", 688=>x"6c00", 689=>x"6600", 690=>x"6200", 691=>x"6200", 692=>x"6c00", 693=>x"8700",
---- 694=>x"9700", 695=>x"7400", 696=>x"8900", 697=>x"7700", 698=>x"7400", 699=>x"6a00", 700=>x"6300",
---- 701=>x"5900", 702=>x"6700", 703=>x"6200", 704=>x"7e00", 705=>x"7a00", 706=>x"7200", 707=>x"6c00",
---- 708=>x"6b00", 709=>x"5d00", 710=>x"4500", 711=>x"5300", 712=>x"6300", 713=>x"6900", 714=>x"5f00",
---- 715=>x"4c00", 716=>x"4300", 717=>x"4800", 718=>x"3f00", 719=>x"4a00", 720=>x"6c00", 721=>x"9700",
---- 722=>x"5700", 723=>x"5e00", 724=>x"6600", 725=>x"5200", 726=>x"5000", 727=>x"6700", 728=>x"7b00",
---- 729=>x"6500", 730=>x"7200", 731=>x"8b00", 732=>x"7e00", 733=>x"6700", 734=>x"5100", 735=>x"5e00",
---- 736=>x"6f00", 737=>x"6c00", 738=>x"7b00", 739=>x"7000", 740=>x"5d00", 741=>x"4500", 742=>x"4500",
---- 743=>x"4e00", 744=>x"7400", 745=>x"5700", 746=>x"4500", 747=>x"3a00", 748=>x"3900", 749=>x"3900",
---- 750=>x"3700", 751=>x"3a00", 752=>x"5000", 753=>x"4700", 754=>x"4700", 755=>x"3c00", 756=>x"3600",
---- 757=>x"3c00", 758=>x"3b00", 759=>x"3b00", 760=>x"5d00", 761=>x"4f00", 762=>x"4600", 763=>x"3500",
---- 764=>x"3300", 765=>x"3500", 766=>x"3300", 767=>x"5200", 768=>x"4200", 769=>x"3700", 770=>x"3600",
---- 771=>x"2f00", 772=>x"3700", 773=>x"2d00", 774=>x"3e00", 775=>x"7a00", 776=>x"2b00", 777=>x"3300",
---- 778=>x"3900", 779=>x"2e00", 780=>x"3400", 781=>x"2b00", 782=>x"5700", 783=>x"7c00", 784=>x"3400",
---- 785=>x"3f00", 786=>x"2b00", 787=>x"2a00", 788=>x"3100", 789=>x"3a00", 790=>x"7c00", 791=>x"6500",
---- 792=>x"4a00", 793=>x"3700", 794=>x"2400", 795=>x"2800", 796=>x"3700", 797=>x"5c00", 798=>x"8d00",
---- 799=>x"4000", 800=>x"4900", 801=>x"2400", 802=>x"2500", 803=>x"2a00", 804=>x"4a00", 805=>x"5b00",
---- 806=>x"5900", 807=>x"2f00", 808=>x"2c00", 809=>x"2600", 810=>x"2700", 811=>x"3400", 812=>x"5d00",
---- 813=>x"5000", 814=>x"4500", 815=>x"2700", 816=>x"2000", 817=>x"2800", 818=>x"2900", 819=>x"3900",
---- 820=>x"6100", 821=>x"4b00", 822=>x"3900", 823=>x"2c00", 824=>x"2300", 825=>x"2b00", 826=>x"2e00",
---- 827=>x"c500", 828=>x"5300", 829=>x"4b00", 830=>x"3b00", 831=>x"2a00", 832=>x"2100", 833=>x"2d00",
---- 834=>x"4f00", 835=>x"4000", 836=>x"3400", 837=>x"3900", 838=>x"3900", 839=>x"3b00", 840=>x"2d00",
---- 841=>x"3f00", 842=>x"5300", 843=>x"3000", 844=>x"2e00", 845=>x"3200", 846=>x"3200", 847=>x"3800",
---- 848=>x"4d00", 849=>x"4600", 850=>x"2f00", 851=>x"2e00", 852=>x"2f00", 853=>x"2f00", 854=>x"2f00",
---- 855=>x"3100", 856=>x"6800", 857=>x"4600", 858=>x"2a00", 859=>x"2e00", 860=>x"3200", 861=>x"2e00",
---- 862=>x"3000", 863=>x"3100", 864=>x"7e00", 865=>x"5700", 866=>x"2700", 867=>x"2c00", 868=>x"3200",
---- 869=>x"3100", 870=>x"3000", 871=>x"2c00", 872=>x"7d00", 873=>x"7c00", 874=>x"4300", 875=>x"2b00",
---- 876=>x"2900", 877=>x"2e00", 878=>x"2d00", 879=>x"2a00", 880=>x"5100", 881=>x"8a00", 882=>x"6f00",
---- 883=>x"5700", 884=>x"5700", 885=>x"3c00", 886=>x"2400", 887=>x"2700", 888=>x"3600", 889=>x"8600",
---- 890=>x"5e00", 891=>x"3900", 892=>x"4d00", 893=>x"3e00", 894=>x"2700", 895=>x"2400", 896=>x"3300",
---- 897=>x"8200", 898=>x"5f00", 899=>x"2000", 900=>x"2500", 901=>x"2400", 902=>x"2300", 903=>x"2200",
---- 904=>x"2400", 905=>x"5f00", 906=>x"7600", 907=>x"2700", 908=>x"2700", 909=>x"2300", 910=>x"2300",
---- 911=>x"1d00", 912=>x"d300", 913=>x"3f00", 914=>x"7c00", 915=>x"3300", 916=>x"1f00", 917=>x"2100",
---- 918=>x"2000", 919=>x"3600", 920=>x"5300", 921=>x"4d00", 922=>x"9400", 923=>x"5e00", 924=>x"1e00",
---- 925=>x"1c00", 926=>x"2e00", 927=>x"7f00", 928=>x"3e00", 929=>x"3b00", 930=>x"8a00", 931=>x"5d00",
---- 932=>x"1700", 933=>x"2500", 934=>x"7000", 935=>x"9e00", 936=>x"2100", 937=>x"1b00", 938=>x"5500",
---- 939=>x"7a00", 940=>x"2200", 941=>x"5d00", 942=>x"9c00", 943=>x"7e00", 944=>x"1d00", 945=>x"1f00",
---- 946=>x"2e00", 947=>x"6e00", 948=>x"6400", 949=>x"9500", 950=>x"8900", 951=>x"9400", 952=>x"1b00",
---- 953=>x"1f00", 954=>x"1e00", 955=>x"4500", 956=>x"8c00", 957=>x"8800", 958=>x"6c00", 959=>x"8700",
---- 960=>x"2800", 961=>x"2000", 962=>x"2d00", 963=>x"7200", 964=>x"7700", 965=>x"5a00", 966=>x"7a00",
---- 967=>x"b100", 968=>x"3400", 969=>x"2200", 970=>x"6300", 971=>x"9700", 972=>x"5d00", 973=>x"6a00",
---- 974=>x"b300", 975=>x"ae00", 976=>x"2100", 977=>x"4c00", 978=>x"9b00", 979=>x"7600", 980=>x"5d00",
---- 981=>x"a900", 982=>x"bb00", 983=>x"a300", 984=>x"3400", 985=>x"8e00", 986=>x"8300", 987=>x"a500",
---- 988=>x"9200", 989=>x"bc00", 990=>x"a700", 991=>x"ac00", 992=>x"7300", 993=>x"9600", 994=>x"5b00",
---- 995=>x"8000", 996=>x"b600", 997=>x"a800", 998=>x"ad00", 999=>x"b400", 1000=>x"a100", 1001=>x"7300",
---- 1002=>x"7300", 1003=>x"b900", 1004=>x"ab00", 1005=>x"a700", 1006=>x"b400", 1007=>x"4200", 1008=>x"9600",
---- 1009=>x"7100", 1010=>x"a900", 1011=>x"b700", 1012=>x"a400", 1013=>x"af00", 1014=>x"b700", 1015=>x"c400",
---- 1016=>x"6900", 1017=>x"9d00", 1018=>x"bd00", 1019=>x"a500", 1020=>x"ac00", 1021=>x"b600", 1022=>x"bf00",
---- 1023=>x"c700", 1024=>x"8000", 1025=>x"c000", 1026=>x"aa00", 1027=>x"a900", 1028=>x"b400", 1029=>x"c000",
---- 1030=>x"c900", 1031=>x"c700", 1032=>x"b500", 1033=>x"b200", 1034=>x"aa00", 1035=>x"b000", 1036=>x"bb00",
---- 1037=>x"c700", 1038=>x"ca00", 1039=>x"c100", 1040=>x"bf00", 1041=>x"a500", 1042=>x"b000", 1043=>x"b400",
---- 1044=>x"bc00", 1045=>x"c900", 1046=>x"c500", 1047=>x"bf00", 1048=>x"ac00", 1049=>x"a800", 1050=>x"b000",
---- 1051=>x"b600", 1052=>x"c100", 1053=>x"cc00", 1054=>x"c500", 1055=>x"be00", 1056=>x"a700", 1057=>x"b200",
---- 1058=>x"b200", 1059=>x"b600", 1060=>x"c700", 1061=>x"ca00", 1062=>x"c300", 1063=>x"c500", 1064=>x"b200",
---- 1065=>x"b800", 1066=>x"b600", 1067=>x"c100", 1068=>x"cd00", 1069=>x"c700", 1070=>x"c700", 1071=>x"cc00",
---- 1072=>x"a000", 1073=>x"b100", 1074=>x"bd00", 1075=>x"c900", 1076=>x"c800", 1077=>x"c300", 1078=>x"cc00",
---- 1079=>x"9300", 1080=>x"b100", 1081=>x"be00", 1082=>x"c600", 1083=>x"c700", 1084=>x"c300", 1085=>x"ca00",
---- 1086=>x"9600", 1087=>x"6500", 1088=>x"bd00", 1089=>x"c600", 1090=>x"c800", 1091=>x"c400", 1092=>x"c600",
---- 1093=>x"9700", 1094=>x"6900", 1095=>x"7800", 1096=>x"c200", 1097=>x"c900", 1098=>x"c500", 1099=>x"c500",
---- 1100=>x"7100", 1101=>x"6200", 1102=>x"7a00", 1103=>x"7e00", 1104=>x"c900", 1105=>x"c700", 1106=>x"c800",
---- 1107=>x"8f00", 1108=>x"5b00", 1109=>x"7200", 1110=>x"7e00", 1111=>x"7f00", 1112=>x"c800", 1113=>x"cb00",
---- 1114=>x"9100", 1115=>x"5600", 1116=>x"6b00", 1117=>x"7a00", 1118=>x"8200", 1119=>x"8700", 1120=>x"ce00",
---- 1121=>x"9600", 1122=>x"4c00", 1123=>x"5f00", 1124=>x"7200", 1125=>x"7e00", 1126=>x"8300", 1127=>x"8800",
---- 1128=>x"9e00", 1129=>x"4b00", 1130=>x"5a00", 1131=>x"6c00", 1132=>x"7700", 1133=>x"7f00", 1134=>x"8600",
---- 1135=>x"8c00", 1136=>x"4900", 1137=>x"5400", 1138=>x"9500", 1139=>x"6f00", 1140=>x"7600", 1141=>x"8000",
---- 1142=>x"8600", 1143=>x"8b00", 1144=>x"4700", 1145=>x"6200", 1146=>x"7000", 1147=>x"7400", 1148=>x"7900",
---- 1149=>x"8400", 1150=>x"8700", 1151=>x"8900", 1152=>x"5700", 1153=>x"6600", 1154=>x"7000", 1155=>x"7800",
---- 1156=>x"7c00", 1157=>x"7d00", 1158=>x"8900", 1159=>x"8b00", 1160=>x"5800", 1161=>x"6d00", 1162=>x"7200",
---- 1163=>x"7700", 1164=>x"7d00", 1165=>x"8100", 1166=>x"8400", 1167=>x"8b00", 1168=>x"5b00", 1169=>x"6f00",
---- 1170=>x"7600", 1171=>x"7800", 1172=>x"7e00", 1173=>x"8000", 1174=>x"8400", 1175=>x"8c00", 1176=>x"6400",
---- 1177=>x"7100", 1178=>x"7900", 1179=>x"8400", 1180=>x"7d00", 1181=>x"8000", 1182=>x"8500", 1183=>x"8a00",
---- 1184=>x"6600", 1185=>x"7500", 1186=>x"7900", 1187=>x"7b00", 1188=>x"7c00", 1189=>x"7c00", 1190=>x"8300",
---- 1191=>x"8b00", 1192=>x"6b00", 1193=>x"7500", 1194=>x"7700", 1195=>x"7d00", 1196=>x"8000", 1197=>x"7d00",
---- 1198=>x"8400", 1199=>x"8600", 1200=>x"6a00", 1201=>x"7500", 1202=>x"7800", 1203=>x"7800", 1204=>x"8000",
---- 1205=>x"8500", 1206=>x"8500", 1207=>x"8300", 1208=>x"6700", 1209=>x"7300", 1210=>x"7b00", 1211=>x"7a00",
---- 1212=>x"7d00", 1213=>x"8300", 1214=>x"8400", 1215=>x"8800", 1216=>x"6500", 1217=>x"6f00", 1218=>x"7600",
---- 1219=>x"7d00", 1220=>x"8000", 1221=>x"8000", 1222=>x"8400", 1223=>x"8800", 1224=>x"6200", 1225=>x"6c00",
---- 1226=>x"7300", 1227=>x"7900", 1228=>x"8100", 1229=>x"8100", 1230=>x"8500", 1231=>x"7a00", 1232=>x"6400",
---- 1233=>x"6b00", 1234=>x"7400", 1235=>x"7b00", 1236=>x"7e00", 1237=>x"7e00", 1238=>x"8200", 1239=>x"8300",
---- 1240=>x"6200", 1241=>x"6c00", 1242=>x"7200", 1243=>x"7d00", 1244=>x"7c00", 1245=>x"7f00", 1246=>x"8300",
---- 1247=>x"8300", 1248=>x"6000", 1249=>x"6900", 1250=>x"7600", 1251=>x"7900", 1252=>x"7d00", 1253=>x"8100",
---- 1254=>x"8100", 1255=>x"8500", 1256=>x"5c00", 1257=>x"6900", 1258=>x"7200", 1259=>x"7600", 1260=>x"7e00",
---- 1261=>x"8000", 1262=>x"8200", 1263=>x"8500", 1264=>x"5900", 1265=>x"6b00", 1266=>x"7200", 1267=>x"7700",
---- 1268=>x"7c00", 1269=>x"7e00", 1270=>x"8000", 1271=>x"8300", 1272=>x"5d00", 1273=>x"6d00", 1274=>x"7400",
---- 1275=>x"7a00", 1276=>x"7c00", 1277=>x"8000", 1278=>x"8000", 1279=>x"8200", 1280=>x"6000", 1281=>x"6e00",
---- 1282=>x"7400", 1283=>x"7900", 1284=>x"7e00", 1285=>x"8000", 1286=>x"8200", 1287=>x"8000", 1288=>x"6000",
---- 1289=>x"6b00", 1290=>x"7400", 1291=>x"7900", 1292=>x"7b00", 1293=>x"7c00", 1294=>x"8100", 1295=>x"8000",
---- 1296=>x"6300", 1297=>x"6900", 1298=>x"7200", 1299=>x"7700", 1300=>x"7800", 1301=>x"7c00", 1302=>x"8000",
---- 1303=>x"8200", 1304=>x"6800", 1305=>x"7000", 1306=>x"7200", 1307=>x"7700", 1308=>x"7c00", 1309=>x"7a00",
---- 1310=>x"7f00", 1311=>x"8200", 1312=>x"6b00", 1313=>x"7000", 1314=>x"7400", 1315=>x"7800", 1316=>x"7d00",
---- 1317=>x"7c00", 1318=>x"7d00", 1319=>x"8300", 1320=>x"6c00", 1321=>x"7300", 1322=>x"7500", 1323=>x"7800",
---- 1324=>x"7b00", 1325=>x"7d00", 1326=>x"7f00", 1327=>x"8200", 1328=>x"6a00", 1329=>x"7000", 1330=>x"7700",
---- 1331=>x"7900", 1332=>x"7b00", 1333=>x"7c00", 1334=>x"7a00", 1335=>x"7f00", 1336=>x"6b00", 1337=>x"7300",
---- 1338=>x"7900", 1339=>x"7d00", 1340=>x"7d00", 1341=>x"7e00", 1342=>x"7f00", 1343=>x"8100", 1344=>x"6f00",
---- 1345=>x"7100", 1346=>x"7800", 1347=>x"7d00", 1348=>x"7d00", 1349=>x"7f00", 1350=>x"8000", 1351=>x"7f00",
---- 1352=>x"6900", 1353=>x"7100", 1354=>x"7500", 1355=>x"7800", 1356=>x"7d00", 1357=>x"7e00", 1358=>x"8200",
---- 1359=>x"8200", 1360=>x"6700", 1361=>x"7000", 1362=>x"7400", 1363=>x"7a00", 1364=>x"7d00", 1365=>x"8100",
---- 1366=>x"8100", 1367=>x"8200", 1368=>x"5e00", 1369=>x"6c00", 1370=>x"7300", 1371=>x"7b00", 1372=>x"7c00",
---- 1373=>x"8000", 1374=>x"7d00", 1375=>x"8000", 1376=>x"5900", 1377=>x"6900", 1378=>x"7200", 1379=>x"7600",
---- 1380=>x"7b00", 1381=>x"7f00", 1382=>x"7f00", 1383=>x"8200", 1384=>x"5300", 1385=>x"6400", 1386=>x"7000",
---- 1387=>x"7700", 1388=>x"7c00", 1389=>x"7d00", 1390=>x"8200", 1391=>x"8200", 1392=>x"4f00", 1393=>x"6300",
---- 1394=>x"6c00", 1395=>x"7100", 1396=>x"7900", 1397=>x"8000", 1398=>x"8300", 1399=>x"8100", 1400=>x"4800",
---- 1401=>x"5c00", 1402=>x"6b00", 1403=>x"7500", 1404=>x"7700", 1405=>x"7e00", 1406=>x"8500", 1407=>x"8100",
---- 1408=>x"4d00", 1409=>x"5a00", 1410=>x"6400", 1411=>x"7100", 1412=>x"7900", 1413=>x"7b00", 1414=>x"7f00",
---- 1415=>x"7f00", 1416=>x"4d00", 1417=>x"5800", 1418=>x"6400", 1419=>x"6e00", 1420=>x"7500", 1421=>x"7800",
---- 1422=>x"7d00", 1423=>x"7c00", 1424=>x"4b00", 1425=>x"4c00", 1426=>x"5e00", 1427=>x"6b00", 1428=>x"7300",
---- 1429=>x"7300", 1430=>x"7700", 1431=>x"7a00", 1432=>x"4200", 1433=>x"4b00", 1434=>x"5a00", 1435=>x"6700",
---- 1436=>x"6e00", 1437=>x"7100", 1438=>x"7400", 1439=>x"7500", 1440=>x"3f00", 1441=>x"4900", 1442=>x"5700",
---- 1443=>x"6300", 1444=>x"6b00", 1445=>x"6f00", 1446=>x"7400", 1447=>x"8c00", 1448=>x"4000", 1449=>x"4300",
---- 1450=>x"4f00", 1451=>x"5c00", 1452=>x"6800", 1453=>x"6900", 1454=>x"6a00", 1455=>x"6e00", 1456=>x"4100",
---- 1457=>x"4200", 1458=>x"4a00", 1459=>x"5100", 1460=>x"5f00", 1461=>x"6900", 1462=>x"6900", 1463=>x"6900",
---- 1464=>x"4200", 1465=>x"3a00", 1466=>x"4900", 1467=>x"5000", 1468=>x"5600", 1469=>x"9d00", 1470=>x"6700",
---- 1471=>x"6600", 1472=>x"4700", 1473=>x"3700", 1474=>x"4700", 1475=>x"5100", 1476=>x"5400", 1477=>x"5900",
---- 1478=>x"5d00", 1479=>x"6600", 1480=>x"4500", 1481=>x"3700", 1482=>x"3b00", 1483=>x"4700", 1484=>x"4600",
---- 1485=>x"5600", 1486=>x"5900", 1487=>x"6100", 1488=>x"4600", 1489=>x"3a00", 1490=>x"3500", 1491=>x"4600",
---- 1492=>x"4000", 1493=>x"4700", 1494=>x"5300", 1495=>x"5b00", 1496=>x"3e00", 1497=>x"3800", 1498=>x"3200",
---- 1499=>x"4900", 1500=>x"4600", 1501=>x"3300", 1502=>x"3f00", 1503=>x"5000", 1504=>x"3e00", 1505=>x"3e00",
---- 1506=>x"3400", 1507=>x"4500", 1508=>x"4b00", 1509=>x"3500", 1510=>x"3000", 1511=>x"3d00", 1512=>x"3800",
---- 1513=>x"4300", 1514=>x"3600", 1515=>x"3d00", 1516=>x"4c00", 1517=>x"3d00", 1518=>x"2e00", 1519=>x"2e00",
---- 1520=>x"3900", 1521=>x"4400", 1522=>x"3700", 1523=>x"3900", 1524=>x"4800", 1525=>x"4500", 1526=>x"3500",
---- 1527=>x"2d00", 1528=>x"3c00", 1529=>x"3f00", 1530=>x"3600", 1531=>x"3900", 1532=>x"4a00", 1533=>x"4a00",
---- 1534=>x"4200", 1535=>x"3300", 1536=>x"4000", 1537=>x"3f00", 1538=>x"3b00", 1539=>x"3700", 1540=>x"bb00",
---- 1541=>x"4900", 1542=>x"4800", 1543=>x"3d00", 1544=>x"4200", 1545=>x"4100", 1546=>x"3e00", 1547=>x"3600",
---- 1548=>x"3d00", 1549=>x"4600", 1550=>x"5100", 1551=>x"5000", 1552=>x"3b00", 1553=>x"3b00", 1554=>x"3d00",
---- 1555=>x"3500", 1556=>x"3400", 1557=>x"4000", 1558=>x"b300", 1559=>x"5000", 1560=>x"3b00", 1561=>x"3a00",
---- 1562=>x"3600", 1563=>x"3300", 1564=>x"2e00", 1565=>x"3900", 1566=>x"4600", 1567=>x"4e00", 1568=>x"3700",
---- 1569=>x"3f00", 1570=>x"3500", 1571=>x"3200", 1572=>x"3200", 1573=>x"3400", 1574=>x"4900", 1575=>x"5100",
---- 1576=>x"3900", 1577=>x"3900", 1578=>x"3400", 1579=>x"3900", 1580=>x"3400", 1581=>x"3500", 1582=>x"4900",
---- 1583=>x"5500", 1584=>x"3900", 1585=>x"3b00", 1586=>x"3b00", 1587=>x"3600", 1588=>x"3600", 1589=>x"3200",
---- 1590=>x"4300", 1591=>x"5300", 1592=>x"3a00", 1593=>x"3a00", 1594=>x"3a00", 1595=>x"3800", 1596=>x"3800",
---- 1597=>x"2f00", 1598=>x"3f00", 1599=>x"5200", 1600=>x"3b00", 1601=>x"4300", 1602=>x"4000", 1603=>x"3700",
---- 1604=>x"3600", 1605=>x"2e00", 1606=>x"3800", 1607=>x"4d00", 1608=>x"3f00", 1609=>x"4800", 1610=>x"4400",
---- 1611=>x"3900", 1612=>x"3900", 1613=>x"3200", 1614=>x"3800", 1615=>x"4900", 1616=>x"3c00", 1617=>x"4100",
---- 1618=>x"5000", 1619=>x"4000", 1620=>x"3900", 1621=>x"3300", 1622=>x"3800", 1623=>x"4d00", 1624=>x"4000",
---- 1625=>x"3c00", 1626=>x"5200", 1627=>x"4600", 1628=>x"3400", 1629=>x"3900", 1630=>x"3600", 1631=>x"4e00",
---- 1632=>x"4300", 1633=>x"4100", 1634=>x"5600", 1635=>x"5400", 1636=>x"3800", 1637=>x"3300", 1638=>x"3400",
---- 1639=>x"5000", 1640=>x"3e00", 1641=>x"4600", 1642=>x"5a00", 1643=>x"6200", 1644=>x"4400", 1645=>x"2e00",
---- 1646=>x"2b00", 1647=>x"4800", 1648=>x"3e00", 1649=>x"4900", 1650=>x"6000", 1651=>x"6a00", 1652=>x"5400",
---- 1653=>x"3400", 1654=>x"2d00", 1655=>x"3d00", 1656=>x"4000", 1657=>x"4b00", 1658=>x"6700", 1659=>x"6e00",
---- 1660=>x"5c00", 1661=>x"3800", 1662=>x"2b00", 1663=>x"3d00", 1664=>x"4100", 1665=>x"4c00", 1666=>x"6d00",
---- 1667=>x"7700", 1668=>x"6700", 1669=>x"3f00", 1670=>x"2900", 1671=>x"3600", 1672=>x"3d00", 1673=>x"5800",
---- 1674=>x"7400", 1675=>x"7600", 1676=>x"6b00", 1677=>x"4800", 1678=>x"2a00", 1679=>x"3600", 1680=>x"3a00",
---- 1681=>x"5d00", 1682=>x"7500", 1683=>x"7800", 1684=>x"6f00", 1685=>x"5000", 1686=>x"2800", 1687=>x"2f00",
---- 1688=>x"4400", 1689=>x"6700", 1690=>x"7500", 1691=>x"7600", 1692=>x"6e00", 1693=>x"4e00", 1694=>x"2900",
---- 1695=>x"2b00", 1696=>x"4e00", 1697=>x"6500", 1698=>x"6c00", 1699=>x"7200", 1700=>x"9200", 1701=>x"5000",
---- 1702=>x"2b00", 1703=>x"2d00", 1704=>x"5600", 1705=>x"6a00", 1706=>x"6f00", 1707=>x"6700", 1708=>x"9b00",
---- 1709=>x"5a00", 1710=>x"3200", 1711=>x"2f00", 1712=>x"6300", 1713=>x"7100", 1714=>x"6500", 1715=>x"6200",
---- 1716=>x"7000", 1717=>x"6000", 1718=>x"3200", 1719=>x"2f00", 1720=>x"5f00", 1721=>x"6300", 1722=>x"6300",
---- 1723=>x"7300", 1724=>x"7b00", 1725=>x"6000", 1726=>x"3400", 1727=>x"3000", 1728=>x"6200", 1729=>x"6c00",
---- 1730=>x"7600", 1731=>x"7b00", 1732=>x"7800", 1733=>x"6400", 1734=>x"3200", 1735=>x"3200", 1736=>x"7200",
---- 1737=>x"7800", 1738=>x"7b00", 1739=>x"7d00", 1740=>x"7800", 1741=>x"6800", 1742=>x"3100", 1743=>x"3900",
---- 1744=>x"7900", 1745=>x"7b00", 1746=>x"7d00", 1747=>x"7a00", 1748=>x"7a00", 1749=>x"6000", 1750=>x"3200",
---- 1751=>x"4200", 1752=>x"7c00", 1753=>x"7d00", 1754=>x"7b00", 1755=>x"7800", 1756=>x"7600", 1757=>x"5700",
---- 1758=>x"2d00", 1759=>x"4800", 1760=>x"7e00", 1761=>x"7d00", 1762=>x"7b00", 1763=>x"7c00", 1764=>x"7700",
---- 1765=>x"4f00", 1766=>x"2d00", 1767=>x"4b00", 1768=>x"7d00", 1769=>x"7c00", 1770=>x"7d00", 1771=>x"7b00",
---- 1772=>x"7a00", 1773=>x"4900", 1774=>x"2e00", 1775=>x"4e00", 1776=>x"7c00", 1777=>x"7a00", 1778=>x"8000",
---- 1779=>x"7f00", 1780=>x"7300", 1781=>x"4a00", 1782=>x"3400", 1783=>x"5500", 1784=>x"7c00", 1785=>x"8000",
---- 1786=>x"8100", 1787=>x"8100", 1788=>x"6e00", 1789=>x"4300", 1790=>x"3a00", 1791=>x"5a00", 1792=>x"8100",
---- 1793=>x"7f00", 1794=>x"8100", 1795=>x"8300", 1796=>x"6800", 1797=>x"3a00", 1798=>x"4200", 1799=>x"5f00",
---- 1800=>x"7e00", 1801=>x"8100", 1802=>x"8100", 1803=>x"7e00", 1804=>x"5d00", 1805=>x"3700", 1806=>x"4b00",
---- 1807=>x"6500", 1808=>x"7d00", 1809=>x"8100", 1810=>x"8000", 1811=>x"7800", 1812=>x"4f00", 1813=>x"3400",
---- 1814=>x"5100", 1815=>x"6500", 1816=>x"7f00", 1817=>x"7d00", 1818=>x"7d00", 1819=>x"7300", 1820=>x"4200",
---- 1821=>x"3a00", 1822=>x"5a00", 1823=>x"6500", 1824=>x"7d00", 1825=>x"7c00", 1826=>x"7b00", 1827=>x"6300",
---- 1828=>x"3700", 1829=>x"4200", 1830=>x"6000", 1831=>x"6b00", 1832=>x"7b00", 1833=>x"7b00", 1834=>x"7700",
---- 1835=>x"4e00", 1836=>x"3200", 1837=>x"5300", 1838=>x"6100", 1839=>x"7400", 1840=>x"7b00", 1841=>x"7d00",
---- 1842=>x"6900", 1843=>x"3c00", 1844=>x"3700", 1845=>x"5700", 1846=>x"6700", 1847=>x"7e00", 1848=>x"7c00",
---- 1849=>x"7a00", 1850=>x"5900", 1851=>x"3200", 1852=>x"4100", 1853=>x"5a00", 1854=>x"7000", 1855=>x"8800",
---- 1856=>x"7b00", 1857=>x"6c00", 1858=>x"3800", 1859=>x"3100", 1860=>x"5100", 1861=>x"6000", 1862=>x"7c00",
---- 1863=>x"8300", 1864=>x"7700", 1865=>x"4d00", 1866=>x"2900", 1867=>x"4000", 1868=>x"5a00", 1869=>x"6c00",
---- 1870=>x"8100", 1871=>x"8500", 1872=>x"6100", 1873=>x"3000", 1874=>x"2800", 1875=>x"4a00", 1876=>x"6800",
---- 1877=>x"7700", 1878=>x"8400", 1879=>x"8700", 1880=>x"3900", 1881=>x"2200", 1882=>x"3900", 1883=>x"5a00",
---- 1884=>x"6f00", 1885=>x"8100", 1886=>x"8600", 1887=>x"8700", 1888=>x"2700", 1889=>x"2a00", 1890=>x"4c00",
---- 1891=>x"6600", 1892=>x"7b00", 1893=>x"8300", 1894=>x"8400", 1895=>x"8900", 1896=>x"2900", 1897=>x"3e00",
---- 1898=>x"5d00", 1899=>x"7800", 1900=>x"8200", 1901=>x"8100", 1902=>x"8600", 1903=>x"8a00", 1904=>x"2e00",
---- 1905=>x"5300", 1906=>x"7100", 1907=>x"8100", 1908=>x"8100", 1909=>x"8200", 1910=>x"8900", 1911=>x"8600",
---- 1912=>x"4900", 1913=>x"6600", 1914=>x"7c00", 1915=>x"8100", 1916=>x"8100", 1917=>x"8500", 1918=>x"8800",
---- 1919=>x"8600", 1920=>x"6400", 1921=>x"7a00", 1922=>x"7f00", 1923=>x"7f00", 1924=>x"8300", 1925=>x"8400",
---- 1926=>x"8600", 1927=>x"8800", 1928=>x"7200", 1929=>x"7b00", 1930=>x"7d00", 1931=>x"8100", 1932=>x"8400",
---- 1933=>x"8100", 1934=>x"8700", 1935=>x"8700", 1936=>x"7a00", 1937=>x"7c00", 1938=>x"7f00", 1939=>x"7f00",
---- 1940=>x"8300", 1941=>x"8300", 1942=>x"8700", 1943=>x"8800", 1944=>x"7a00", 1945=>x"7c00", 1946=>x"7f00",
---- 1947=>x"8300", 1948=>x"8400", 1949=>x"8500", 1950=>x"8600", 1951=>x"8900", 1952=>x"7d00", 1953=>x"7d00",
---- 1954=>x"8000", 1955=>x"8300", 1956=>x"8200", 1957=>x"8400", 1958=>x"8800", 1959=>x"8700", 1960=>x"7a00",
---- 1961=>x"7d00", 1962=>x"8300", 1963=>x"8200", 1964=>x"8400", 1965=>x"8100", 1966=>x"8600", 1967=>x"8800",
---- 1968=>x"8000", 1969=>x"7f00", 1970=>x"8000", 1971=>x"7e00", 1972=>x"8200", 1973=>x"8300", 1974=>x"8500",
---- 1975=>x"8600", 1976=>x"7f00", 1977=>x"8000", 1978=>x"8000", 1979=>x"8100", 1980=>x"8200", 1981=>x"7f00",
---- 1982=>x"8200", 1983=>x"8600", 1984=>x"8200", 1985=>x"8300", 1986=>x"7d00", 1987=>x"8000", 1988=>x"7e00",
---- 1989=>x"7f00", 1990=>x"8200", 1991=>x"8700", 1992=>x"7f00", 1993=>x"8100", 1994=>x"8000", 1995=>x"8000",
---- 1996=>x"8000", 1997=>x"8000", 1998=>x"8700", 1999=>x"8400", 2000=>x"8000", 2001=>x"8100", 2002=>x"8000",
---- 2003=>x"8100", 2004=>x"8100", 2005=>x"8100", 2006=>x"8700", 2007=>x"8400", 2008=>x"8000", 2009=>x"8100",
---- 2010=>x"8000", 2011=>x"8500", 2012=>x"8500", 2013=>x"8100", 2014=>x"8300", 2015=>x"8300", 2016=>x"8000",
---- 2017=>x"8300", 2018=>x"8300", 2019=>x"8300", 2020=>x"8500", 2021=>x"8300", 2022=>x"8200", 2023=>x"8400",
---- 2024=>x"8100", 2025=>x"8400", 2026=>x"8300", 2027=>x"8200", 2028=>x"8400", 2029=>x"8500", 2030=>x"8100",
---- 2031=>x"8100", 2032=>x"8000", 2033=>x"8200", 2034=>x"8000", 2035=>x"8200", 2036=>x"8400", 2037=>x"8300",
---- 2038=>x"8200", 2039=>x"8200", 2040=>x"7e00", 2041=>x"8000", 2042=>x"8100", 2043=>x"8400", 2044=>x"8300",
---- 2045=>x"8500", 2046=>x"8400", 2047=>x"8200"),
---- 15 => (0=>x"8600", 1=>x"8500", 2=>x"8500", 3=>x"8700", 4=>x"8500", 5=>x"8400", 6=>x"8200", 7=>x"8500",
---- 8=>x"8600", 9=>x"8400", 10=>x"8600", 11=>x"8800", 12=>x"8500", 13=>x"8400", 14=>x"8100",
---- 15=>x"8500", 16=>x"8700", 17=>x"8500", 18=>x"8500", 19=>x"8700", 20=>x"8500", 21=>x"8400",
---- 22=>x"8200", 23=>x"8500", 24=>x"8400", 25=>x"8500", 26=>x"8600", 27=>x"8200", 28=>x"8400",
---- 29=>x"8300", 30=>x"8300", 31=>x"8400", 32=>x"8300", 33=>x"8400", 34=>x"8300", 35=>x"8300",
---- 36=>x"8000", 37=>x"8200", 38=>x"8300", 39=>x"8400", 40=>x"8200", 41=>x"8100", 42=>x"8400",
---- 43=>x"8400", 44=>x"8200", 45=>x"8200", 46=>x"8000", 47=>x"7f00", 48=>x"8500", 49=>x"8700",
---- 50=>x"8800", 51=>x"8500", 52=>x"8400", 53=>x"8300", 54=>x"8300", 55=>x"8100", 56=>x"8400",
---- 57=>x"8600", 58=>x"8600", 59=>x"8600", 60=>x"8500", 61=>x"8100", 62=>x"8400", 63=>x"8400",
---- 64=>x"8400", 65=>x"8800", 66=>x"8500", 67=>x"8900", 68=>x"8700", 69=>x"8100", 70=>x"8600",
---- 71=>x"8200", 72=>x"8600", 73=>x"8800", 74=>x"8700", 75=>x"8800", 76=>x"8700", 77=>x"8400",
---- 78=>x"8400", 79=>x"8300", 80=>x"8200", 81=>x"8400", 82=>x"8700", 83=>x"8900", 84=>x"8c00",
---- 85=>x"8700", 86=>x"8400", 87=>x"8300", 88=>x"8300", 89=>x"8300", 90=>x"8500", 91=>x"8600",
---- 92=>x"8800", 93=>x"8300", 94=>x"8400", 95=>x"8200", 96=>x"8400", 97=>x"8200", 98=>x"8200",
---- 99=>x"8200", 100=>x"8300", 101=>x"8500", 102=>x"8300", 103=>x"8200", 104=>x"7c00", 105=>x"8000",
---- 106=>x"8000", 107=>x"8200", 108=>x"8400", 109=>x"8300", 110=>x"8400", 111=>x"8200", 112=>x"7f00",
---- 113=>x"8200", 114=>x"8100", 115=>x"7e00", 116=>x"8200", 117=>x"8200", 118=>x"8200", 119=>x"8400",
---- 120=>x"7f00", 121=>x"8200", 122=>x"8400", 123=>x"8100", 124=>x"8000", 125=>x"8000", 126=>x"8000",
---- 127=>x"8300", 128=>x"7d00", 129=>x"7e00", 130=>x"8300", 131=>x"8000", 132=>x"8100", 133=>x"8100",
---- 134=>x"8000", 135=>x"7f00", 136=>x"7b00", 137=>x"7e00", 138=>x"8100", 139=>x"8000", 140=>x"8100",
---- 141=>x"8300", 142=>x"8100", 143=>x"8000", 144=>x"7c00", 145=>x"7c00", 146=>x"8200", 147=>x"8100",
---- 148=>x"7f00", 149=>x"8100", 150=>x"8400", 151=>x"8200", 152=>x"7d00", 153=>x"7d00", 154=>x"7d00",
---- 155=>x"7f00", 156=>x"8000", 157=>x"7e00", 158=>x"8100", 159=>x"8100", 160=>x"7a00", 161=>x"7900",
---- 162=>x"7d00", 163=>x"8000", 164=>x"7e00", 165=>x"7f00", 166=>x"8500", 167=>x"8100", 168=>x"7800",
---- 169=>x"7800", 170=>x"7c00", 171=>x"7d00", 172=>x"7d00", 173=>x"8000", 174=>x"8100", 175=>x"8100",
---- 176=>x"7500", 177=>x"7400", 178=>x"7900", 179=>x"7c00", 180=>x"7900", 181=>x"7900", 182=>x"7d00",
---- 183=>x"7f00", 184=>x"8b00", 185=>x"8300", 186=>x"7500", 187=>x"7300", 188=>x"7300", 189=>x"7500",
---- 190=>x"7700", 191=>x"7800", 192=>x"bd00", 193=>x"b100", 194=>x"a100", 195=>x"9900", 196=>x"8400",
---- 197=>x"7900", 198=>x"7200", 199=>x"7300", 200=>x"b200", 201=>x"b600", 202=>x"c300", 203=>x"c200",
---- 204=>x"ba00", 205=>x"aa00", 206=>x"9500", 207=>x"8400", 208=>x"b100", 209=>x"b700", 210=>x"b400",
---- 211=>x"ba00", 212=>x"ba00", 213=>x"c200", 214=>x"c500", 215=>x"b700", 216=>x"5000", 217=>x"b600",
---- 218=>x"b400", 219=>x"b600", 220=>x"b800", 221=>x"be00", 222=>x"bb00", 223=>x"c300", 224=>x"b200",
---- 225=>x"b400", 226=>x"b400", 227=>x"b400", 228=>x"b400", 229=>x"ba00", 230=>x"bf00", 231=>x"bd00",
---- 232=>x"ad00", 233=>x"b500", 234=>x"b700", 235=>x"ba00", 236=>x"bc00", 237=>x"b900", 238=>x"c000",
---- 239=>x"bf00", 240=>x"5200", 241=>x"b700", 242=>x"ba00", 243=>x"bb00", 244=>x"bb00", 245=>x"bd00",
---- 246=>x"bf00", 247=>x"4000", 248=>x"b700", 249=>x"b900", 250=>x"b800", 251=>x"bc00", 252=>x"4800",
---- 253=>x"b700", 254=>x"bf00", 255=>x"bc00", 256=>x"be00", 257=>x"ba00", 258=>x"b600", 259=>x"b700",
---- 260=>x"b700", 261=>x"bd00", 262=>x"c000", 263=>x"bb00", 264=>x"b300", 265=>x"b900", 266=>x"bb00",
---- 267=>x"b800", 268=>x"bb00", 269=>x"be00", 270=>x"bd00", 271=>x"b800", 272=>x"b500", 273=>x"b900",
---- 274=>x"bb00", 275=>x"b600", 276=>x"bd00", 277=>x"bb00", 278=>x"bb00", 279=>x"bf00", 280=>x"b000",
---- 281=>x"ba00", 282=>x"b400", 283=>x"b200", 284=>x"b800", 285=>x"bf00", 286=>x"be00", 287=>x"3f00",
---- 288=>x"b900", 289=>x"b500", 290=>x"b500", 291=>x"bc00", 292=>x"c000", 293=>x"bf00", 294=>x"bf00",
---- 295=>x"c400", 296=>x"b700", 297=>x"b700", 298=>x"bb00", 299=>x"bc00", 300=>x"c000", 301=>x"c100",
---- 302=>x"bf00", 303=>x"bd00", 304=>x"b800", 305=>x"b800", 306=>x"bc00", 307=>x"b900", 308=>x"ba00",
---- 309=>x"c000", 310=>x"c000", 311=>x"be00", 312=>x"bd00", 313=>x"be00", 314=>x"b300", 315=>x"bc00",
---- 316=>x"be00", 317=>x"b700", 318=>x"be00", 319=>x"be00", 320=>x"b600", 321=>x"ba00", 322=>x"bb00",
---- 323=>x"b700", 324=>x"b900", 325=>x"be00", 326=>x"be00", 327=>x"c000", 328=>x"bc00", 329=>x"bb00",
---- 330=>x"b400", 331=>x"bc00", 332=>x"be00", 333=>x"b800", 334=>x"b900", 335=>x"c100", 336=>x"bb00",
---- 337=>x"b800", 338=>x"3c00", 339=>x"c100", 340=>x"b800", 341=>x"bd00", 342=>x"bd00", 343=>x"b800",
---- 344=>x"4400", 345=>x"ba00", 346=>x"bb00", 347=>x"c000", 348=>x"c200", 349=>x"ac00", 350=>x"a300",
---- 351=>x"a800", 352=>x"af00", 353=>x"b700", 354=>x"bc00", 355=>x"b300", 356=>x"aa00", 357=>x"9d00",
---- 358=>x"ac00", 359=>x"c200", 360=>x"b600", 361=>x"bd00", 362=>x"a000", 363=>x"9700", 364=>x"a400",
---- 365=>x"b800", 366=>x"ce00", 367=>x"d000", 368=>x"a700", 369=>x"9d00", 370=>x"9900", 371=>x"b700",
---- 372=>x"ca00", 373=>x"cd00", 374=>x"cb00", 375=>x"d000", 376=>x"8d00", 377=>x"9d00", 378=>x"bf00",
---- 379=>x"d200", 380=>x"cf00", 381=>x"d000", 382=>x"cb00", 383=>x"c600", 384=>x"aa00", 385=>x"c700",
---- 386=>x"cb00", 387=>x"cb00", 388=>x"ca00", 389=>x"ca00", 390=>x"cb00", 391=>x"c800", 392=>x"c400",
---- 393=>x"c400", 394=>x"cb00", 395=>x"c900", 396=>x"c300", 397=>x"cb00", 398=>x"d000", 399=>x"d100",
---- 400=>x"c000", 401=>x"c200", 402=>x"c100", 403=>x"cc00", 404=>x"ca00", 405=>x"c500", 406=>x"cf00",
---- 407=>x"ce00", 408=>x"bf00", 409=>x"c200", 410=>x"c700", 411=>x"c000", 412=>x"c600", 413=>x"c300",
---- 414=>x"c300", 415=>x"c400", 416=>x"c800", 417=>x"be00", 418=>x"c300", 419=>x"c200", 420=>x"bb00",
---- 421=>x"c100", 422=>x"c100", 423=>x"be00", 424=>x"c100", 425=>x"c200", 426=>x"bb00", 427=>x"c300",
---- 428=>x"c100", 429=>x"b800", 430=>x"c400", 431=>x"c300", 432=>x"be00", 433=>x"bf00", 434=>x"c300",
---- 435=>x"b900", 436=>x"c000", 437=>x"c200", 438=>x"b800", 439=>x"b800", 440=>x"c000", 441=>x"c200",
---- 442=>x"c200", 443=>x"c100", 444=>x"b100", 445=>x"ba00", 446=>x"be00", 447=>x"c200", 448=>x"c100",
---- 449=>x"be00", 450=>x"b500", 451=>x"ac00", 452=>x"b700", 453=>x"c400", 454=>x"ca00", 455=>x"c200",
---- 456=>x"af00", 457=>x"a700", 458=>x"b200", 459=>x"bc00", 460=>x"c200", 461=>x"c300", 462=>x"c500",
---- 463=>x"c800", 464=>x"a800", 465=>x"b800", 466=>x"ba00", 467=>x"bf00", 468=>x"bc00", 469=>x"c200",
---- 470=>x"c200", 471=>x"3b00", 472=>x"c100", 473=>x"be00", 474=>x"bc00", 475=>x"b700", 476=>x"bd00",
---- 477=>x"c300", 478=>x"c600", 479=>x"c100", 480=>x"bd00", 481=>x"b600", 482=>x"b900", 483=>x"bc00",
---- 484=>x"b700", 485=>x"c000", 486=>x"c400", 487=>x"bf00", 488=>x"b600", 489=>x"bc00", 490=>x"bf00",
---- 491=>x"bc00", 492=>x"bf00", 493=>x"bf00", 494=>x"c200", 495=>x"bb00", 496=>x"bc00", 497=>x"bf00",
---- 498=>x"c200", 499=>x"bd00", 500=>x"b900", 501=>x"bf00", 502=>x"ba00", 503=>x"c100", 504=>x"b800",
---- 505=>x"c500", 506=>x"bc00", 507=>x"c300", 508=>x"ba00", 509=>x"b600", 510=>x"4700", 511=>x"b900",
---- 512=>x"ba00", 513=>x"b700", 514=>x"bd00", 515=>x"b700", 516=>x"c100", 517=>x"ba00", 518=>x"bc00",
---- 519=>x"b700", 520=>x"b800", 521=>x"b800", 522=>x"b500", 523=>x"b800", 524=>x"b600", 525=>x"bd00",
---- 526=>x"ba00", 527=>x"b200", 528=>x"b900", 529=>x"b600", 530=>x"b500", 531=>x"b300", 532=>x"bb00",
---- 533=>x"b400", 534=>x"aa00", 535=>x"a300", 536=>x"b900", 537=>x"b300", 538=>x"b400", 539=>x"b700",
---- 540=>x"b100", 541=>x"a100", 542=>x"a600", 543=>x"b700", 544=>x"b300", 545=>x"ba00", 546=>x"ba00",
---- 547=>x"ab00", 548=>x"9c00", 549=>x"a400", 550=>x"be00", 551=>x"bd00", 552=>x"b300", 553=>x"b100",
---- 554=>x"ad00", 555=>x"a100", 556=>x"ae00", 557=>x"b600", 558=>x"b200", 559=>x"ba00", 560=>x"a800",
---- 561=>x"9b00", 562=>x"9f00", 563=>x"b800", 564=>x"b600", 565=>x"b100", 566=>x"af00", 567=>x"ad00",
---- 568=>x"9900", 569=>x"9c00", 570=>x"b400", 571=>x"b500", 572=>x"ae00", 573=>x"ac00", 574=>x"ad00",
---- 575=>x"b000", 576=>x"a800", 577=>x"b200", 578=>x"ad00", 579=>x"af00", 580=>x"b200", 581=>x"b200",
---- 582=>x"b200", 583=>x"ae00", 584=>x"b100", 585=>x"b300", 586=>x"ae00", 587=>x"a600", 588=>x"af00",
---- 589=>x"b500", 590=>x"b300", 591=>x"ad00", 592=>x"b100", 593=>x"a800", 594=>x"ae00", 595=>x"b000",
---- 596=>x"a800", 597=>x"ab00", 598=>x"b200", 599=>x"5100", 600=>x"b000", 601=>x"a800", 602=>x"a800",
---- 603=>x"af00", 604=>x"b400", 605=>x"5300", 606=>x"a500", 607=>x"b000", 608=>x"a100", 609=>x"b000",
---- 610=>x"ae00", 611=>x"ac00", 612=>x"b100", 613=>x"b800", 614=>x"ae00", 615=>x"a700", 616=>x"a100",
---- 617=>x"a500", 618=>x"4d00", 619=>x"b100", 620=>x"ad00", 621=>x"b000", 622=>x"b600", 623=>x"ae00",
---- 624=>x"a800", 625=>x"a300", 626=>x"a100", 627=>x"aa00", 628=>x"b100", 629=>x"aa00", 630=>x"a500",
---- 631=>x"a800", 632=>x"a900", 633=>x"ac00", 634=>x"a700", 635=>x"9f00", 636=>x"a400", 637=>x"ae00",
---- 638=>x"a400", 639=>x"9d00", 640=>x"ac00", 641=>x"a900", 642=>x"ab00", 643=>x"a200", 644=>x"9c00",
---- 645=>x"9d00", 646=>x"b100", 647=>x"a800", 648=>x"a400", 649=>x"9f00", 650=>x"9f00", 651=>x"a400",
---- 652=>x"a500", 653=>x"9f00", 654=>x"9f00", 655=>x"ac00", 656=>x"9b00", 657=>x"6000", 658=>x"a000",
---- 659=>x"a200", 660=>x"a400", 661=>x"ae00", 662=>x"a600", 663=>x"9b00", 664=>x"9700", 665=>x"a600",
---- 666=>x"a700", 667=>x"aa00", 668=>x"aa00", 669=>x"a500", 670=>x"9d00", 671=>x"9000", 672=>x"8300",
---- 673=>x"8300", 674=>x"8700", 675=>x"8400", 676=>x"8900", 677=>x"9300", 678=>x"9c00", 679=>x"9e00",
---- 680=>x"8400", 681=>x"8a00", 682=>x"8100", 683=>x"6700", 684=>x"4a00", 685=>x"8500", 686=>x"ae00",
---- 687=>x"9e00", 688=>x"8c00", 689=>x"9600", 690=>x"9800", 691=>x"9100", 692=>x"6100", 693=>x"6a00",
---- 694=>x"9c00", 695=>x"9c00", 696=>x"8d00", 697=>x"a200", 698=>x"a600", 699=>x"a200", 700=>x"9000",
---- 701=>x"7100", 702=>x"6c00", 703=>x"6c00", 704=>x"9900", 705=>x"ab00", 706=>x"a500", 707=>x"a700",
---- 708=>x"9600", 709=>x"7f00", 710=>x"8200", 711=>x"7700", 712=>x"9000", 713=>x"9c00", 714=>x"a400",
---- 715=>x"9e00", 716=>x"8500", 717=>x"8300", 718=>x"8300", 719=>x"7a00", 720=>x"8200", 721=>x"8a00",
---- 722=>x"8d00", 723=>x"8a00", 724=>x"8900", 725=>x"7900", 726=>x"5900", 727=>x"4600", 728=>x"6b00",
---- 729=>x"5800", 730=>x"7400", 731=>x"8400", 732=>x"5f00", 733=>x"4e00", 734=>x"5100", 735=>x"3d00",
---- 736=>x"4b00", 737=>x"5000", 738=>x"7300", 739=>x"6400", 740=>x"6400", 741=>x"5500", 742=>x"4c00",
---- 743=>x"4800", 744=>x"4200", 745=>x"5e00", 746=>x"6400", 747=>x"7900", 748=>x"6d00", 749=>x"6a00",
---- 750=>x"6300", 751=>x"7b00", 752=>x"5b00", 753=>x"6800", 754=>x"7300", 755=>x"7500", 756=>x"5a00",
---- 757=>x"4d00", 758=>x"4e00", 759=>x"6500", 760=>x"7b00", 761=>x"6800", 762=>x"7400", 763=>x"5700",
---- 764=>x"3b00", 765=>x"3000", 766=>x"3800", 767=>x"6000", 768=>x"7c00", 769=>x"7400", 770=>x"6100",
---- 771=>x"3400", 772=>x"2a00", 773=>x"2800", 774=>x"4f00", 775=>x"7600", 776=>x"7000", 777=>x"5f00",
---- 778=>x"3600", 779=>x"3200", 780=>x"2c00", 781=>x"4800", 782=>x"8200", 783=>x"4e00", 784=>x"4c00",
---- 785=>x"4400", 786=>x"2b00", 787=>x"3200", 788=>x"5000", 789=>x"8300", 790=>x"6b00", 791=>x"4c00",
---- 792=>x"3a00", 793=>x"3700", 794=>x"3100", 795=>x"4600", 796=>x"7600", 797=>x"5800", 798=>x"6200",
---- 799=>x"7900", 800=>x"3400", 801=>x"3500", 802=>x"3700", 803=>x"6a00", 804=>x"5300", 805=>x"4d00",
---- 806=>x"7000", 807=>x"5e00", 808=>x"2e00", 809=>x"3800", 810=>x"3f00", 811=>x"5100", 812=>x"3d00",
---- 813=>x"4000", 814=>x"6100", 815=>x"4400", 816=>x"3b00", 817=>x"3d00", 818=>x"3c00", 819=>x"3600",
---- 820=>x"2a00", 821=>x"4200", 822=>x"6d00", 823=>x"2e00", 824=>x"3e00", 825=>x"2f00", 826=>x"3000",
---- 827=>x"3400", 828=>x"2500", 829=>x"4900", 830=>x"6900", 831=>x"2800", 832=>x"4e00", 833=>x"5500",
---- 834=>x"4f00", 835=>x"5400", 836=>x"3c00", 837=>x"5b00", 838=>x"6100", 839=>x"3b00", 840=>x"3d00",
---- 841=>x"4400", 842=>x"4a00", 843=>x"4300", 844=>x"3e00", 845=>x"5700", 846=>x"5200", 847=>x"4400",
---- 848=>x"3100", 849=>x"2e00", 850=>x"2f00", 851=>x"2800", 852=>x"2300", 853=>x"c100", 854=>x"4400",
---- 855=>x"4e00", 856=>x"3600", 857=>x"3100", 858=>x"2c00", 859=>x"2e00", 860=>x"2700", 861=>x"3d00",
---- 862=>x"6100", 863=>x"7000", 864=>x"2f00", 865=>x"2f00", 866=>x"2600", 867=>x"2500", 868=>x"2d00",
---- 869=>x"5400", 870=>x"7f00", 871=>x"a200", 872=>x"2800", 873=>x"2400", 874=>x"2300", 875=>x"2500",
---- 876=>x"5c00", 877=>x"7c00", 878=>x"6d00", 879=>x"5100", 880=>x"2300", 881=>x"2400", 882=>x"2100",
---- 883=>x"a600", 884=>x"9c00", 885=>x"7500", 886=>x"5700", 887=>x"7b00", 888=>x"2100", 889=>x"e200",
---- 890=>x"5400", 891=>x"9d00", 892=>x"8b00", 893=>x"6600", 894=>x"7e00", 895=>x"b500", 896=>x"1900",
---- 897=>x"4200", 898=>x"a000", 899=>x"8e00", 900=>x"6700", 901=>x"8600", 902=>x"b700", 903=>x"b200",
---- 904=>x"3b00", 905=>x"9500", 906=>x"9400", 907=>x"6900", 908=>x"8100", 909=>x"b200", 910=>x"b100",
---- 911=>x"a600", 912=>x"8a00", 913=>x"9b00", 914=>x"7600", 915=>x"7e00", 916=>x"4d00", 917=>x"b100",
---- 918=>x"af00", 919=>x"af00", 920=>x"9a00", 921=>x"7700", 922=>x"7800", 923=>x"af00", 924=>x"b500",
---- 925=>x"ac00", 926=>x"b900", 927=>x"b400", 928=>x"7800", 929=>x"7300", 930=>x"a000", 931=>x"b400",
---- 932=>x"a800", 933=>x"b000", 934=>x"bb00", 935=>x"bc00", 936=>x"7500", 937=>x"9800", 938=>x"ac00",
---- 939=>x"5c00", 940=>x"ae00", 941=>x"af00", 942=>x"bc00", 943=>x"bd00", 944=>x"8e00", 945=>x"b000",
---- 946=>x"9f00", 947=>x"a200", 948=>x"a700", 949=>x"b300", 950=>x"bc00", 951=>x"b900", 952=>x"b300",
---- 953=>x"a100", 954=>x"a000", 955=>x"a000", 956=>x"a200", 957=>x"5400", 958=>x"ba00", 959=>x"bc00",
---- 960=>x"a500", 961=>x"a100", 962=>x"a400", 963=>x"a100", 964=>x"9f00", 965=>x"a600", 966=>x"ba00",
---- 967=>x"c000", 968=>x"a400", 969=>x"ac00", 970=>x"ac00", 971=>x"a300", 972=>x"9d00", 973=>x"a800",
---- 974=>x"bc00", 975=>x"bf00", 976=>x"ad00", 977=>x"b500", 978=>x"af00", 979=>x"9e00", 980=>x"9800",
---- 981=>x"5900", 982=>x"bb00", 983=>x"c100", 984=>x"b500", 985=>x"c000", 986=>x"ac00", 987=>x"6600",
---- 988=>x"9800", 989=>x"ac00", 990=>x"be00", 991=>x"c100", 992=>x"bf00", 993=>x"c100", 994=>x"a500",
---- 995=>x"9700", 996=>x"a000", 997=>x"b600", 998=>x"bc00", 999=>x"c000", 1000=>x"c600", 1001=>x"b600",
---- 1002=>x"9800", 1003=>x"9b00", 1004=>x"ac00", 1005=>x"ba00", 1006=>x"c100", 1007=>x"c800", 1008=>x"c400",
---- 1009=>x"a800", 1010=>x"9700", 1011=>x"a500", 1012=>x"b800", 1013=>x"c500", 1014=>x"c800", 1015=>x"9a00",
---- 1016=>x"ba00", 1017=>x"a500", 1018=>x"a200", 1019=>x"b000", 1020=>x"c400", 1021=>x"c800", 1022=>x"8800",
---- 1023=>x"6200", 1024=>x"b800", 1025=>x"ac00", 1026=>x"ae00", 1027=>x"c300", 1028=>x"c400", 1029=>x"7400",
---- 1030=>x"5200", 1031=>x"6100", 1032=>x"b900", 1033=>x"b400", 1034=>x"c100", 1035=>x"c000", 1036=>x"6700",
---- 1037=>x"4700", 1038=>x"5100", 1039=>x"4b00", 1040=>x"ba00", 1041=>x"be00", 1042=>x"c100", 1043=>x"6600",
---- 1044=>x"3900", 1045=>x"4600", 1046=>x"3a00", 1047=>x"c900", 1048=>x"c200", 1049=>x"c200", 1050=>x"6800",
---- 1051=>x"4400", 1052=>x"4600", 1053=>x"3b00", 1054=>x"3000", 1055=>x"3000", 1056=>x"c300", 1057=>x"7300",
---- 1058=>x"4900", 1059=>x"5400", 1060=>x"4500", 1061=>x"3300", 1062=>x"2900", 1063=>x"2f00", 1064=>x"8200",
---- 1065=>x"5300", 1066=>x"5b00", 1067=>x"4800", 1068=>x"3500", 1069=>x"3000", 1070=>x"2c00", 1071=>x"3800",
---- 1072=>x"5e00", 1073=>x"7100", 1074=>x"6900", 1075=>x"5700", 1076=>x"4a00", 1077=>x"3a00", 1078=>x"2c00",
---- 1079=>x"4000", 1080=>x"7200", 1081=>x"7d00", 1082=>x"7d00", 1083=>x"7400", 1084=>x"7100", 1085=>x"5c00",
---- 1086=>x"3400", 1087=>x"3400", 1088=>x"7700", 1089=>x"7c00", 1090=>x"8500", 1091=>x"8900", 1092=>x"8600",
---- 1093=>x"7600", 1094=>x"5100", 1095=>x"4200", 1096=>x"7e00", 1097=>x"7d00", 1098=>x"8500", 1099=>x"9200",
---- 1100=>x"8d00", 1101=>x"8a00", 1102=>x"7a00", 1103=>x"6b00", 1104=>x"8600", 1105=>x"8300", 1106=>x"8700",
---- 1107=>x"9100", 1108=>x"9000", 1109=>x"9000", 1110=>x"8d00", 1111=>x"7b00", 1112=>x"8b00", 1113=>x"8b00",
---- 1114=>x"8c00", 1115=>x"9000", 1116=>x"9000", 1117=>x"9000", 1118=>x"9200", 1119=>x"8d00", 1120=>x"9100",
---- 1121=>x"8f00", 1122=>x"9000", 1123=>x"9400", 1124=>x"9500", 1125=>x"9100", 1126=>x"8d00", 1127=>x"9000",
---- 1128=>x"9300", 1129=>x"6800", 1130=>x"9900", 1131=>x"9600", 1132=>x"9700", 1133=>x"9700", 1134=>x"9700",
---- 1135=>x"9400", 1136=>x"9600", 1137=>x"9900", 1138=>x"9900", 1139=>x"9700", 1140=>x"9d00", 1141=>x"a000",
---- 1142=>x"a200", 1143=>x"a000", 1144=>x"9400", 1145=>x"9600", 1146=>x"9a00", 1147=>x"9d00", 1148=>x"a300",
---- 1149=>x"a700", 1150=>x"a400", 1151=>x"a300", 1152=>x"9100", 1153=>x"9600", 1154=>x"9a00", 1155=>x"9e00",
---- 1156=>x"a100", 1157=>x"aa00", 1158=>x"a400", 1159=>x"a400", 1160=>x"8f00", 1161=>x"9700", 1162=>x"9900",
---- 1163=>x"9d00", 1164=>x"a100", 1165=>x"a600", 1166=>x"aa00", 1167=>x"a700", 1168=>x"9000", 1169=>x"9600",
---- 1170=>x"9700", 1171=>x"9b00", 1172=>x"a100", 1173=>x"a400", 1174=>x"ad00", 1175=>x"ab00", 1176=>x"9100",
---- 1177=>x"9400", 1178=>x"9600", 1179=>x"9b00", 1180=>x"9f00", 1181=>x"a600", 1182=>x"a800", 1183=>x"ab00",
---- 1184=>x"8f00", 1185=>x"9200", 1186=>x"9800", 1187=>x"9900", 1188=>x"9d00", 1189=>x"a200", 1190=>x"a900",
---- 1191=>x"ae00", 1192=>x"8800", 1193=>x"9100", 1194=>x"9500", 1195=>x"9300", 1196=>x"9900", 1197=>x"a000",
---- 1198=>x"a800", 1199=>x"ab00", 1200=>x"8a00", 1201=>x"9100", 1202=>x"9000", 1203=>x"9200", 1204=>x"6700",
---- 1205=>x"9c00", 1206=>x"9e00", 1207=>x"a300", 1208=>x"8b00", 1209=>x"8f00", 1210=>x"9300", 1211=>x"9600",
---- 1212=>x"9900", 1213=>x"9800", 1214=>x"9b00", 1215=>x"a100", 1216=>x"8c00", 1217=>x"8e00", 1218=>x"9300",
---- 1219=>x"9700", 1220=>x"9800", 1221=>x"9b00", 1222=>x"9d00", 1223=>x"a000", 1224=>x"8800", 1225=>x"8c00",
---- 1226=>x"9000", 1227=>x"9400", 1228=>x"9700", 1229=>x"9b00", 1230=>x"9e00", 1231=>x"a000", 1232=>x"8700",
---- 1233=>x"8b00", 1234=>x"8d00", 1235=>x"9300", 1236=>x"9800", 1237=>x"9c00", 1238=>x"9b00", 1239=>x"9f00",
---- 1240=>x"8a00", 1241=>x"8800", 1242=>x"8b00", 1243=>x"9500", 1244=>x"6d00", 1245=>x"9800", 1246=>x"9800",
---- 1247=>x"9d00", 1248=>x"8500", 1249=>x"8a00", 1250=>x"8f00", 1251=>x"8f00", 1252=>x"9200", 1253=>x"9600",
---- 1254=>x"9600", 1255=>x"9800", 1256=>x"8700", 1257=>x"8500", 1258=>x"8a00", 1259=>x"8c00", 1260=>x"9300",
---- 1261=>x"9400", 1262=>x"9600", 1263=>x"9700", 1264=>x"8700", 1265=>x"8a00", 1266=>x"8b00", 1267=>x"8f00",
---- 1268=>x"9200", 1269=>x"9100", 1270=>x"9a00", 1271=>x"9800", 1272=>x"8400", 1273=>x"8800", 1274=>x"8b00",
---- 1275=>x"8f00", 1276=>x"8f00", 1277=>x"8f00", 1278=>x"6c00", 1279=>x"9600", 1280=>x"8400", 1281=>x"8500",
---- 1282=>x"8d00", 1283=>x"8b00", 1284=>x"8f00", 1285=>x"9000", 1286=>x"9200", 1287=>x"9600", 1288=>x"8400",
---- 1289=>x"8900", 1290=>x"8b00", 1291=>x"8a00", 1292=>x"8f00", 1293=>x"8f00", 1294=>x"9600", 1295=>x"9600",
---- 1296=>x"8200", 1297=>x"8700", 1298=>x"8800", 1299=>x"8b00", 1300=>x"6e00", 1301=>x"9100", 1302=>x"9300",
---- 1303=>x"9700", 1304=>x"8300", 1305=>x"8700", 1306=>x"8800", 1307=>x"8d00", 1308=>x"9100", 1309=>x"9100",
---- 1310=>x"9100", 1311=>x"9400", 1312=>x"8200", 1313=>x"8500", 1314=>x"8800", 1315=>x"8900", 1316=>x"8d00",
---- 1317=>x"9300", 1318=>x"9100", 1319=>x"9400", 1320=>x"7f00", 1321=>x"8400", 1322=>x"8600", 1323=>x"8900",
---- 1324=>x"8a00", 1325=>x"8f00", 1326=>x"9000", 1327=>x"9000", 1328=>x"8200", 1329=>x"8200", 1330=>x"8600",
---- 1331=>x"8800", 1332=>x"8900", 1333=>x"8e00", 1334=>x"9100", 1335=>x"8f00", 1336=>x"8200", 1337=>x"8600",
---- 1338=>x"8b00", 1339=>x"8b00", 1340=>x"8d00", 1341=>x"8d00", 1342=>x"8b00", 1343=>x"8d00", 1344=>x"8200",
---- 1345=>x"8500", 1346=>x"8800", 1347=>x"8a00", 1348=>x"8d00", 1349=>x"8d00", 1350=>x"8d00", 1351=>x"8a00",
---- 1352=>x"8100", 1353=>x"8400", 1354=>x"8900", 1355=>x"8800", 1356=>x"8c00", 1357=>x"8b00", 1358=>x"8d00",
---- 1359=>x"8b00", 1360=>x"8000", 1361=>x"8400", 1362=>x"8800", 1363=>x"8700", 1364=>x"8b00", 1365=>x"8e00",
---- 1366=>x"8c00", 1367=>x"8900", 1368=>x"8100", 1369=>x"8600", 1370=>x"8900", 1371=>x"8900", 1372=>x"7500",
---- 1373=>x"8f00", 1374=>x"8b00", 1375=>x"8e00", 1376=>x"8300", 1377=>x"8300", 1378=>x"8800", 1379=>x"8900",
---- 1380=>x"8b00", 1381=>x"8a00", 1382=>x"8d00", 1383=>x"8a00", 1384=>x"7f00", 1385=>x"8300", 1386=>x"8600",
---- 1387=>x"8700", 1388=>x"8600", 1389=>x"8a00", 1390=>x"8d00", 1391=>x"8d00", 1392=>x"7c00", 1393=>x"8100",
---- 1394=>x"8300", 1395=>x"8500", 1396=>x"8600", 1397=>x"8500", 1398=>x"8b00", 1399=>x"9100", 1400=>x"7d00",
---- 1401=>x"7f00", 1402=>x"8100", 1403=>x"8200", 1404=>x"8700", 1405=>x"8a00", 1406=>x"8b00", 1407=>x"8d00",
---- 1408=>x"7d00", 1409=>x"7d00", 1410=>x"8100", 1411=>x"8300", 1412=>x"8700", 1413=>x"8b00", 1414=>x"8800",
---- 1415=>x"8b00", 1416=>x"8600", 1417=>x"7e00", 1418=>x"7f00", 1419=>x"8000", 1420=>x"8400", 1421=>x"8800",
---- 1422=>x"8800", 1423=>x"8700", 1424=>x"7800", 1425=>x"7c00", 1426=>x"7d00", 1427=>x"7f00", 1428=>x"8100",
---- 1429=>x"8200", 1430=>x"8600", 1431=>x"8800", 1432=>x"7700", 1433=>x"7a00", 1434=>x"7a00", 1435=>x"7b00",
---- 1436=>x"7f00", 1437=>x"8200", 1438=>x"7e00", 1439=>x"8500", 1440=>x"7300", 1441=>x"7700", 1442=>x"7800",
---- 1443=>x"7c00", 1444=>x"7d00", 1445=>x"8100", 1446=>x"8000", 1447=>x"8200", 1448=>x"7400", 1449=>x"7600",
---- 1450=>x"7800", 1451=>x"7c00", 1452=>x"7c00", 1453=>x"8200", 1454=>x"8400", 1455=>x"8400", 1456=>x"6f00",
---- 1457=>x"7300", 1458=>x"7700", 1459=>x"7700", 1460=>x"7800", 1461=>x"7f00", 1462=>x"8300", 1463=>x"8100",
---- 1464=>x"6b00", 1465=>x"6900", 1466=>x"7200", 1467=>x"7400", 1468=>x"7800", 1469=>x"7c00", 1470=>x"8100",
---- 1471=>x"8100", 1472=>x"6900", 1473=>x"6c00", 1474=>x"6e00", 1475=>x"7500", 1476=>x"7a00", 1477=>x"7e00",
---- 1478=>x"8000", 1479=>x"7f00", 1480=>x"6800", 1481=>x"6a00", 1482=>x"6f00", 1483=>x"7100", 1484=>x"7700",
---- 1485=>x"7e00", 1486=>x"7e00", 1487=>x"7f00", 1488=>x"6300", 1489=>x"6600", 1490=>x"6b00", 1491=>x"6e00",
---- 1492=>x"7100", 1493=>x"7c00", 1494=>x"7f00", 1495=>x"7f00", 1496=>x"5600", 1497=>x"5c00", 1498=>x"6600",
---- 1499=>x"6800", 1500=>x"6f00", 1501=>x"7600", 1502=>x"7c00", 1503=>x"8300", 1504=>x"4800", 1505=>x"5300",
---- 1506=>x"5e00", 1507=>x"5e00", 1508=>x"6800", 1509=>x"7000", 1510=>x"7600", 1511=>x"7f00", 1512=>x"3500",
---- 1513=>x"4300", 1514=>x"5100", 1515=>x"5800", 1516=>x"5c00", 1517=>x"9600", 1518=>x"7500", 1519=>x"7800",
---- 1520=>x"2c00", 1521=>x"3600", 1522=>x"3f00", 1523=>x"4c00", 1524=>x"5200", 1525=>x"6000", 1526=>x"6f00",
---- 1527=>x"7600", 1528=>x"3000", 1529=>x"2c00", 1530=>x"3200", 1531=>x"3a00", 1532=>x"4a00", 1533=>x"5400",
---- 1534=>x"6000", 1535=>x"6800", 1536=>x"3700", 1537=>x"3600", 1538=>x"3100", 1539=>x"3800", 1540=>x"3b00",
---- 1541=>x"4000", 1542=>x"4300", 1543=>x"4500", 1544=>x"3f00", 1545=>x"3c00", 1546=>x"3d00", 1547=>x"4500",
---- 1548=>x"4500", 1549=>x"4600", 1550=>x"4800", 1551=>x"4d00", 1552=>x"4900", 1553=>x"4b00", 1554=>x"5400",
---- 1555=>x"6600", 1556=>x"6c00", 1557=>x"6d00", 1558=>x"7500", 1559=>x"7c00", 1560=>x"5400", 1561=>x"5a00",
---- 1562=>x"6a00", 1563=>x"6e00", 1564=>x"7700", 1565=>x"7b00", 1566=>x"8200", 1567=>x"8300", 1568=>x"5400",
---- 1569=>x"6300", 1570=>x"6f00", 1571=>x"8900", 1572=>x"8000", 1573=>x"8200", 1574=>x"8100", 1575=>x"7e00",
---- 1576=>x"5700", 1577=>x"6600", 1578=>x"7500", 1579=>x"7b00", 1580=>x"7f00", 1581=>x"8000", 1582=>x"7e00",
---- 1583=>x"7c00", 1584=>x"5b00", 1585=>x"6b00", 1586=>x"7300", 1587=>x"7900", 1588=>x"7c00", 1589=>x"7d00",
---- 1590=>x"7e00", 1591=>x"7c00", 1592=>x"5900", 1593=>x"6b00", 1594=>x"7900", 1595=>x"7900", 1596=>x"7500",
---- 1597=>x"7c00", 1598=>x"7e00", 1599=>x"7d00", 1600=>x"5a00", 1601=>x"6700", 1602=>x"7300", 1603=>x"7400",
---- 1604=>x"7a00", 1605=>x"7c00", 1606=>x"7a00", 1607=>x"7b00", 1608=>x"5e00", 1609=>x"6700", 1610=>x"6f00",
---- 1611=>x"7000", 1612=>x"7200", 1613=>x"7a00", 1614=>x"7b00", 1615=>x"7c00", 1616=>x"5900", 1617=>x"6500",
---- 1618=>x"7100", 1619=>x"7400", 1620=>x"7400", 1621=>x"7700", 1622=>x"7b00", 1623=>x"7e00", 1624=>x"5a00",
---- 1625=>x"6500", 1626=>x"7100", 1627=>x"7500", 1628=>x"8800", 1629=>x"7600", 1630=>x"7b00", 1631=>x"8100",
---- 1632=>x"5500", 1633=>x"6800", 1634=>x"7100", 1635=>x"7400", 1636=>x"7800", 1637=>x"7d00", 1638=>x"7e00",
---- 1639=>x"7e00", 1640=>x"5300", 1641=>x"6b00", 1642=>x"7400", 1643=>x"7200", 1644=>x"7900", 1645=>x"8300",
---- 1646=>x"7e00", 1647=>x"7200", 1648=>x"5200", 1649=>x"6e00", 1650=>x"7900", 1651=>x"7800", 1652=>x"7700",
---- 1653=>x"7c00", 1654=>x"7100", 1655=>x"6f00", 1656=>x"5200", 1657=>x"7000", 1658=>x"7b00", 1659=>x"7b00",
---- 1660=>x"7300", 1661=>x"7000", 1662=>x"7700", 1663=>x"8100", 1664=>x"5200", 1665=>x"6800", 1666=>x"7b00",
---- 1667=>x"7100", 1668=>x"6c00", 1669=>x"7900", 1670=>x"8800", 1671=>x"8300", 1672=>x"5200", 1673=>x"6200",
---- 1674=>x"6f00", 1675=>x"6c00", 1676=>x"7a00", 1677=>x"8500", 1678=>x"8a00", 1679=>x"8200", 1680=>x"4d00",
---- 1681=>x"6000", 1682=>x"6d00", 1683=>x"7900", 1684=>x"7c00", 1685=>x"8300", 1686=>x"8700", 1687=>x"8300",
---- 1688=>x"4a00", 1689=>x"6500", 1690=>x"7300", 1691=>x"7600", 1692=>x"7f00", 1693=>x"8500", 1694=>x"8500",
---- 1695=>x"8300", 1696=>x"4f00", 1697=>x"6600", 1698=>x"7200", 1699=>x"7600", 1700=>x"8000", 1701=>x"8300",
---- 1702=>x"8000", 1703=>x"8000", 1704=>x"5000", 1705=>x"6600", 1706=>x"7700", 1707=>x"7900", 1708=>x"8000",
---- 1709=>x"8200", 1710=>x"7e00", 1711=>x"7d00", 1712=>x"5300", 1713=>x"6000", 1714=>x"7200", 1715=>x"7c00",
---- 1716=>x"8500", 1717=>x"8400", 1718=>x"8100", 1719=>x"8100", 1720=>x"5800", 1721=>x"6300", 1722=>x"7200",
---- 1723=>x"8000", 1724=>x"8300", 1725=>x"8000", 1726=>x"8000", 1727=>x"8200", 1728=>x"5800", 1729=>x"6700",
---- 1730=>x"7200", 1731=>x"8000", 1732=>x"8400", 1733=>x"8300", 1734=>x"8400", 1735=>x"8600", 1736=>x"5b00",
---- 1737=>x"6600", 1738=>x"7300", 1739=>x"8000", 1740=>x"8400", 1741=>x"8500", 1742=>x"8800", 1743=>x"8600",
---- 1744=>x"5d00", 1745=>x"6800", 1746=>x"7700", 1747=>x"7d00", 1748=>x"8200", 1749=>x"8100", 1750=>x"8700",
---- 1751=>x"8a00", 1752=>x"5e00", 1753=>x"6700", 1754=>x"7900", 1755=>x"7c00", 1756=>x"7f00", 1757=>x"8400",
---- 1758=>x"8500", 1759=>x"8800", 1760=>x"5e00", 1761=>x"6700", 1762=>x"7a00", 1763=>x"8400", 1764=>x"8200",
---- 1765=>x"8500", 1766=>x"8300", 1767=>x"8500", 1768=>x"6300", 1769=>x"6e00", 1770=>x"7b00", 1771=>x"7f00",
---- 1772=>x"8400", 1773=>x"8500", 1774=>x"8300", 1775=>x"8700", 1776=>x"6500", 1777=>x"7000", 1778=>x"7e00",
---- 1779=>x"7e00", 1780=>x"8500", 1781=>x"8600", 1782=>x"8600", 1783=>x"8400", 1784=>x"6400", 1785=>x"7300",
---- 1786=>x"8500", 1787=>x"8200", 1788=>x"8400", 1789=>x"8700", 1790=>x"8600", 1791=>x"8700", 1792=>x"6400",
---- 1793=>x"7b00", 1794=>x"8700", 1795=>x"8300", 1796=>x"8600", 1797=>x"8500", 1798=>x"8a00", 1799=>x"8a00",
---- 1800=>x"6c00", 1801=>x"8100", 1802=>x"8400", 1803=>x"8300", 1804=>x"7800", 1805=>x"7500", 1806=>x"8a00",
---- 1807=>x"8a00", 1808=>x"7100", 1809=>x"8100", 1810=>x"8300", 1811=>x"8400", 1812=>x"8a00", 1813=>x"8c00",
---- 1814=>x"8900", 1815=>x"8c00", 1816=>x"7800", 1817=>x"8200", 1818=>x"8600", 1819=>x"8800", 1820=>x"8c00",
---- 1821=>x"8d00", 1822=>x"8c00", 1823=>x"8b00", 1824=>x"7d00", 1825=>x"8500", 1826=>x"8700", 1827=>x"8900",
---- 1828=>x"8900", 1829=>x"8e00", 1830=>x"8e00", 1831=>x"8a00", 1832=>x"8200", 1833=>x"8500", 1834=>x"8700",
---- 1835=>x"8800", 1836=>x"8c00", 1837=>x"8800", 1838=>x"8c00", 1839=>x"8e00", 1840=>x"8200", 1841=>x"8800",
---- 1842=>x"8700", 1843=>x"8800", 1844=>x"8b00", 1845=>x"8a00", 1846=>x"8a00", 1847=>x"8b00", 1848=>x"8600",
---- 1849=>x"8600", 1850=>x"8600", 1851=>x"8700", 1852=>x"8a00", 1853=>x"8c00", 1854=>x"8b00", 1855=>x"8e00",
---- 1856=>x"8600", 1857=>x"8400", 1858=>x"8700", 1859=>x"8900", 1860=>x"8b00", 1861=>x"8d00", 1862=>x"8f00",
---- 1863=>x"8f00", 1864=>x"8300", 1865=>x"8900", 1866=>x"8700", 1867=>x"8500", 1868=>x"8800", 1869=>x"8d00",
---- 1870=>x"8d00", 1871=>x"8e00", 1872=>x"8600", 1873=>x"8600", 1874=>x"8500", 1875=>x"8800", 1876=>x"8800",
---- 1877=>x"8900", 1878=>x"8d00", 1879=>x"8b00", 1880=>x"8a00", 1881=>x"8600", 1882=>x"8700", 1883=>x"8900",
---- 1884=>x"8a00", 1885=>x"8c00", 1886=>x"8d00", 1887=>x"8c00", 1888=>x"8a00", 1889=>x"8700", 1890=>x"8800",
---- 1891=>x"8b00", 1892=>x"8b00", 1893=>x"8b00", 1894=>x"8b00", 1895=>x"8b00", 1896=>x"8800", 1897=>x"8900",
---- 1898=>x"8900", 1899=>x"8900", 1900=>x"8900", 1901=>x"8900", 1902=>x"8b00", 1903=>x"8b00", 1904=>x"8500",
---- 1905=>x"8900", 1906=>x"8c00", 1907=>x"8b00", 1908=>x"8b00", 1909=>x"8b00", 1910=>x"8b00", 1911=>x"8b00",
---- 1912=>x"8600", 1913=>x"8800", 1914=>x"8c00", 1915=>x"8c00", 1916=>x"8a00", 1917=>x"8a00", 1918=>x"8900",
---- 1919=>x"8c00", 1920=>x"8800", 1921=>x"8900", 1922=>x"8b00", 1923=>x"8b00", 1924=>x"8b00", 1925=>x"8a00",
---- 1926=>x"8a00", 1927=>x"8c00", 1928=>x"8700", 1929=>x"8b00", 1930=>x"8a00", 1931=>x"8c00", 1932=>x"8c00",
---- 1933=>x"8b00", 1934=>x"8900", 1935=>x"8a00", 1936=>x"8600", 1937=>x"8c00", 1938=>x"8b00", 1939=>x"8c00",
---- 1940=>x"8b00", 1941=>x"8900", 1942=>x"8c00", 1943=>x"7500", 1944=>x"8800", 1945=>x"8800", 1946=>x"8a00",
---- 1947=>x"8a00", 1948=>x"8900", 1949=>x"8c00", 1950=>x"8f00", 1951=>x"8b00", 1952=>x"8700", 1953=>x"8800",
---- 1954=>x"8900", 1955=>x"8700", 1956=>x"8900", 1957=>x"8e00", 1958=>x"8c00", 1959=>x"8d00", 1960=>x"8800",
---- 1961=>x"8b00", 1962=>x"8800", 1963=>x"8a00", 1964=>x"8a00", 1965=>x"8b00", 1966=>x"8c00", 1967=>x"8a00",
---- 1968=>x"8200", 1969=>x"8a00", 1970=>x"8700", 1971=>x"8800", 1972=>x"8b00", 1973=>x"8c00", 1974=>x"8b00",
---- 1975=>x"8900", 1976=>x"8100", 1977=>x"8600", 1978=>x"8700", 1979=>x"8b00", 1980=>x"8a00", 1981=>x"8800",
---- 1982=>x"8700", 1983=>x"8800", 1984=>x"8600", 1985=>x"8600", 1986=>x"8700", 1987=>x"8800", 1988=>x"8700",
---- 1989=>x"8600", 1990=>x"8800", 1991=>x"8c00", 1992=>x"8500", 1993=>x"8b00", 1994=>x"8a00", 1995=>x"8900",
---- 1996=>x"8700", 1997=>x"8900", 1998=>x"8800", 1999=>x"8b00", 2000=>x"8600", 2001=>x"8800", 2002=>x"8700",
---- 2003=>x"8700", 2004=>x"8600", 2005=>x"8b00", 2006=>x"8900", 2007=>x"8a00", 2008=>x"8400", 2009=>x"8600",
---- 2010=>x"8500", 2011=>x"8700", 2012=>x"8a00", 2013=>x"8a00", 2014=>x"8900", 2015=>x"8900", 2016=>x"8100",
---- 2017=>x"8700", 2018=>x"8500", 2019=>x"8500", 2020=>x"8a00", 2021=>x"8900", 2022=>x"8700", 2023=>x"8700",
---- 2024=>x"8700", 2025=>x"8700", 2026=>x"8b00", 2027=>x"8900", 2028=>x"8800", 2029=>x"8500", 2030=>x"8500",
---- 2031=>x"8700", 2032=>x"8500", 2033=>x"8600", 2034=>x"8800", 2035=>x"8900", 2036=>x"8a00", 2037=>x"8900",
---- 2038=>x"8400", 2039=>x"8600", 2040=>x"8200", 2041=>x"8400", 2042=>x"8800", 2043=>x"8a00", 2044=>x"8b00",
---- 2045=>x"8800", 2046=>x"8500", 2047=>x"8500"),
---- 16 => (0=>x"8c00", 1=>x"8800", 2=>x"8200", 3=>x"8000", 4=>x"8400", 5=>x"8200", 6=>x"8500", 7=>x"8300",
---- 8=>x"8c00", 9=>x"8600", 10=>x"8200", 11=>x"8000", 12=>x"8500", 13=>x"8200", 14=>x"8500",
---- 15=>x"8300", 16=>x"8a00", 17=>x"8800", 18=>x"8300", 19=>x"7f00", 20=>x"8300", 21=>x"8400",
---- 22=>x"8300", 23=>x"8200", 24=>x"8300", 25=>x"8600", 26=>x"8400", 27=>x"8000", 28=>x"8000",
---- 29=>x"7f00", 30=>x"7e00", 31=>x"8300", 32=>x"8300", 33=>x"8500", 34=>x"8200", 35=>x"8200",
---- 36=>x"8000", 37=>x"7f00", 38=>x"8100", 39=>x"8000", 40=>x"8100", 41=>x"8300", 42=>x"8200",
---- 43=>x"8400", 44=>x"8200", 45=>x"8100", 46=>x"7e00", 47=>x"7f00", 48=>x"8100", 49=>x"8200",
---- 50=>x"8200", 51=>x"8300", 52=>x"8300", 53=>x"8400", 54=>x"8100", 55=>x"8100", 56=>x"8100",
---- 57=>x"8300", 58=>x"8200", 59=>x"8200", 60=>x"8100", 61=>x"8200", 62=>x"8200", 63=>x"7f00",
---- 64=>x"8200", 65=>x"8100", 66=>x"8300", 67=>x"8200", 68=>x"8300", 69=>x"8300", 70=>x"8200",
---- 71=>x"7e00", 72=>x"8300", 73=>x"8300", 74=>x"8300", 75=>x"8400", 76=>x"8600", 77=>x"8100",
---- 78=>x"8100", 79=>x"7f00", 80=>x"8400", 81=>x"8300", 82=>x"8200", 83=>x"8000", 84=>x"8900",
---- 85=>x"8000", 86=>x"8100", 87=>x"7e00", 88=>x"8200", 89=>x"8200", 90=>x"8200", 91=>x"8100",
---- 92=>x"8200", 93=>x"8200", 94=>x"8100", 95=>x"8100", 96=>x"8100", 97=>x"8100", 98=>x"8300",
---- 99=>x"8300", 100=>x"8100", 101=>x"8200", 102=>x"8000", 103=>x"7f00", 104=>x"8300", 105=>x"8400",
---- 106=>x"8300", 107=>x"8400", 108=>x"7f00", 109=>x"7f00", 110=>x"7f00", 111=>x"7e00", 112=>x"8200",
---- 113=>x"8400", 114=>x"8500", 115=>x"8400", 116=>x"8100", 117=>x"7e00", 118=>x"7f00", 119=>x"7f00",
---- 120=>x"8500", 121=>x"8100", 122=>x"8400", 123=>x"8200", 124=>x"7f00", 125=>x"7d00", 126=>x"8000",
---- 127=>x"7f00", 128=>x"8500", 129=>x"8300", 130=>x"8300", 131=>x"8100", 132=>x"8000", 133=>x"7d00",
---- 134=>x"7e00", 135=>x"7e00", 136=>x"8300", 137=>x"8500", 138=>x"8300", 139=>x"8100", 140=>x"7f00",
---- 141=>x"8100", 142=>x"8000", 143=>x"8000", 144=>x"8300", 145=>x"8400", 146=>x"8400", 147=>x"8000",
---- 148=>x"7f00", 149=>x"8000", 150=>x"8100", 151=>x"8000", 152=>x"8600", 153=>x"8200", 154=>x"8200",
---- 155=>x"8200", 156=>x"7e00", 157=>x"8100", 158=>x"7f00", 159=>x"7f00", 160=>x"8300", 161=>x"8200",
---- 162=>x"7f00", 163=>x"7e00", 164=>x"7d00", 165=>x"8100", 166=>x"7f00", 167=>x"7c00", 168=>x"8000",
---- 169=>x"8400", 170=>x"8000", 171=>x"8000", 172=>x"8300", 173=>x"8000", 174=>x"7e00", 175=>x"7f00",
---- 176=>x"7c00", 177=>x"7d00", 178=>x"7c00", 179=>x"7e00", 180=>x"7f00", 181=>x"7f00", 182=>x"7e00",
---- 183=>x"8000", 184=>x"7800", 185=>x"7d00", 186=>x"7b00", 187=>x"7c00", 188=>x"7d00", 189=>x"7d00",
---- 190=>x"7c00", 191=>x"7f00", 192=>x"7600", 193=>x"7800", 194=>x"7a00", 195=>x"7c00", 196=>x"7c00",
---- 197=>x"7c00", 198=>x"7d00", 199=>x"7d00", 200=>x"7400", 201=>x"7100", 202=>x"7100", 203=>x"7900",
---- 204=>x"7900", 205=>x"7a00", 206=>x"7c00", 207=>x"7a00", 208=>x"a700", 209=>x"8f00", 210=>x"7700",
---- 211=>x"6f00", 212=>x"7500", 213=>x"7600", 214=>x"7900", 215=>x"7800", 216=>x"c400", 217=>x"c000",
---- 218=>x"b100", 219=>x"8900", 220=>x"7200", 221=>x"7000", 222=>x"7700", 223=>x"7800", 224=>x"c200",
---- 225=>x"c600", 226=>x"c800", 227=>x"c200", 228=>x"a500", 229=>x"7c00", 230=>x"6f00", 231=>x"7300",
---- 232=>x"c100", 233=>x"c400", 234=>x"c200", 235=>x"c500", 236=>x"c600", 237=>x"bb00", 238=>x"8e00",
---- 239=>x"9100", 240=>x"c100", 241=>x"c400", 242=>x"c000", 243=>x"c100", 244=>x"c300", 245=>x"cb00",
---- 246=>x"c400", 247=>x"a200", 248=>x"bc00", 249=>x"c200", 250=>x"c200", 251=>x"c100", 252=>x"c600",
---- 253=>x"c500", 254=>x"ca00", 255=>x"c800", 256=>x"bd00", 257=>x"bb00", 258=>x"bf00", 259=>x"c100",
---- 260=>x"c500", 261=>x"c400", 262=>x"c400", 263=>x"c200", 264=>x"b800", 265=>x"bf00", 266=>x"c200",
---- 267=>x"c100", 268=>x"c500", 269=>x"c300", 270=>x"c400", 271=>x"c500", 272=>x"bd00", 273=>x"bd00",
---- 274=>x"c000", 275=>x"c300", 276=>x"c400", 277=>x"c300", 278=>x"c700", 279=>x"c500", 280=>x"c100",
---- 281=>x"be00", 282=>x"bd00", 283=>x"c300", 284=>x"c300", 285=>x"c600", 286=>x"c500", 287=>x"c400",
---- 288=>x"bf00", 289=>x"bf00", 290=>x"c400", 291=>x"c300", 292=>x"c400", 293=>x"c400", 294=>x"c400",
---- 295=>x"c400", 296=>x"c100", 297=>x"3d00", 298=>x"c100", 299=>x"c700", 300=>x"c400", 301=>x"c400",
---- 302=>x"c400", 303=>x"c000", 304=>x"be00", 305=>x"c100", 306=>x"c400", 307=>x"c500", 308=>x"c300",
---- 309=>x"c300", 310=>x"c500", 311=>x"c000", 312=>x"c400", 313=>x"b900", 314=>x"c300", 315=>x"c500",
---- 316=>x"c300", 317=>x"c000", 318=>x"c000", 319=>x"bc00", 320=>x"c000", 321=>x"c000", 322=>x"c400",
---- 323=>x"bc00", 324=>x"ba00", 325=>x"b900", 326=>x"b900", 327=>x"b900", 328=>x"c100", 329=>x"bc00",
---- 330=>x"b000", 331=>x"b100", 332=>x"b800", 333=>x"bc00", 334=>x"cb00", 335=>x"d300", 336=>x"ab00",
---- 337=>x"ab00", 338=>x"b100", 339=>x"be00", 340=>x"ce00", 341=>x"d400", 342=>x"d300", 343=>x"d500",
---- 344=>x"b400", 345=>x"c500", 346=>x"cf00", 347=>x"d700", 348=>x"d500", 349=>x"d200", 350=>x"cd00",
---- 351=>x"cd00", 352=>x"d100", 353=>x"d500", 354=>x"d500", 355=>x"d500", 356=>x"d200", 357=>x"ce00",
---- 358=>x"c800", 359=>x"3500", 360=>x"d200", 361=>x"d600", 362=>x"ce00", 363=>x"cb00", 364=>x"cb00",
---- 365=>x"cd00", 366=>x"d000", 367=>x"c900", 368=>x"ca00", 369=>x"cb00", 370=>x"c900", 371=>x"ce00",
---- 372=>x"d500", 373=>x"d000", 374=>x"cd00", 375=>x"cb00", 376=>x"c800", 377=>x"c900", 378=>x"cf00",
---- 379=>x"d700", 380=>x"d000", 381=>x"d000", 382=>x"cc00", 383=>x"c900", 384=>x"c900", 385=>x"d200",
---- 386=>x"ca00", 387=>x"ce00", 388=>x"cc00", 389=>x"c500", 390=>x"c500", 391=>x"c400", 392=>x"cb00",
---- 393=>x"c600", 394=>x"ca00", 395=>x"c700", 396=>x"c300", 397=>x"c200", 398=>x"c300", 399=>x"c700",
---- 400=>x"ca00", 401=>x"c300", 402=>x"3a00", 403=>x"ca00", 404=>x"c400", 405=>x"cb00", 406=>x"c600",
---- 407=>x"c200", 408=>x"c500", 409=>x"3a00", 410=>x"c600", 411=>x"c900", 412=>x"ca00", 413=>x"c000",
---- 414=>x"c400", 415=>x"c500", 416=>x"c300", 417=>x"c600", 418=>x"3b00", 419=>x"c100", 420=>x"c400",
---- 421=>x"c800", 422=>x"cc00", 423=>x"cb00", 424=>x"b700", 425=>x"bc00", 426=>x"bc00", 427=>x"c400",
---- 428=>x"cc00", 429=>x"cd00", 430=>x"ce00", 431=>x"cc00", 432=>x"b700", 433=>x"c100", 434=>x"c900",
---- 435=>x"3800", 436=>x"c900", 437=>x"cd00", 438=>x"cc00", 439=>x"ce00", 440=>x"c700", 441=>x"c300",
---- 442=>x"c400", 443=>x"ca00", 444=>x"c500", 445=>x"c900", 446=>x"cc00", 447=>x"cb00", 448=>x"c400",
---- 449=>x"c500", 450=>x"c000", 451=>x"c200", 452=>x"c700", 453=>x"c600", 454=>x"cd00", 455=>x"ce00",
---- 456=>x"c200", 457=>x"c500", 458=>x"ca00", 459=>x"c100", 460=>x"c300", 461=>x"cc00", 462=>x"c700",
---- 463=>x"3100", 464=>x"c900", 465=>x"c200", 466=>x"c500", 467=>x"c700", 468=>x"c400", 469=>x"c600",
---- 470=>x"c500", 471=>x"c400", 472=>x"c400", 473=>x"c400", 474=>x"bd00", 475=>x"c800", 476=>x"c400",
---- 477=>x"c000", 478=>x"c600", 479=>x"c600", 480=>x"c300", 481=>x"c400", 482=>x"c400", 483=>x"4200",
---- 484=>x"c400", 485=>x"c100", 486=>x"c000", 487=>x"c200", 488=>x"bf00", 489=>x"c500", 490=>x"c200",
---- 491=>x"c300", 492=>x"be00", 493=>x"be00", 494=>x"bb00", 495=>x"b700", 496=>x"ba00", 497=>x"c000",
---- 498=>x"c600", 499=>x"c200", 500=>x"ba00", 501=>x"b100", 502=>x"c100", 503=>x"c300", 504=>x"c200",
---- 505=>x"bc00", 506=>x"b600", 507=>x"b300", 508=>x"b400", 509=>x"c600", 510=>x"c900", 511=>x"ca00",
---- 512=>x"b600", 513=>x"b300", 514=>x"ad00", 515=>x"bd00", 516=>x"c000", 517=>x"c400", 518=>x"c800",
---- 519=>x"c700", 520=>x"a400", 521=>x"ac00", 522=>x"c000", 523=>x"c000", 524=>x"bc00", 525=>x"be00",
---- 526=>x"c500", 527=>x"c800", 528=>x"b100", 529=>x"c000", 530=>x"bf00", 531=>x"bc00", 532=>x"b500",
---- 533=>x"bc00", 534=>x"c100", 535=>x"c300", 536=>x"b500", 537=>x"b300", 538=>x"be00", 539=>x"bf00",
---- 540=>x"b800", 541=>x"b400", 542=>x"bc00", 543=>x"bf00", 544=>x"b700", 545=>x"b100", 546=>x"b500",
---- 547=>x"bf00", 548=>x"c100", 549=>x"b900", 550=>x"b800", 551=>x"c000", 552=>x"bb00", 553=>x"b500",
---- 554=>x"b600", 555=>x"b500", 556=>x"b200", 557=>x"bd00", 558=>x"bd00", 559=>x"b500", 560=>x"b900",
---- 561=>x"bb00", 562=>x"b200", 563=>x"b400", 564=>x"af00", 565=>x"ae00", 566=>x"b400", 567=>x"ba00",
---- 568=>x"b000", 569=>x"b500", 570=>x"b500", 571=>x"ac00", 572=>x"b700", 573=>x"b500", 574=>x"a700",
---- 575=>x"b500", 576=>x"af00", 577=>x"b000", 578=>x"ae00", 579=>x"b400", 580=>x"af00", 581=>x"b700",
---- 582=>x"b500", 583=>x"af00", 584=>x"ad00", 585=>x"b200", 586=>x"a900", 587=>x"ad00", 588=>x"b800",
---- 589=>x"ac00", 590=>x"b900", 591=>x"c300", 592=>x"b000", 593=>x"ad00", 594=>x"a900", 595=>x"5800",
---- 596=>x"ac00", 597=>x"b500", 598=>x"4900", 599=>x"bc00", 600=>x"b200", 601=>x"ad00", 602=>x"ae00",
---- 603=>x"aa00", 604=>x"a800", 605=>x"ac00", 606=>x"b200", 607=>x"ae00", 608=>x"b200", 609=>x"b200",
---- 610=>x"ae00", 611=>x"aa00", 612=>x"a900", 613=>x"a800", 614=>x"a900", 615=>x"ad00", 616=>x"a400",
---- 617=>x"a100", 618=>x"a700", 619=>x"b100", 620=>x"a800", 621=>x"a000", 622=>x"a800", 623=>x"ae00",
---- 624=>x"a500", 625=>x"9f00", 626=>x"9d00", 627=>x"a500", 628=>x"ac00", 629=>x"ac00", 630=>x"aa00",
---- 631=>x"a800", 632=>x"a900", 633=>x"a700", 634=>x"a600", 635=>x"a500", 636=>x"a400", 637=>x"ac00",
---- 638=>x"a100", 639=>x"9500", 640=>x"a000", 641=>x"a800", 642=>x"ac00", 643=>x"aa00", 644=>x"9900",
---- 645=>x"9800", 646=>x"a100", 647=>x"a300", 648=>x"ad00", 649=>x"9b00", 650=>x"9800", 651=>x"9a00",
---- 652=>x"a600", 653=>x"a100", 654=>x"a300", 655=>x"a600", 656=>x"9e00", 657=>x"8800", 658=>x"9800",
---- 659=>x"ab00", 660=>x"a800", 661=>x"a700", 662=>x"5c00", 663=>x"a800", 664=>x"9800", 665=>x"a000",
---- 666=>x"5e00", 667=>x"a600", 668=>x"aa00", 669=>x"9d00", 670=>x"a500", 671=>x"a900", 672=>x"a700",
---- 673=>x"a700", 674=>x"a300", 675=>x"a200", 676=>x"a100", 677=>x"a200", 678=>x"a000", 679=>x"9e00",
---- 680=>x"a100", 681=>x"a200", 682=>x"9e00", 683=>x"9d00", 684=>x"9d00", 685=>x"a300", 686=>x"a400",
---- 687=>x"a300", 688=>x"a200", 689=>x"a700", 690=>x"a600", 691=>x"a200", 692=>x"8f00", 693=>x"8900",
---- 694=>x"9300", 695=>x"9900", 696=>x"7b00", 697=>x"8100", 698=>x"8400", 699=>x"a400", 700=>x"a700",
---- 701=>x"9900", 702=>x"6300", 703=>x"9100", 704=>x"7900", 705=>x"7400", 706=>x"6500", 707=>x"6000",
---- 708=>x"7500", 709=>x"8700", 710=>x"9100", 711=>x"9700", 712=>x"7a00", 713=>x"6e00", 714=>x"5900",
---- 715=>x"4900", 716=>x"5600", 717=>x"5d00", 718=>x"4a00", 719=>x"4f00", 720=>x"4600", 721=>x"3f00",
---- 722=>x"3f00", 723=>x"6d00", 724=>x"7800", 725=>x"4000", 726=>x"be00", 727=>x"4900", 728=>x"3400",
---- 729=>x"4f00", 730=>x"7300", 731=>x"5c00", 732=>x"4700", 733=>x"3f00", 734=>x"4600", 735=>x"5400",
---- 736=>x"6100", 737=>x"6500", 738=>x"4d00", 739=>x"4900", 740=>x"4f00", 741=>x"4400", 742=>x"4800",
---- 743=>x"4f00", 744=>x"6a00", 745=>x"5800", 746=>x"7100", 747=>x"4700", 748=>x"3900", 749=>x"3000",
---- 750=>x"4900", 751=>x"6400", 752=>x"5500", 753=>x"7e00", 754=>x"5c00", 755=>x"4100", 756=>x"5700",
---- 757=>x"3800", 758=>x"4400", 759=>x"6d00", 760=>x"5f00", 761=>x"4f00", 762=>x"5500", 763=>x"6200",
---- 764=>x"4900", 765=>x"2500", 766=>x"4000", 767=>x"5b00", 768=>x"3f00", 769=>x"5100", 770=>x"7100",
---- 771=>x"4200", 772=>x"2700", 773=>x"2100", 774=>x"4e00", 775=>x"6100", 776=>x"4500", 777=>x"6200",
---- 778=>x"4a00", 779=>x"2200", 780=>x"2b00", 781=>x"2500", 782=>x"5d00", 783=>x"5a00", 784=>x"6100",
---- 785=>x"4700", 786=>x"1f00", 787=>x"3600", 788=>x"2f00", 789=>x"2600", 790=>x"6400", 791=>x"4100",
---- 792=>x"5d00", 793=>x"2000", 794=>x"3700", 795=>x"6b00", 796=>x"1d00", 797=>x"2b00", 798=>x"7d00",
---- 799=>x"7000", 800=>x"2f00", 801=>x"3100", 802=>x"7d00", 803=>x"a900", 804=>x"1400", 805=>x"5200",
---- 806=>x"a700", 807=>x"a700", 808=>x"2000", 809=>x"6a00", 810=>x"9500", 811=>x"2800", 812=>x"2600",
---- 813=>x"8900", 814=>x"6a00", 815=>x"7400", 816=>x"2200", 817=>x"7e00", 818=>x"6800", 819=>x"3700",
---- 820=>x"6d00", 821=>x"8000", 822=>x"6a00", 823=>x"6a00", 824=>x"3f00", 825=>x"8100", 826=>x"6b00",
---- 827=>x"8800", 828=>x"8d00", 829=>x"5400", 830=>x"6600", 831=>x"8a00", 832=>x"5b00", 833=>x"7500",
---- 834=>x"7200", 835=>x"8e00", 836=>x"7d00", 837=>x"6000", 838=>x"9800", 839=>x"a800", 840=>x"4f00",
---- 841=>x"6800", 842=>x"5700", 843=>x"8500", 844=>x"7900", 845=>x"9300", 846=>x"b100", 847=>x"a900",
---- 848=>x"5700", 849=>x"5000", 850=>x"5100", 851=>x"7a00", 852=>x"7700", 853=>x"8f00", 854=>x"9500",
---- 855=>x"a800", 856=>x"5b00", 857=>x"4c00", 858=>x"5e00", 859=>x"8600", 860=>x"8a00", 861=>x"9f00",
---- 862=>x"a500", 863=>x"b000", 864=>x"ae00", 865=>x"6400", 866=>x"8800", 867=>x"9c00", 868=>x"a000",
---- 869=>x"bb00", 870=>x"b000", 871=>x"b500", 872=>x"7900", 873=>x"9900", 874=>x"8c00", 875=>x"9e00",
---- 876=>x"ac00", 877=>x"b800", 878=>x"b600", 879=>x"b600", 880=>x"af00", 881=>x"a400", 882=>x"7b00",
---- 883=>x"9900", 884=>x"bb00", 885=>x"b300", 886=>x"b400", 887=>x"bb00", 888=>x"a800", 889=>x"a100",
---- 890=>x"8300", 891=>x"8700", 892=>x"b700", 893=>x"b600", 894=>x"ab00", 895=>x"bc00", 896=>x"a200",
---- 897=>x"a600", 898=>x"8e00", 899=>x"8700", 900=>x"a600", 901=>x"a900", 902=>x"a700", 903=>x"be00",
---- 904=>x"a500", 905=>x"a800", 906=>x"9200", 907=>x"8f00", 908=>x"b000", 909=>x"a100", 910=>x"ac00",
---- 911=>x"bf00", 912=>x"a500", 913=>x"ac00", 914=>x"9500", 915=>x"6d00", 916=>x"b100", 917=>x"ad00",
---- 918=>x"b400", 919=>x"bf00", 920=>x"af00", 921=>x"b200", 922=>x"9e00", 923=>x"9200", 924=>x"a500",
---- 925=>x"a600", 926=>x"b900", 927=>x"c300", 928=>x"b500", 929=>x"b400", 930=>x"9c00", 931=>x"6f00",
---- 932=>x"a000", 933=>x"a600", 934=>x"ba00", 935=>x"c900", 936=>x"ba00", 937=>x"b700", 938=>x"9700",
---- 939=>x"8300", 940=>x"a100", 941=>x"b300", 942=>x"c000", 943=>x"c000", 944=>x"bb00", 945=>x"b900",
---- 946=>x"5900", 947=>x"7f00", 948=>x"9d00", 949=>x"bc00", 950=>x"c000", 951=>x"5200", 952=>x"ba00",
---- 953=>x"ba00", 954=>x"b500", 955=>x"9500", 956=>x"a700", 957=>x"4500", 958=>x"ab00", 959=>x"a800",
---- 960=>x"b700", 961=>x"4500", 962=>x"b600", 963=>x"aa00", 964=>x"b400", 965=>x"b100", 966=>x"a900",
---- 967=>x"a200", 968=>x"ba00", 969=>x"bd00", 970=>x"b600", 971=>x"b300", 972=>x"b900", 973=>x"a900",
---- 974=>x"8a00", 975=>x"8400", 976=>x"c000", 977=>x"bf00", 978=>x"be00", 979=>x"bb00", 980=>x"9100",
---- 981=>x"5600", 982=>x"5300", 983=>x"9200", 984=>x"c200", 985=>x"c500", 986=>x"b800", 987=>x"8000",
---- 988=>x"5200", 989=>x"5800", 990=>x"6300", 991=>x"6300", 992=>x"c600", 993=>x"b300", 994=>x"8200",
---- 995=>x"7400", 996=>x"8800", 997=>x"8e00", 998=>x"8a00", 999=>x"8000", 1000=>x"a800", 1001=>x"7a00",
---- 1002=>x"7f00", 1003=>x"9100", 1004=>x"9a00", 1005=>x"9700", 1006=>x"9500", 1007=>x"9f00", 1008=>x"7000",
---- 1009=>x"7d00", 1010=>x"8300", 1011=>x"8c00", 1012=>x"9100", 1013=>x"8f00", 1014=>x"7900", 1015=>x"8e00",
---- 1016=>x"7100", 1017=>x"7300", 1018=>x"7100", 1019=>x"7800", 1020=>x"7700", 1021=>x"7d00", 1022=>x"5000",
---- 1023=>x"5800", 1024=>x"5f00", 1025=>x"6000", 1026=>x"5100", 1027=>x"4b00", 1028=>x"4d00", 1029=>x"4c00",
---- 1030=>x"3200", 1031=>x"3800", 1032=>x"3a00", 1033=>x"3e00", 1034=>x"3b00", 1035=>x"3600", 1036=>x"3300",
---- 1037=>x"3100", 1038=>x"3100", 1039=>x"3300", 1040=>x"3300", 1041=>x"3300", 1042=>x"3500", 1043=>x"3200",
---- 1044=>x"3000", 1045=>x"2e00", 1046=>x"2d00", 1047=>x"3400", 1048=>x"2f00", 1049=>x"3100", 1050=>x"3200",
---- 1051=>x"3000", 1052=>x"2c00", 1053=>x"3000", 1054=>x"3400", 1055=>x"4c00", 1056=>x"4100", 1057=>x"3d00",
---- 1058=>x"3300", 1059=>x"3b00", 1060=>x"2300", 1061=>x"3000", 1062=>x"4c00", 1063=>x"5000", 1064=>x"5e00",
---- 1065=>x"5500", 1066=>x"3f00", 1067=>x"5d00", 1068=>x"3200", 1069=>x"3000", 1070=>x"6000", 1071=>x"3300",
---- 1072=>x"6000", 1073=>x"7500", 1074=>x"4500", 1075=>x"4f00", 1076=>x"5900", 1077=>x"5600", 1078=>x"4600",
---- 1079=>x"4c00", 1080=>x"5d00", 1081=>x"7800", 1082=>x"6c00", 1083=>x"4300", 1084=>x"3e00", 1085=>x"4000",
---- 1086=>x"4d00", 1087=>x"9c00", 1088=>x"6100", 1089=>x"7100", 1090=>x"8000", 1091=>x"7a00", 1092=>x"6100",
---- 1093=>x"6e00", 1094=>x"a200", 1095=>x"c600", 1096=>x"5f00", 1097=>x"5f00", 1098=>x"7c00", 1099=>x"8700",
---- 1100=>x"9400", 1101=>x"9d00", 1102=>x"a900", 1103=>x"b400", 1104=>x"7b00", 1105=>x"7e00", 1106=>x"6d00",
---- 1107=>x"7100", 1108=>x"7100", 1109=>x"7900", 1110=>x"8c00", 1111=>x"8d00", 1112=>x"9000", 1113=>x"8800",
---- 1114=>x"8d00", 1115=>x"7b00", 1116=>x"6700", 1117=>x"7200", 1118=>x"8800", 1119=>x"7e00", 1120=>x"9700",
---- 1121=>x"8e00", 1122=>x"8500", 1123=>x"8a00", 1124=>x"7e00", 1125=>x"8300", 1126=>x"8800", 1127=>x"8a00",
---- 1128=>x"6c00", 1129=>x"9100", 1130=>x"9000", 1131=>x"9200", 1132=>x"8d00", 1133=>x"8d00", 1134=>x"8d00",
---- 1135=>x"9400", 1136=>x"9c00", 1137=>x"9600", 1138=>x"9500", 1139=>x"9800", 1140=>x"9600", 1141=>x"9900",
---- 1142=>x"9c00", 1143=>x"a100", 1144=>x"aa00", 1145=>x"aa00", 1146=>x"a300", 1147=>x"a400", 1148=>x"a400",
---- 1149=>x"a300", 1150=>x"ab00", 1151=>x"ad00", 1152=>x"ac00", 1153=>x"b000", 1154=>x"ab00", 1155=>x"a600",
---- 1156=>x"a700", 1157=>x"a700", 1158=>x"ac00", 1159=>x"af00", 1160=>x"ac00", 1161=>x"af00", 1162=>x"ab00",
---- 1163=>x"b000", 1164=>x"b000", 1165=>x"ad00", 1166=>x"ad00", 1167=>x"ab00", 1168=>x"ac00", 1169=>x"b400",
---- 1170=>x"af00", 1171=>x"ab00", 1172=>x"b200", 1173=>x"b100", 1174=>x"b200", 1175=>x"af00", 1176=>x"ad00",
---- 1177=>x"b100", 1178=>x"b300", 1179=>x"b000", 1180=>x"b000", 1181=>x"b200", 1182=>x"b100", 1183=>x"b000",
---- 1184=>x"ae00", 1185=>x"b300", 1186=>x"b300", 1187=>x"b300", 1188=>x"b300", 1189=>x"b000", 1190=>x"ae00",
---- 1191=>x"af00", 1192=>x"ae00", 1193=>x"b200", 1194=>x"b200", 1195=>x"b200", 1196=>x"b700", 1197=>x"b800",
---- 1198=>x"af00", 1199=>x"ac00", 1200=>x"a700", 1201=>x"ad00", 1202=>x"b200", 1203=>x"b300", 1204=>x"af00",
---- 1205=>x"b400", 1206=>x"b100", 1207=>x"ad00", 1208=>x"a600", 1209=>x"a800", 1210=>x"ac00", 1211=>x"af00",
---- 1212=>x"af00", 1213=>x"b300", 1214=>x"b100", 1215=>x"ab00", 1216=>x"a700", 1217=>x"a900", 1218=>x"ad00",
---- 1219=>x"af00", 1220=>x"ad00", 1221=>x"af00", 1222=>x"b000", 1223=>x"5500", 1224=>x"9f00", 1225=>x"a300",
---- 1226=>x"a900", 1227=>x"ae00", 1228=>x"a800", 1229=>x"aa00", 1230=>x"ac00", 1231=>x"ac00", 1232=>x"a200",
---- 1233=>x"9f00", 1234=>x"a100", 1235=>x"a900", 1236=>x"a700", 1237=>x"a800", 1238=>x"a800", 1239=>x"a900",
---- 1240=>x"a100", 1241=>x"9f00", 1242=>x"9d00", 1243=>x"a100", 1244=>x"a400", 1245=>x"a600", 1246=>x"a500",
---- 1247=>x"a800", 1248=>x"9a00", 1249=>x"9d00", 1250=>x"9c00", 1251=>x"9b00", 1252=>x"9e00", 1253=>x"a300",
---- 1254=>x"a500", 1255=>x"a400", 1256=>x"6900", 1257=>x"9800", 1258=>x"9a00", 1259=>x"9c00", 1260=>x"9f00",
---- 1261=>x"a100", 1262=>x"a300", 1263=>x"a000", 1264=>x"9700", 1265=>x"9800", 1266=>x"9900", 1267=>x"9c00",
---- 1268=>x"9d00", 1269=>x"9e00", 1270=>x"9f00", 1271=>x"a000", 1272=>x"9700", 1273=>x"9700", 1274=>x"9e00",
---- 1275=>x"9c00", 1276=>x"9d00", 1277=>x"9d00", 1278=>x"9f00", 1279=>x"a100", 1280=>x"9700", 1281=>x"9600",
---- 1282=>x"9600", 1283=>x"9800", 1284=>x"9c00", 1285=>x"9b00", 1286=>x"9c00", 1287=>x"a000", 1288=>x"9600",
---- 1289=>x"9800", 1290=>x"9900", 1291=>x"9700", 1292=>x"9a00", 1293=>x"9b00", 1294=>x"9d00", 1295=>x"9e00",
---- 1296=>x"9700", 1297=>x"9700", 1298=>x"9900", 1299=>x"9500", 1300=>x"9b00", 1301=>x"9b00", 1302=>x"9f00",
---- 1303=>x"9d00", 1304=>x"9700", 1305=>x"9300", 1306=>x"9600", 1307=>x"9800", 1308=>x"9b00", 1309=>x"9900",
---- 1310=>x"9c00", 1311=>x"9c00", 1312=>x"9400", 1313=>x"9000", 1314=>x"9500", 1315=>x"9300", 1316=>x"9b00",
---- 1317=>x"9600", 1318=>x"9700", 1319=>x"6200", 1320=>x"9000", 1321=>x"9200", 1322=>x"9700", 1323=>x"9400",
---- 1324=>x"9b00", 1325=>x"9900", 1326=>x"9b00", 1327=>x"9b00", 1328=>x"9000", 1329=>x"9000", 1330=>x"9000",
---- 1331=>x"9400", 1332=>x"9a00", 1333=>x"9a00", 1334=>x"9b00", 1335=>x"9c00", 1336=>x"8f00", 1337=>x"9000",
---- 1338=>x"9400", 1339=>x"9800", 1340=>x"9900", 1341=>x"9900", 1342=>x"9a00", 1343=>x"9c00", 1344=>x"8a00",
---- 1345=>x"8c00", 1346=>x"9000", 1347=>x"9300", 1348=>x"9700", 1349=>x"9700", 1350=>x"9800", 1351=>x"6600",
---- 1352=>x"8e00", 1353=>x"8d00", 1354=>x"8e00", 1355=>x"8e00", 1356=>x"9200", 1357=>x"9600", 1358=>x"9500",
---- 1359=>x"9700", 1360=>x"8f00", 1361=>x"8c00", 1362=>x"8d00", 1363=>x"8e00", 1364=>x"8c00", 1365=>x"9100",
---- 1366=>x"9400", 1367=>x"9500", 1368=>x"8c00", 1369=>x"8800", 1370=>x"8a00", 1371=>x"8b00", 1372=>x"8c00",
---- 1373=>x"8e00", 1374=>x"9000", 1375=>x"9100", 1376=>x"8a00", 1377=>x"8700", 1378=>x"8900", 1379=>x"8c00",
---- 1380=>x"8f00", 1381=>x"8e00", 1382=>x"8900", 1383=>x"8c00", 1384=>x"8c00", 1385=>x"8700", 1386=>x"8800",
---- 1387=>x"8d00", 1388=>x"8a00", 1389=>x"8a00", 1390=>x"8700", 1391=>x"8400", 1392=>x"8e00", 1393=>x"8c00",
---- 1394=>x"8c00", 1395=>x"9200", 1396=>x"8800", 1397=>x"6d00", 1398=>x"6300", 1399=>x"8f00", 1400=>x"8f00",
---- 1401=>x"9000", 1402=>x"8f00", 1403=>x"9200", 1404=>x"8200", 1405=>x"5c00", 1406=>x"5000", 1407=>x"5100",
---- 1408=>x"9000", 1409=>x"9400", 1410=>x"9100", 1411=>x"9100", 1412=>x"8300", 1413=>x"7600", 1414=>x"7a00",
---- 1415=>x"7400", 1416=>x"9100", 1417=>x"9300", 1418=>x"9200", 1419=>x"9100", 1420=>x"8e00", 1421=>x"8b00",
---- 1422=>x"8100", 1423=>x"8100", 1424=>x"8f00", 1425=>x"9300", 1426=>x"9100", 1427=>x"8f00", 1428=>x"9600",
---- 1429=>x"8f00", 1430=>x"8500", 1431=>x"8100", 1432=>x"8a00", 1433=>x"8e00", 1434=>x"8f00", 1435=>x"9300",
---- 1436=>x"9300", 1437=>x"9000", 1438=>x"8a00", 1439=>x"8800", 1440=>x"8700", 1441=>x"8c00", 1442=>x"8d00",
---- 1443=>x"9000", 1444=>x"9300", 1445=>x"9000", 1446=>x"8c00", 1447=>x"8800", 1448=>x"8800", 1449=>x"8900",
---- 1450=>x"8a00", 1451=>x"8b00", 1452=>x"8c00", 1453=>x"8e00", 1454=>x"8e00", 1455=>x"8900", 1456=>x"8600",
---- 1457=>x"8900", 1458=>x"8a00", 1459=>x"8c00", 1460=>x"8b00", 1461=>x"8f00", 1462=>x"8d00", 1463=>x"8b00",
---- 1464=>x"8300", 1465=>x"7900", 1466=>x"8a00", 1467=>x"8900", 1468=>x"8c00", 1469=>x"8e00", 1470=>x"8c00",
---- 1471=>x"8b00", 1472=>x"8400", 1473=>x"8500", 1474=>x"8700", 1475=>x"8a00", 1476=>x"8900", 1477=>x"8d00",
---- 1478=>x"8900", 1479=>x"8900", 1480=>x"8600", 1481=>x"8400", 1482=>x"8800", 1483=>x"7600", 1484=>x"8800",
---- 1485=>x"8b00", 1486=>x"8900", 1487=>x"8a00", 1488=>x"8300", 1489=>x"8700", 1490=>x"8800", 1491=>x"8900",
---- 1492=>x"8a00", 1493=>x"8b00", 1494=>x"8b00", 1495=>x"7100", 1496=>x"8400", 1497=>x"8400", 1498=>x"8400",
---- 1499=>x"8900", 1500=>x"8a00", 1501=>x"8a00", 1502=>x"8e00", 1503=>x"8d00", 1504=>x"8100", 1505=>x"8200",
---- 1506=>x"8400", 1507=>x"8600", 1508=>x"8900", 1509=>x"8b00", 1510=>x"9100", 1511=>x"9200", 1512=>x"7d00",
---- 1513=>x"8100", 1514=>x"8400", 1515=>x"8700", 1516=>x"8600", 1517=>x"8c00", 1518=>x"9100", 1519=>x"9100",
---- 1520=>x"7900", 1521=>x"7c00", 1522=>x"7f00", 1523=>x"8400", 1524=>x"8700", 1525=>x"8900", 1526=>x"8b00",
---- 1527=>x"9200", 1528=>x"6900", 1529=>x"7000", 1530=>x"7b00", 1531=>x"7c00", 1532=>x"8100", 1533=>x"8000",
---- 1534=>x"8800", 1535=>x"8a00", 1536=>x"4600", 1537=>x"4f00", 1538=>x"5c00", 1539=>x"6200", 1540=>x"6b00",
---- 1541=>x"7100", 1542=>x"7800", 1543=>x"7c00", 1544=>x"5900", 1545=>x"5d00", 1546=>x"6200", 1547=>x"6400",
---- 1548=>x"6600", 1549=>x"7200", 1550=>x"7900", 1551=>x"7900", 1552=>x"7f00", 1553=>x"8400", 1554=>x"8900",
---- 1555=>x"8b00", 1556=>x"8500", 1557=>x"8400", 1558=>x"8700", 1559=>x"8900", 1560=>x"8300", 1561=>x"8600",
---- 1562=>x"8c00", 1563=>x"8d00", 1564=>x"8a00", 1565=>x"8900", 1566=>x"8800", 1567=>x"8e00", 1568=>x"7d00",
---- 1569=>x"8000", 1570=>x"8400", 1571=>x"8500", 1572=>x"8600", 1573=>x"8400", 1574=>x"8600", 1575=>x"8800",
---- 1576=>x"7e00", 1577=>x"8000", 1578=>x"8400", 1579=>x"8400", 1580=>x"8500", 1581=>x"8500", 1582=>x"8a00",
---- 1583=>x"8a00", 1584=>x"7c00", 1585=>x"7e00", 1586=>x"8100", 1587=>x"8300", 1588=>x"8500", 1589=>x"8900",
---- 1590=>x"8a00", 1591=>x"8b00", 1592=>x"7d00", 1593=>x"8100", 1594=>x"7d00", 1595=>x"8200", 1596=>x"8a00",
---- 1597=>x"8900", 1598=>x"8800", 1599=>x"8800", 1600=>x"7c00", 1601=>x"7f00", 1602=>x"8000", 1603=>x"8200",
---- 1604=>x"8700", 1605=>x"8700", 1606=>x"8700", 1607=>x"8800", 1608=>x"7e00", 1609=>x"8100", 1610=>x"8300",
---- 1611=>x"7e00", 1612=>x"8100", 1613=>x"8700", 1614=>x"8600", 1615=>x"8b00", 1616=>x"7c00", 1617=>x"8200",
---- 1618=>x"7b00", 1619=>x"7c00", 1620=>x"8400", 1621=>x"8800", 1622=>x"8b00", 1623=>x"8d00", 1624=>x"7f00",
---- 1625=>x"7b00", 1626=>x"7c00", 1627=>x"8400", 1628=>x"8700", 1629=>x"8900", 1630=>x"8d00", 1631=>x"8f00",
---- 1632=>x"7a00", 1633=>x"7800", 1634=>x"8400", 1635=>x"8800", 1636=>x"8800", 1637=>x"8800", 1638=>x"8c00",
---- 1639=>x"8d00", 1640=>x"7200", 1641=>x"8000", 1642=>x"8800", 1643=>x"8b00", 1644=>x"8b00", 1645=>x"8700",
---- 1646=>x"8700", 1647=>x"8a00", 1648=>x"7c00", 1649=>x"8700", 1650=>x"8500", 1651=>x"8b00", 1652=>x"8b00",
---- 1653=>x"8800", 1654=>x"8a00", 1655=>x"8d00", 1656=>x"8400", 1657=>x"8600", 1658=>x"8800", 1659=>x"8b00",
---- 1660=>x"8a00", 1661=>x"8a00", 1662=>x"8c00", 1663=>x"8c00", 1664=>x"7f00", 1665=>x"8800", 1666=>x"8a00",
---- 1667=>x"8b00", 1668=>x"8a00", 1669=>x"8a00", 1670=>x"8c00", 1671=>x"8a00", 1672=>x"8000", 1673=>x"8600",
---- 1674=>x"8900", 1675=>x"8800", 1676=>x"8d00", 1677=>x"8a00", 1678=>x"8d00", 1679=>x"8a00", 1680=>x"8500",
---- 1681=>x"8300", 1682=>x"8600", 1683=>x"8900", 1684=>x"8a00", 1685=>x"8d00", 1686=>x"8d00", 1687=>x"8c00",
---- 1688=>x"8500", 1689=>x"8500", 1690=>x"8600", 1691=>x"8700", 1692=>x"8a00", 1693=>x"8b00", 1694=>x"8d00",
---- 1695=>x"8b00", 1696=>x"8800", 1697=>x"8800", 1698=>x"8300", 1699=>x"8300", 1700=>x"8a00", 1701=>x"8700",
---- 1702=>x"8d00", 1703=>x"8d00", 1704=>x"8600", 1705=>x"8600", 1706=>x"8600", 1707=>x"8700", 1708=>x"8b00",
---- 1709=>x"8800", 1710=>x"7400", 1711=>x"8d00", 1712=>x"8400", 1713=>x"8900", 1714=>x"8a00", 1715=>x"8a00",
---- 1716=>x"8c00", 1717=>x"8900", 1718=>x"8900", 1719=>x"8b00", 1720=>x"8800", 1721=>x"8900", 1722=>x"8800",
---- 1723=>x"8a00", 1724=>x"8b00", 1725=>x"8b00", 1726=>x"8400", 1727=>x"8900", 1728=>x"8800", 1729=>x"8900",
---- 1730=>x"8700", 1731=>x"8900", 1732=>x"7500", 1733=>x"8a00", 1734=>x"8900", 1735=>x"8700", 1736=>x"8600",
---- 1737=>x"8a00", 1738=>x"8a00", 1739=>x"8800", 1740=>x"8800", 1741=>x"8700", 1742=>x"8800", 1743=>x"8b00",
---- 1744=>x"8900", 1745=>x"8800", 1746=>x"8c00", 1747=>x"8900", 1748=>x"8800", 1749=>x"8800", 1750=>x"8700",
---- 1751=>x"8900", 1752=>x"8900", 1753=>x"8b00", 1754=>x"8a00", 1755=>x"8a00", 1756=>x"8a00", 1757=>x"8900",
---- 1758=>x"8700", 1759=>x"8900", 1760=>x"8a00", 1761=>x"8a00", 1762=>x"8c00", 1763=>x"8c00", 1764=>x"8900",
---- 1765=>x"8800", 1766=>x"8800", 1767=>x"8900", 1768=>x"8a00", 1769=>x"8b00", 1770=>x"9000", 1771=>x"8f00",
---- 1772=>x"8a00", 1773=>x"8800", 1774=>x"8900", 1775=>x"8800", 1776=>x"8900", 1777=>x"8c00", 1778=>x"8e00",
---- 1779=>x"8d00", 1780=>x"8a00", 1781=>x"8b00", 1782=>x"8b00", 1783=>x"8900", 1784=>x"8b00", 1785=>x"8900",
---- 1786=>x"8d00", 1787=>x"8b00", 1788=>x"8a00", 1789=>x"8800", 1790=>x"8a00", 1791=>x"8b00", 1792=>x"8b00",
---- 1793=>x"8c00", 1794=>x"8900", 1795=>x"8b00", 1796=>x"8c00", 1797=>x"8b00", 1798=>x"8c00", 1799=>x"8800",
---- 1800=>x"8a00", 1801=>x"8c00", 1802=>x"8c00", 1803=>x"8c00", 1804=>x"8f00", 1805=>x"8d00", 1806=>x"8900",
---- 1807=>x"8700", 1808=>x"8a00", 1809=>x"8a00", 1810=>x"8d00", 1811=>x"8f00", 1812=>x"8d00", 1813=>x"8c00",
---- 1814=>x"8d00", 1815=>x"8a00", 1816=>x"8c00", 1817=>x"9000", 1818=>x"8d00", 1819=>x"8a00", 1820=>x"8a00",
---- 1821=>x"8a00", 1822=>x"8a00", 1823=>x"7600", 1824=>x"8d00", 1825=>x"9200", 1826=>x"9000", 1827=>x"8b00",
---- 1828=>x"8b00", 1829=>x"8a00", 1830=>x"8a00", 1831=>x"8a00", 1832=>x"8c00", 1833=>x"8f00", 1834=>x"9500",
---- 1835=>x"8f00", 1836=>x"8b00", 1837=>x"8a00", 1838=>x"8c00", 1839=>x"8d00", 1840=>x"8d00", 1841=>x"9000",
---- 1842=>x"8f00", 1843=>x"9000", 1844=>x"8c00", 1845=>x"8c00", 1846=>x"8d00", 1847=>x"7100", 1848=>x"8f00",
---- 1849=>x"8f00", 1850=>x"8f00", 1851=>x"9100", 1852=>x"8f00", 1853=>x"8d00", 1854=>x"8c00", 1855=>x"8e00",
---- 1856=>x"8e00", 1857=>x"9200", 1858=>x"8f00", 1859=>x"8b00", 1860=>x"8b00", 1861=>x"8e00", 1862=>x"8f00",
---- 1863=>x"8d00", 1864=>x"8e00", 1865=>x"9200", 1866=>x"9000", 1867=>x"8a00", 1868=>x"8c00", 1869=>x"8f00",
---- 1870=>x"8d00", 1871=>x"8900", 1872=>x"8d00", 1873=>x"9000", 1874=>x"8e00", 1875=>x"8b00", 1876=>x"8c00",
---- 1877=>x"8e00", 1878=>x"8e00", 1879=>x"8c00", 1880=>x"8e00", 1881=>x"8c00", 1882=>x"8d00", 1883=>x"8e00",
---- 1884=>x"8f00", 1885=>x"8f00", 1886=>x"9000", 1887=>x"8b00", 1888=>x"8900", 1889=>x"8c00", 1890=>x"8d00",
---- 1891=>x"8e00", 1892=>x"8e00", 1893=>x"9000", 1894=>x"8e00", 1895=>x"8d00", 1896=>x"8a00", 1897=>x"8d00",
---- 1898=>x"8b00", 1899=>x"9000", 1900=>x"9000", 1901=>x"9000", 1902=>x"9000", 1903=>x"8e00", 1904=>x"8b00",
---- 1905=>x"8d00", 1906=>x"8a00", 1907=>x"9000", 1908=>x"8f00", 1909=>x"9100", 1910=>x"9000", 1911=>x"8e00",
---- 1912=>x"8b00", 1913=>x"8c00", 1914=>x"8a00", 1915=>x"9100", 1916=>x"8f00", 1917=>x"8e00", 1918=>x"8f00",
---- 1919=>x"8f00", 1920=>x"8c00", 1921=>x"8c00", 1922=>x"8c00", 1923=>x"8e00", 1924=>x"8f00", 1925=>x"8e00",
---- 1926=>x"8e00", 1927=>x"8d00", 1928=>x"8c00", 1929=>x"8900", 1930=>x"8900", 1931=>x"8a00", 1932=>x"9000",
---- 1933=>x"9100", 1934=>x"8d00", 1935=>x"8b00", 1936=>x"8c00", 1937=>x"8b00", 1938=>x"8c00", 1939=>x"8c00",
---- 1940=>x"9100", 1941=>x"9000", 1942=>x"8d00", 1943=>x"8c00", 1944=>x"8b00", 1945=>x"8c00", 1946=>x"8d00",
---- 1947=>x"8e00", 1948=>x"8e00", 1949=>x"8e00", 1950=>x"8f00", 1951=>x"9100", 1952=>x"8b00", 1953=>x"8b00",
---- 1954=>x"8e00", 1955=>x"8f00", 1956=>x"8f00", 1957=>x"8f00", 1958=>x"9000", 1959=>x"9100", 1960=>x"8800",
---- 1961=>x"8b00", 1962=>x"9000", 1963=>x"8e00", 1964=>x"8d00", 1965=>x"8f00", 1966=>x"8f00", 1967=>x"8f00",
---- 1968=>x"8a00", 1969=>x"8c00", 1970=>x"8c00", 1971=>x"8a00", 1972=>x"8c00", 1973=>x"8d00", 1974=>x"9200",
---- 1975=>x"8f00", 1976=>x"8c00", 1977=>x"8d00", 1978=>x"8e00", 1979=>x"8d00", 1980=>x"8e00", 1981=>x"8d00",
---- 1982=>x"9100", 1983=>x"8f00", 1984=>x"8e00", 1985=>x"8d00", 1986=>x"8c00", 1987=>x"8d00", 1988=>x"8f00",
---- 1989=>x"8d00", 1990=>x"8b00", 1991=>x"8e00", 1992=>x"8d00", 1993=>x"8c00", 1994=>x"8b00", 1995=>x"8c00",
---- 1996=>x"8f00", 1997=>x"8c00", 1998=>x"8d00", 1999=>x"8d00", 2000=>x"8b00", 2001=>x"8900", 2002=>x"8800",
---- 2003=>x"8c00", 2004=>x"8d00", 2005=>x"8d00", 2006=>x"8e00", 2007=>x"8d00", 2008=>x"8800", 2009=>x"8a00",
---- 2010=>x"8c00", 2011=>x"8c00", 2012=>x"8c00", 2013=>x"8b00", 2014=>x"8d00", 2015=>x"8a00", 2016=>x"8b00",
---- 2017=>x"7200", 2018=>x"8b00", 2019=>x"8a00", 2020=>x"8d00", 2021=>x"8b00", 2022=>x"8d00", 2023=>x"8c00",
---- 2024=>x"8d00", 2025=>x"8d00", 2026=>x"8a00", 2027=>x"8d00", 2028=>x"7100", 2029=>x"8a00", 2030=>x"8c00",
---- 2031=>x"8f00", 2032=>x"8800", 2033=>x"8800", 2034=>x"8b00", 2035=>x"8c00", 2036=>x"8c00", 2037=>x"8d00",
---- 2038=>x"8b00", 2039=>x"8e00", 2040=>x"8700", 2041=>x"8600", 2042=>x"8900", 2043=>x"8b00", 2044=>x"8b00",
---- 2045=>x"8d00", 2046=>x"8d00", 2047=>x"8b00"),
---- 17 => (0=>x"8000", 1=>x"8200", 2=>x"8100", 3=>x"8600", 4=>x"8200", 5=>x"7f00", 6=>x"8200", 7=>x"8300",
---- 8=>x"8000", 9=>x"8200", 10=>x"8100", 11=>x"8600", 12=>x"8200", 13=>x"7f00", 14=>x"8200",
---- 15=>x"8300", 16=>x"8000", 17=>x"8200", 18=>x"8000", 19=>x"8600", 20=>x"8100", 21=>x"7e00",
---- 22=>x"8100", 23=>x"8200", 24=>x"7f00", 25=>x"8000", 26=>x"8000", 27=>x"8000", 28=>x"7e00",
---- 29=>x"7e00", 30=>x"8100", 31=>x"8300", 32=>x"7f00", 33=>x"7f00", 34=>x"7f00", 35=>x"8000",
---- 36=>x"7d00", 37=>x"7e00", 38=>x"7f00", 39=>x"7f00", 40=>x"8000", 41=>x"8000", 42=>x"8000",
---- 43=>x"8000", 44=>x"7f00", 45=>x"8000", 46=>x"7e00", 47=>x"7f00", 48=>x"8000", 49=>x"8100",
---- 50=>x"8200", 51=>x"8100", 52=>x"7f00", 53=>x"8100", 54=>x"8000", 55=>x"8200", 56=>x"8000",
---- 57=>x"8100", 58=>x"7f00", 59=>x"7f00", 60=>x"8000", 61=>x"7f00", 62=>x"7f00", 63=>x"8100",
---- 64=>x"8200", 65=>x"8100", 66=>x"7f00", 67=>x"7f00", 68=>x"7f00", 69=>x"7b00", 70=>x"8000",
---- 71=>x"8100", 72=>x"7f00", 73=>x"8300", 74=>x"8200", 75=>x"8200", 76=>x"8100", 77=>x"7e00",
---- 78=>x"7f00", 79=>x"7e00", 80=>x"8100", 81=>x"8000", 82=>x"8000", 83=>x"8200", 84=>x"8300",
---- 85=>x"7e00", 86=>x"7d00", 87=>x"7f00", 88=>x"8000", 89=>x"8200", 90=>x"7e00", 91=>x"7c00",
---- 92=>x"7d00", 93=>x"7f00", 94=>x"7d00", 95=>x"8000", 96=>x"7f00", 97=>x"8200", 98=>x"8000",
---- 99=>x"7f00", 100=>x"7e00", 101=>x"7d00", 102=>x"7c00", 103=>x"7e00", 104=>x"7d00", 105=>x"7f00",
---- 106=>x"8000", 107=>x"7e00", 108=>x"8000", 109=>x"7e00", 110=>x"7e00", 111=>x"7f00", 112=>x"8000",
---- 113=>x"8000", 114=>x"8000", 115=>x"8000", 116=>x"7d00", 117=>x"7f00", 118=>x"7f00", 119=>x"7d00",
---- 120=>x"7d00", 121=>x"8200", 122=>x"7f00", 123=>x"8000", 124=>x"8100", 125=>x"7e00", 126=>x"7c00",
---- 127=>x"7f00", 128=>x"7c00", 129=>x"8200", 130=>x"8000", 131=>x"7d00", 132=>x"8000", 133=>x"7e00",
---- 134=>x"7c00", 135=>x"7f00", 136=>x"8000", 137=>x"8300", 138=>x"7e00", 139=>x"7e00", 140=>x"8100",
---- 141=>x"7d00", 142=>x"7d00", 143=>x"7e00", 144=>x"8000", 145=>x"7f00", 146=>x"8000", 147=>x"7e00",
---- 148=>x"7e00", 149=>x"7e00", 150=>x"7c00", 151=>x"7d00", 152=>x"8000", 153=>x"8200", 154=>x"8100",
---- 155=>x"7f00", 156=>x"7e00", 157=>x"8000", 158=>x"7e00", 159=>x"7d00", 160=>x"7f00", 161=>x"8000",
---- 162=>x"7f00", 163=>x"7f00", 164=>x"7e00", 165=>x"7d00", 166=>x"7e00", 167=>x"7f00", 168=>x"7b00",
---- 169=>x"7e00", 170=>x"8200", 171=>x"7a00", 172=>x"7f00", 173=>x"7c00", 174=>x"8200", 175=>x"8200",
---- 176=>x"7e00", 177=>x"8100", 178=>x"8100", 179=>x"8200", 180=>x"8200", 181=>x"7e00", 182=>x"8000",
---- 183=>x"8000", 184=>x"7f00", 185=>x"8100", 186=>x"8200", 187=>x"8100", 188=>x"8300", 189=>x"7f00",
---- 190=>x"8000", 191=>x"7d00", 192=>x"7f00", 193=>x"8200", 194=>x"8200", 195=>x"8100", 196=>x"8300",
---- 197=>x"8300", 198=>x"8200", 199=>x"7d00", 200=>x"7e00", 201=>x"8200", 202=>x"8300", 203=>x"8200",
---- 204=>x"8100", 205=>x"8100", 206=>x"8000", 207=>x"7d00", 208=>x"7d00", 209=>x"7d00", 210=>x"7f00",
---- 211=>x"7f00", 212=>x"7d00", 213=>x"7f00", 214=>x"7f00", 215=>x"7e00", 216=>x"7800", 217=>x"7b00",
---- 218=>x"7c00", 219=>x"7e00", 220=>x"7d00", 221=>x"7f00", 222=>x"7f00", 223=>x"8100", 224=>x"7500",
---- 225=>x"7600", 226=>x"7e00", 227=>x"7c00", 228=>x"7e00", 229=>x"8100", 230=>x"7f00", 231=>x"7e00",
---- 232=>x"6c00", 233=>x"7600", 234=>x"7c00", 235=>x"7900", 236=>x"7a00", 237=>x"7d00", 238=>x"8000",
---- 239=>x"7b00", 240=>x"7800", 241=>x"6c00", 242=>x"8800", 243=>x"7300", 244=>x"7600", 245=>x"7500",
---- 246=>x"7700", 247=>x"7900", 248=>x"b800", 249=>x"8f00", 250=>x"7000", 251=>x"6d00", 252=>x"7100",
---- 253=>x"7100", 254=>x"7600", 255=>x"7800", 256=>x"c900", 257=>x"c400", 258=>x"9f00", 259=>x"7400",
---- 260=>x"6a00", 261=>x"6d00", 262=>x"7200", 263=>x"7200", 264=>x"c300", 265=>x"c100", 266=>x"c500",
---- 267=>x"b500", 268=>x"8500", 269=>x"9700", 270=>x"6700", 271=>x"6b00", 272=>x"c100", 273=>x"c300",
---- 274=>x"c200", 275=>x"c900", 276=>x"c300", 277=>x"9e00", 278=>x"6c00", 279=>x"6300", 280=>x"c300",
---- 281=>x"c500", 282=>x"c600", 283=>x"c900", 284=>x"cc00", 285=>x"ca00", 286=>x"ab00", 287=>x"7200",
---- 288=>x"c300", 289=>x"c300", 290=>x"c500", 291=>x"ca00", 292=>x"ca00", 293=>x"ca00", 294=>x"d000",
---- 295=>x"b100", 296=>x"c300", 297=>x"c600", 298=>x"c800", 299=>x"c600", 300=>x"c400", 301=>x"c100",
---- 302=>x"c400", 303=>x"cc00", 304=>x"c100", 305=>x"c100", 306=>x"bc00", 307=>x"b800", 308=>x"bc00",
---- 309=>x"c100", 310=>x"cb00", 311=>x"d500", 312=>x"b800", 313=>x"bc00", 314=>x"be00", 315=>x"cb00",
---- 316=>x"d300", 317=>x"d700", 318=>x"d900", 319=>x"db00", 320=>x"c500", 321=>x"d100", 322=>x"d400",
---- 323=>x"d400", 324=>x"d800", 325=>x"d600", 326=>x"d500", 327=>x"d700", 328=>x"d800", 329=>x"d300",
---- 330=>x"d300", 331=>x"d200", 332=>x"d200", 333=>x"d600", 334=>x"d200", 335=>x"d300", 336=>x"d300",
---- 337=>x"cf00", 338=>x"cf00", 339=>x"d300", 340=>x"d000", 341=>x"d200", 342=>x"d300", 343=>x"ce00",
---- 344=>x"ce00", 345=>x"d000", 346=>x"d100", 347=>x"cf00", 348=>x"cf00", 349=>x"cd00", 350=>x"d200",
---- 351=>x"d500", 352=>x"d000", 353=>x"ce00", 354=>x"cf00", 355=>x"d000", 356=>x"3200", 357=>x"cf00",
---- 358=>x"cf00", 359=>x"d200", 360=>x"ce00", 361=>x"d100", 362=>x"ce00", 363=>x"cf00", 364=>x"ce00",
---- 365=>x"cb00", 366=>x"cf00", 367=>x"3200", 368=>x"c900", 369=>x"cf00", 370=>x"ce00", 371=>x"cb00",
---- 372=>x"cc00", 373=>x"ca00", 374=>x"ca00", 375=>x"cf00", 376=>x"c500", 377=>x"c100", 378=>x"c400",
---- 379=>x"cb00", 380=>x"ca00", 381=>x"ce00", 382=>x"d600", 383=>x"d900", 384=>x"ca00", 385=>x"c700",
---- 386=>x"c700", 387=>x"cf00", 388=>x"d100", 389=>x"cb00", 390=>x"cf00", 391=>x"ce00", 392=>x"2e00",
---- 393=>x"d100", 394=>x"c900", 395=>x"c700", 396=>x"c800", 397=>x"c500", 398=>x"c700", 399=>x"c800",
---- 400=>x"c700", 401=>x"c800", 402=>x"c900", 403=>x"ca00", 404=>x"c900", 405=>x"cb00", 406=>x"d000",
---- 407=>x"cd00", 408=>x"cd00", 409=>x"c400", 410=>x"cb00", 411=>x"d300", 412=>x"cf00", 413=>x"ce00",
---- 414=>x"cd00", 415=>x"cf00", 416=>x"ce00", 417=>x"d100", 418=>x"c500", 419=>x"cd00", 420=>x"d200",
---- 421=>x"cf00", 422=>x"cf00", 423=>x"cf00", 424=>x"c500", 425=>x"ce00", 426=>x"d100", 427=>x"c800",
---- 428=>x"ce00", 429=>x"cd00", 430=>x"d000", 431=>x"cc00", 432=>x"cd00", 433=>x"c800", 434=>x"d400",
---- 435=>x"ce00", 436=>x"c300", 437=>x"cf00", 438=>x"d000", 439=>x"cf00", 440=>x"cf00", 441=>x"ca00",
---- 442=>x"c900", 443=>x"d100", 444=>x"c800", 445=>x"cc00", 446=>x"cd00", 447=>x"cc00", 448=>x"cd00",
---- 449=>x"cc00", 450=>x"c600", 451=>x"3300", 452=>x"ce00", 453=>x"ca00", 454=>x"cd00", 455=>x"cf00",
---- 456=>x"cd00", 457=>x"ca00", 458=>x"c800", 459=>x"cc00", 460=>x"ca00", 461=>x"cc00", 462=>x"c700",
---- 463=>x"c600", 464=>x"ca00", 465=>x"ce00", 466=>x"c700", 467=>x"c500", 468=>x"c400", 469=>x"c100",
---- 470=>x"ca00", 471=>x"cb00", 472=>x"c700", 473=>x"c800", 474=>x"bf00", 475=>x"be00", 476=>x"c400",
---- 477=>x"c800", 478=>x"ce00", 479=>x"cf00", 480=>x"bf00", 481=>x"bb00", 482=>x"c200", 483=>x"cb00",
---- 484=>x"cc00", 485=>x"ca00", 486=>x"ca00", 487=>x"cd00", 488=>x"be00", 489=>x"c700", 490=>x"c900",
---- 491=>x"cb00", 492=>x"cc00", 493=>x"c800", 494=>x"ca00", 495=>x"cc00", 496=>x"c400", 497=>x"c900",
---- 498=>x"c800", 499=>x"c300", 500=>x"c500", 501=>x"3900", 502=>x"cb00", 503=>x"cb00", 504=>x"c400",
---- 505=>x"c400", 506=>x"c600", 507=>x"c500", 508=>x"c000", 509=>x"bb00", 510=>x"c400", 511=>x"cb00",
---- 512=>x"c900", 513=>x"c200", 514=>x"c000", 515=>x"c800", 516=>x"c800", 517=>x"c100", 518=>x"bc00",
---- 519=>x"c700", 520=>x"c800", 521=>x"c500", 522=>x"bd00", 523=>x"c100", 524=>x"c500", 525=>x"c700",
---- 526=>x"c300", 527=>x"c000", 528=>x"c300", 529=>x"c600", 530=>x"c600", 531=>x"c300", 532=>x"c300",
---- 533=>x"c300", 534=>x"c400", 535=>x"c900", 536=>x"c000", 537=>x"c600", 538=>x"c500", 539=>x"c100",
---- 540=>x"c500", 541=>x"c900", 542=>x"c500", 543=>x"c600", 544=>x"c100", 545=>x"bc00", 546=>x"c200",
---- 547=>x"be00", 548=>x"c000", 549=>x"ca00", 550=>x"c800", 551=>x"c600", 552=>x"b600", 553=>x"c000",
---- 554=>x"be00", 555=>x"c000", 556=>x"be00", 557=>x"c700", 558=>x"3200", 559=>x"cd00", 560=>x"ac00",
---- 561=>x"b400", 562=>x"c100", 563=>x"c600", 564=>x"c300", 565=>x"be00", 566=>x"c400", 567=>x"be00",
---- 568=>x"ba00", 569=>x"b400", 570=>x"bd00", 571=>x"b900", 572=>x"b200", 573=>x"a200", 574=>x"ab00",
---- 575=>x"ad00", 576=>x"bf00", 577=>x"bc00", 578=>x"c100", 579=>x"b000", 580=>x"a100", 581=>x"ae00",
---- 582=>x"ba00", 583=>x"b800", 584=>x"c100", 585=>x"bc00", 586=>x"b400", 587=>x"af00", 588=>x"b300",
---- 589=>x"b400", 590=>x"b600", 591=>x"b900", 592=>x"b700", 593=>x"b000", 594=>x"b200", 595=>x"b800",
---- 596=>x"b700", 597=>x"b600", 598=>x"b900", 599=>x"b300", 600=>x"af00", 601=>x"b900", 602=>x"bc00",
---- 603=>x"b700", 604=>x"b200", 605=>x"b400", 606=>x"b800", 607=>x"ad00", 608=>x"b300", 609=>x"b600",
---- 610=>x"ba00", 611=>x"b800", 612=>x"b000", 613=>x"b200", 614=>x"b800", 615=>x"b700", 616=>x"b200",
---- 617=>x"b300", 618=>x"a900", 619=>x"a800", 620=>x"af00", 621=>x"b200", 622=>x"b700", 623=>x"bc00",
---- 624=>x"a400", 625=>x"a100", 626=>x"ab00", 627=>x"aa00", 628=>x"b000", 629=>x"b200", 630=>x"b000",
---- 631=>x"ba00", 632=>x"a100", 633=>x"a900", 634=>x"af00", 635=>x"af00", 636=>x"ac00", 637=>x"af00",
---- 638=>x"ae00", 639=>x"ae00", 640=>x"a900", 641=>x"a900", 642=>x"a800", 643=>x"af00", 644=>x"b000",
---- 645=>x"ad00", 646=>x"a700", 647=>x"a900", 648=>x"a500", 649=>x"aa00", 650=>x"aa00", 651=>x"a700",
---- 652=>x"b100", 653=>x"a900", 654=>x"a300", 655=>x"ab00", 656=>x"a300", 657=>x"9f00", 658=>x"aa00",
---- 659=>x"aa00", 660=>x"ac00", 661=>x"ab00", 662=>x"a400", 663=>x"a400", 664=>x"ab00", 665=>x"a400",
---- 666=>x"a100", 667=>x"a700", 668=>x"a600", 669=>x"a600", 670=>x"a600", 671=>x"a800", 672=>x"a400",
---- 673=>x"a900", 674=>x"a500", 675=>x"9d00", 676=>x"a700", 677=>x"a200", 678=>x"a600", 679=>x"a600",
---- 680=>x"a100", 681=>x"a400", 682=>x"a600", 683=>x"9c00", 684=>x"9e00", 685=>x"a300", 686=>x"a100",
---- 687=>x"a500", 688=>x"9b00", 689=>x"a500", 690=>x"a300", 691=>x"a300", 692=>x"9600", 693=>x"8f00",
---- 694=>x"8700", 695=>x"6700", 696=>x"7400", 697=>x"8d00", 698=>x"9300", 699=>x"9500", 700=>x"a600",
---- 701=>x"7a00", 702=>x"7a00", 703=>x"5000", 704=>x"7e00", 705=>x"6a00", 706=>x"6b00", 707=>x"5200",
---- 708=>x"6700", 709=>x"4f00", 710=>x"6700", 711=>x"7500", 712=>x"5000", 713=>x"4d00", 714=>x"4a00",
---- 715=>x"3800", 716=>x"2900", 717=>x"3400", 718=>x"2c00", 719=>x"3c00", 720=>x"3500", 721=>x"3300",
---- 722=>x"3400", 723=>x"3000", 724=>x"2b00", 725=>x"2f00", 726=>x"2d00", 727=>x"2200", 728=>x"3400",
---- 729=>x"2b00", 730=>x"2900", 731=>x"2200", 732=>x"2d00", 733=>x"3700", 734=>x"2600", 735=>x"4f00",
---- 736=>x"3800", 737=>x"3300", 738=>x"2800", 739=>x"2200", 740=>x"2300", 741=>x"1e00", 742=>x"3300",
---- 743=>x"9600", 744=>x"2b00", 745=>x"2a00", 746=>x"2c00", 747=>x"2300", 748=>x"1d00", 749=>x"4000",
---- 750=>x"9100", 751=>x"ba00", 752=>x"2300", 753=>x"2100", 754=>x"2100", 755=>x"2d00", 756=>x"5600",
---- 757=>x"a600", 758=>x"b900", 759=>x"8400", 760=>x"1e00", 761=>x"1f00", 762=>x"1e00", 763=>x"5c00",
---- 764=>x"ac00", 765=>x"b000", 766=>x"8100", 767=>x"7400", 768=>x"2c00", 769=>x"2200", 770=>x"9b00",
---- 771=>x"ae00", 772=>x"a400", 773=>x"7b00", 774=>x"8300", 775=>x"ad00", 776=>x"4000", 777=>x"7300",
---- 778=>x"b200", 779=>x"9b00", 780=>x"7600", 781=>x"8700", 782=>x"b500", 783=>x"c700", 784=>x"8100",
---- 785=>x"b100", 786=>x"9500", 787=>x"7500", 788=>x"8e00", 789=>x"b100", 790=>x"c400", 791=>x"c700",
---- 792=>x"a900", 793=>x"8800", 794=>x"7500", 795=>x"8f00", 796=>x"bd00", 797=>x"be00", 798=>x"c300",
---- 799=>x"c700", 800=>x"7b00", 801=>x"7000", 802=>x"9100", 803=>x"bb00", 804=>x"c800", 805=>x"c200",
---- 806=>x"c000", 807=>x"c100", 808=>x"7700", 809=>x"9a00", 810=>x"bd00", 811=>x"c400", 812=>x"c600",
---- 813=>x"c200", 814=>x"bf00", 815=>x"be00", 816=>x"a400", 817=>x"c200", 818=>x"c600", 819=>x"c200",
---- 820=>x"c200", 821=>x"c100", 822=>x"be00", 823=>x"bb00", 824=>x"c100", 825=>x"bf00", 826=>x"c300",
---- 827=>x"c100", 828=>x"c100", 829=>x"c100", 830=>x"b900", 831=>x"b800", 832=>x"bb00", 833=>x"be00",
---- 834=>x"bd00", 835=>x"ba00", 836=>x"bf00", 837=>x"bc00", 838=>x"ba00", 839=>x"b700", 840=>x"ba00",
---- 841=>x"b700", 842=>x"b300", 843=>x"b800", 844=>x"bb00", 845=>x"b800", 846=>x"b500", 847=>x"af00",
---- 848=>x"b600", 849=>x"ae00", 850=>x"5000", 851=>x"b500", 852=>x"b600", 853=>x"b300", 854=>x"ac00",
---- 855=>x"ab00", 856=>x"b200", 857=>x"b000", 858=>x"b600", 859=>x"b900", 860=>x"b300", 861=>x"ad00",
---- 862=>x"ab00", 863=>x"a800", 864=>x"b400", 865=>x"b900", 866=>x"bd00", 867=>x"b900", 868=>x"b300",
---- 869=>x"aa00", 870=>x"a300", 871=>x"a500", 872=>x"ba00", 873=>x"bc00", 874=>x"bb00", 875=>x"b400",
---- 876=>x"ac00", 877=>x"a300", 878=>x"5f00", 879=>x"a500", 880=>x"bf00", 881=>x"c300", 882=>x"bb00",
---- 883=>x"af00", 884=>x"5900", 885=>x"a200", 886=>x"9e00", 887=>x"a300", 888=>x"bf00", 889=>x"bc00",
---- 890=>x"b300", 891=>x"a800", 892=>x"a400", 893=>x"a200", 894=>x"a000", 895=>x"a100", 896=>x"b500",
---- 897=>x"b200", 898=>x"b100", 899=>x"a900", 900=>x"a800", 901=>x"a500", 902=>x"a400", 903=>x"a700",
---- 904=>x"ba00", 905=>x"b600", 906=>x"ab00", 907=>x"aa00", 908=>x"aa00", 909=>x"ab00", 910=>x"aa00",
---- 911=>x"ae00", 912=>x"c200", 913=>x"b500", 914=>x"a800", 915=>x"a900", 916=>x"ab00", 917=>x"aa00",
---- 918=>x"a900", 919=>x"9e00", 920=>x"c500", 921=>x"b100", 922=>x"a700", 923=>x"ac00", 924=>x"a600",
---- 925=>x"a300", 926=>x"9b00", 927=>x"9400", 928=>x"bc00", 929=>x"a900", 930=>x"a400", 931=>x"a400",
---- 932=>x"a500", 933=>x"9b00", 934=>x"9700", 935=>x"9e00", 936=>x"ae00", 937=>x"a200", 938=>x"9d00",
---- 939=>x"a400", 940=>x"9c00", 941=>x"9b00", 942=>x"a100", 943=>x"a100", 944=>x"a200", 945=>x"9b00",
---- 946=>x"9800", 947=>x"9c00", 948=>x"9a00", 949=>x"9d00", 950=>x"a200", 951=>x"a200", 952=>x"9e00",
---- 953=>x"9a00", 954=>x"9c00", 955=>x"a300", 956=>x"a200", 957=>x"9f00", 958=>x"a300", 959=>x"a500",
---- 960=>x"9a00", 961=>x"9e00", 962=>x"a600", 963=>x"a600", 964=>x"a400", 965=>x"a300", 966=>x"a500",
---- 967=>x"a700", 968=>x"9200", 969=>x"9a00", 970=>x"9d00", 971=>x"a300", 972=>x"a600", 973=>x"a600",
---- 974=>x"aa00", 975=>x"aa00", 976=>x"7600", 977=>x"8200", 978=>x"8e00", 979=>x"9400", 980=>x"9800",
---- 981=>x"9d00", 982=>x"a700", 983=>x"ac00", 984=>x"5f00", 985=>x"6600", 986=>x"6100", 987=>x"6500",
---- 988=>x"7400", 989=>x"8000", 990=>x"9100", 991=>x"a200", 992=>x"7400", 993=>x"6c00", 994=>x"5900",
---- 995=>x"4400", 996=>x"4300", 997=>x"4c00", 998=>x"5b00", 999=>x"7100", 1000=>x"9a00", 1001=>x"8d00",
---- 1002=>x"7800", 1003=>x"6300", 1004=>x"4e00", 1005=>x"4700", 1006=>x"4000", 1007=>x"4000", 1008=>x"a500",
---- 1009=>x"9b00", 1010=>x"8400", 1011=>x"7800", 1012=>x"6900", 1013=>x"5f00", 1014=>x"5800", 1015=>x"4d00",
---- 1016=>x"9a00", 1017=>x"8800", 1018=>x"6800", 1019=>x"7400", 1020=>x"6100", 1021=>x"7500", 1022=>x"6d00",
---- 1023=>x"6600", 1024=>x"6300", 1025=>x"4d00", 1026=>x"cb00", 1027=>x"4400", 1028=>x"5200", 1029=>x"7d00",
---- 1030=>x"6700", 1031=>x"7600", 1032=>x"2e00", 1033=>x"2d00", 1034=>x"2c00", 1035=>x"2700", 1036=>x"2d00",
---- 1037=>x"4500", 1038=>x"6a00", 1039=>x"8e00", 1040=>x"4500", 1041=>x"4c00", 1042=>x"3300", 1043=>x"2a00",
---- 1044=>x"2b00", 1045=>x"2700", 1046=>x"3f00", 1047=>x"7200", 1048=>x"8800", 1049=>x"9e00", 1050=>x"6b00",
---- 1051=>x"3900", 1052=>x"2700", 1053=>x"2900", 1054=>x"2300", 1055=>x"4000", 1056=>x"a800", 1057=>x"cf00",
---- 1058=>x"b300", 1059=>x"8d00", 1060=>x"4300", 1061=>x"2b00", 1062=>x"4800", 1063=>x"4200", 1064=>x"9400",
---- 1065=>x"d200", 1066=>x"c700", 1067=>x"c500", 1068=>x"8d00", 1069=>x"4600", 1070=>x"6400", 1071=>x"6c00",
---- 1072=>x"ba00", 1073=>x"d400", 1074=>x"cf00", 1075=>x"cc00", 1076=>x"b800", 1077=>x"6900", 1078=>x"4f00",
---- 1079=>x"7700", 1080=>x"d100", 1081=>x"ce00", 1082=>x"ce00", 1083=>x"c900", 1084=>x"b200", 1085=>x"8500",
---- 1086=>x"6300", 1087=>x"7600", 1088=>x"c900", 1089=>x"ce00", 1090=>x"cf00", 1091=>x"be00", 1092=>x"6b00",
---- 1093=>x"8e00", 1094=>x"8600", 1095=>x"6f00", 1096=>x"be00", 1097=>x"c500", 1098=>x"be00", 1099=>x"b200",
---- 1100=>x"9e00", 1101=>x"9100", 1102=>x"8500", 1103=>x"7a00", 1104=>x"9200", 1105=>x"9400", 1106=>x"9600",
---- 1107=>x"ae00", 1108=>x"b100", 1109=>x"ad00", 1110=>x"a600", 1111=>x"9200", 1112=>x"6f00", 1113=>x"7200",
---- 1114=>x"8100", 1115=>x"9d00", 1116=>x"9b00", 1117=>x"a700", 1118=>x"9e00", 1119=>x"8b00", 1120=>x"8100",
---- 1121=>x"9000", 1122=>x"9400", 1123=>x"9b00", 1124=>x"9700", 1125=>x"9300", 1126=>x"9200", 1127=>x"9300",
---- 1128=>x"9800", 1129=>x"9a00", 1130=>x"a100", 1131=>x"a200", 1132=>x"a200", 1133=>x"9b00", 1134=>x"a400",
---- 1135=>x"9800", 1136=>x"a200", 1137=>x"a800", 1138=>x"a800", 1139=>x"a600", 1140=>x"a300", 1141=>x"a500",
---- 1142=>x"a500", 1143=>x"9000", 1144=>x"ab00", 1145=>x"ad00", 1146=>x"a400", 1147=>x"aa00", 1148=>x"a700",
---- 1149=>x"a800", 1150=>x"9e00", 1151=>x"8d00", 1152=>x"aa00", 1153=>x"a600", 1154=>x"a900", 1155=>x"a900",
---- 1156=>x"a800", 1157=>x"a100", 1158=>x"9a00", 1159=>x"8e00", 1160=>x"a700", 1161=>x"af00", 1162=>x"b000",
---- 1163=>x"af00", 1164=>x"a800", 1165=>x"9d00", 1166=>x"9800", 1167=>x"9400", 1168=>x"ad00", 1169=>x"af00",
---- 1170=>x"b100", 1171=>x"ad00", 1172=>x"a800", 1173=>x"a300", 1174=>x"9900", 1175=>x"9200", 1176=>x"b100",
---- 1177=>x"b200", 1178=>x"b000", 1179=>x"aa00", 1180=>x"a500", 1181=>x"a000", 1182=>x"9b00", 1183=>x"9600",
---- 1184=>x"af00", 1185=>x"b000", 1186=>x"aa00", 1187=>x"a900", 1188=>x"a400", 1189=>x"9f00", 1190=>x"9900",
---- 1191=>x"9600", 1192=>x"ab00", 1193=>x"ac00", 1194=>x"ab00", 1195=>x"a700", 1196=>x"a000", 1197=>x"9d00",
---- 1198=>x"9900", 1199=>x"9300", 1200=>x"ad00", 1201=>x"ae00", 1202=>x"a800", 1203=>x"a400", 1204=>x"a000",
---- 1205=>x"9b00", 1206=>x"9100", 1207=>x"8e00", 1208=>x"aa00", 1209=>x"ab00", 1210=>x"a800", 1211=>x"a300",
---- 1212=>x"9f00", 1213=>x"9a00", 1214=>x"9200", 1215=>x"8f00", 1216=>x"aa00", 1217=>x"a900", 1218=>x"a600",
---- 1219=>x"a300", 1220=>x"9d00", 1221=>x"9600", 1222=>x"9200", 1223=>x"8800", 1224=>x"aa00", 1225=>x"a800",
---- 1226=>x"a400", 1227=>x"a300", 1228=>x"9b00", 1229=>x"9800", 1230=>x"8e00", 1231=>x"8500", 1232=>x"a900",
---- 1233=>x"a600", 1234=>x"a300", 1235=>x"a000", 1236=>x"9b00", 1237=>x"9700", 1238=>x"8c00", 1239=>x"8600",
---- 1240=>x"a500", 1241=>x"a400", 1242=>x"5b00", 1243=>x"a100", 1244=>x"9b00", 1245=>x"9400", 1246=>x"8c00",
---- 1247=>x"8600", 1248=>x"a000", 1249=>x"a300", 1250=>x"a100", 1251=>x"9e00", 1252=>x"9700", 1253=>x"9000",
---- 1254=>x"8900", 1255=>x"8100", 1256=>x"5b00", 1257=>x"a200", 1258=>x"9d00", 1259=>x"6600", 1260=>x"9400",
---- 1261=>x"9000", 1262=>x"8900", 1263=>x"7b00", 1264=>x"a100", 1265=>x"a100", 1266=>x"9c00", 1267=>x"9800",
---- 1268=>x"9200", 1269=>x"8f00", 1270=>x"8100", 1271=>x"7100", 1272=>x"9e00", 1273=>x"9e00", 1274=>x"9e00",
---- 1275=>x"9400", 1276=>x"6e00", 1277=>x"8f00", 1278=>x"7f00", 1279=>x"6b00", 1280=>x"9f00", 1281=>x"9f00",
---- 1282=>x"9c00", 1283=>x"9700", 1284=>x"9200", 1285=>x"9100", 1286=>x"8100", 1287=>x"6c00", 1288=>x"9e00",
---- 1289=>x"9c00", 1290=>x"9d00", 1291=>x"9a00", 1292=>x"9200", 1293=>x"8e00", 1294=>x"8500", 1295=>x"7500",
---- 1296=>x"9e00", 1297=>x"9d00", 1298=>x"9f00", 1299=>x"9800", 1300=>x"9500", 1301=>x"9300", 1302=>x"8b00",
---- 1303=>x"7a00", 1304=>x"9f00", 1305=>x"9c00", 1306=>x"9d00", 1307=>x"9c00", 1308=>x"9500", 1309=>x"9400",
---- 1310=>x"9200", 1311=>x"8400", 1312=>x"9e00", 1313=>x"6000", 1314=>x"9d00", 1315=>x"9d00", 1316=>x"9800",
---- 1317=>x"9500", 1318=>x"9400", 1319=>x"8e00", 1320=>x"9b00", 1321=>x"9f00", 1322=>x"9f00", 1323=>x"9c00",
---- 1324=>x"9b00", 1325=>x"9a00", 1326=>x"9700", 1327=>x"9400", 1328=>x"a000", 1329=>x"9f00", 1330=>x"9d00",
---- 1331=>x"9e00", 1332=>x"9b00", 1333=>x"9e00", 1334=>x"9900", 1335=>x"9500", 1336=>x"9d00", 1337=>x"9f00",
---- 1338=>x"9d00", 1339=>x"9d00", 1340=>x"9a00", 1341=>x"9600", 1342=>x"9900", 1343=>x"9600", 1344=>x"9600",
---- 1345=>x"9a00", 1346=>x"9a00", 1347=>x"9c00", 1348=>x"9900", 1349=>x"9500", 1350=>x"9600", 1351=>x"9700",
---- 1352=>x"9400", 1353=>x"9900", 1354=>x"9800", 1355=>x"9a00", 1356=>x"9a00", 1357=>x"9200", 1358=>x"9100",
---- 1359=>x"9600", 1360=>x"9400", 1361=>x"9400", 1362=>x"9400", 1363=>x"9a00", 1364=>x"9600", 1365=>x"9600",
---- 1366=>x"9200", 1367=>x"9300", 1368=>x"9100", 1369=>x"9100", 1370=>x"8f00", 1371=>x"9400", 1372=>x"9100",
---- 1373=>x"9100", 1374=>x"9200", 1375=>x"9200", 1376=>x"9000", 1377=>x"8f00", 1378=>x"8c00", 1379=>x"8f00",
---- 1380=>x"9100", 1381=>x"8f00", 1382=>x"8f00", 1383=>x"7000", 1384=>x"8700", 1385=>x"8700", 1386=>x"8900",
---- 1387=>x"8e00", 1388=>x"8e00", 1389=>x"8f00", 1390=>x"8f00", 1391=>x"9000", 1392=>x"7a00", 1393=>x"7f00",
---- 1394=>x"8400", 1395=>x"8900", 1396=>x"8600", 1397=>x"8400", 1398=>x"8300", 1399=>x"7f00", 1400=>x"5200",
---- 1401=>x"5900", 1402=>x"6300", 1403=>x"6800", 1404=>x"9500", 1405=>x"6900", 1406=>x"7000", 1407=>x"6a00",
---- 1408=>x"6700", 1409=>x"5e00", 1410=>x"5b00", 1411=>x"6000", 1412=>x"6600", 1413=>x"6b00", 1414=>x"7300",
---- 1415=>x"7000", 1416=>x"7f00", 1417=>x"7d00", 1418=>x"7c00", 1419=>x"7900", 1420=>x"7900", 1421=>x"7d00",
---- 1422=>x"8400", 1423=>x"8700", 1424=>x"7c00", 1425=>x"7f00", 1426=>x"7f00", 1427=>x"8100", 1428=>x"7900",
---- 1429=>x"7900", 1430=>x"7f00", 1431=>x"8600", 1432=>x"8000", 1433=>x"7d00", 1434=>x"8600", 1435=>x"8000",
---- 1436=>x"8000", 1437=>x"7f00", 1438=>x"7f00", 1439=>x"7e00", 1440=>x"8500", 1441=>x"8400", 1442=>x"7c00",
---- 1443=>x"7a00", 1444=>x"7b00", 1445=>x"8100", 1446=>x"8300", 1447=>x"8000", 1448=>x"8600", 1449=>x"8400",
---- 1450=>x"8300", 1451=>x"7e00", 1452=>x"7e00", 1453=>x"7c00", 1454=>x"7b00", 1455=>x"7c00", 1456=>x"8700",
---- 1457=>x"8500", 1458=>x"8500", 1459=>x"8200", 1460=>x"8500", 1461=>x"8000", 1462=>x"7c00", 1463=>x"7700",
---- 1464=>x"8900", 1465=>x"8700", 1466=>x"8500", 1467=>x"8100", 1468=>x"8400", 1469=>x"8000", 1470=>x"8200",
---- 1471=>x"8300", 1472=>x"8800", 1473=>x"8900", 1474=>x"8700", 1475=>x"8800", 1476=>x"8700", 1477=>x"8500",
---- 1478=>x"8900", 1479=>x"8e00", 1480=>x"8b00", 1481=>x"8c00", 1482=>x"8900", 1483=>x"8b00", 1484=>x"8e00",
---- 1485=>x"8d00", 1486=>x"9500", 1487=>x"9900", 1488=>x"8b00", 1489=>x"8e00", 1490=>x"9300", 1491=>x"9700",
---- 1492=>x"9700", 1493=>x"9300", 1494=>x"9500", 1495=>x"9b00", 1496=>x"8d00", 1497=>x"9300", 1498=>x"9500",
---- 1499=>x"9c00", 1500=>x"9f00", 1501=>x"9c00", 1502=>x"9900", 1503=>x"a000", 1504=>x"9000", 1505=>x"9600",
---- 1506=>x"9800", 1507=>x"a000", 1508=>x"a600", 1509=>x"a700", 1510=>x"a300", 1511=>x"a200", 1512=>x"9100",
---- 1513=>x"9400", 1514=>x"9a00", 1515=>x"9c00", 1516=>x"5900", 1517=>x"ac00", 1518=>x"a800", 1519=>x"a600",
---- 1520=>x"9100", 1521=>x"9300", 1522=>x"9600", 1523=>x"9600", 1524=>x"9e00", 1525=>x"a700", 1526=>x"a400",
---- 1527=>x"a700", 1528=>x"8e00", 1529=>x"9200", 1530=>x"9300", 1531=>x"9400", 1532=>x"9c00", 1533=>x"9c00",
---- 1534=>x"a200", 1535=>x"a800", 1536=>x"8400", 1537=>x"7700", 1538=>x"8d00", 1539=>x"9400", 1540=>x"9900",
---- 1541=>x"6b00", 1542=>x"9900", 1543=>x"a300", 1544=>x"8000", 1545=>x"8700", 1546=>x"8700", 1547=>x"9000",
---- 1548=>x"9600", 1549=>x"9400", 1550=>x"9700", 1551=>x"9d00", 1552=>x"8700", 1553=>x"9200", 1554=>x"8e00",
---- 1555=>x"9d00", 1556=>x"9e00", 1557=>x"a100", 1558=>x"a000", 1559=>x"a000", 1560=>x"8c00", 1561=>x"8d00",
---- 1562=>x"9100", 1563=>x"9900", 1564=>x"9b00", 1565=>x"9e00", 1566=>x"9a00", 1567=>x"9900", 1568=>x"8d00",
---- 1569=>x"8e00", 1570=>x"9300", 1571=>x"9600", 1572=>x"9400", 1573=>x"9900", 1574=>x"9700", 1575=>x"9600",
---- 1576=>x"8a00", 1577=>x"8c00", 1578=>x"9100", 1579=>x"9300", 1580=>x"9500", 1581=>x"9300", 1582=>x"9200",
---- 1583=>x"9100", 1584=>x"8a00", 1585=>x"8c00", 1586=>x"8e00", 1587=>x"6b00", 1588=>x"9100", 1589=>x"8d00",
---- 1590=>x"8f00", 1591=>x"8d00", 1592=>x"7300", 1593=>x"8b00", 1594=>x"8d00", 1595=>x"8e00", 1596=>x"8c00",
---- 1597=>x"8c00", 1598=>x"8d00", 1599=>x"8c00", 1600=>x"8700", 1601=>x"8b00", 1602=>x"8d00", 1603=>x"8b00",
---- 1604=>x"8e00", 1605=>x"8d00", 1606=>x"8900", 1607=>x"8d00", 1608=>x"8a00", 1609=>x"8d00", 1610=>x"8c00",
---- 1611=>x"8b00", 1612=>x"8d00", 1613=>x"8a00", 1614=>x"8a00", 1615=>x"9000", 1616=>x"8d00", 1617=>x"8f00",
---- 1618=>x"8c00", 1619=>x"7500", 1620=>x"8c00", 1621=>x"8900", 1622=>x"8b00", 1623=>x"9100", 1624=>x"8e00",
---- 1625=>x"8c00", 1626=>x"8d00", 1627=>x"8800", 1628=>x"8700", 1629=>x"8700", 1630=>x"8b00", 1631=>x"9100",
---- 1632=>x"8c00", 1633=>x"8d00", 1634=>x"8e00", 1635=>x"8900", 1636=>x"8800", 1637=>x"8a00", 1638=>x"8c00",
---- 1639=>x"9000", 1640=>x"8900", 1641=>x"8d00", 1642=>x"8d00", 1643=>x"8900", 1644=>x"8a00", 1645=>x"8d00",
---- 1646=>x"8e00", 1647=>x"9300", 1648=>x"8e00", 1649=>x"8c00", 1650=>x"8900", 1651=>x"8d00", 1652=>x"8a00",
---- 1653=>x"8f00", 1654=>x"9400", 1655=>x"9600", 1656=>x"9000", 1657=>x"8a00", 1658=>x"7100", 1659=>x"8c00",
---- 1660=>x"8c00", 1661=>x"8f00", 1662=>x"6a00", 1663=>x"9600", 1664=>x"8900", 1665=>x"8b00", 1666=>x"8c00",
---- 1667=>x"8b00", 1668=>x"9100", 1669=>x"8f00", 1670=>x"9200", 1671=>x"9500", 1672=>x"8b00", 1673=>x"8b00",
---- 1674=>x"8a00", 1675=>x"8f00", 1676=>x"8f00", 1677=>x"9100", 1678=>x"9100", 1679=>x"9400", 1680=>x"8d00",
---- 1681=>x"8d00", 1682=>x"8c00", 1683=>x"8c00", 1684=>x"8e00", 1685=>x"8f00", 1686=>x"9200", 1687=>x"9700",
---- 1688=>x"8c00", 1689=>x"8d00", 1690=>x"8d00", 1691=>x"8f00", 1692=>x"8d00", 1693=>x"9000", 1694=>x"9200",
---- 1695=>x"9600", 1696=>x"7100", 1697=>x"8e00", 1698=>x"8d00", 1699=>x"8d00", 1700=>x"9100", 1701=>x"9400",
---- 1702=>x"9500", 1703=>x"9700", 1704=>x"8b00", 1705=>x"8c00", 1706=>x"8d00", 1707=>x"8e00", 1708=>x"9100",
---- 1709=>x"9500", 1710=>x"9400", 1711=>x"9100", 1712=>x"8b00", 1713=>x"8d00", 1714=>x"8d00", 1715=>x"8e00",
---- 1716=>x"8f00", 1717=>x"8f00", 1718=>x"9400", 1719=>x"9000", 1720=>x"8a00", 1721=>x"8c00", 1722=>x"8a00",
---- 1723=>x"8d00", 1724=>x"8d00", 1725=>x"9100", 1726=>x"9200", 1727=>x"8f00", 1728=>x"8800", 1729=>x"8a00",
---- 1730=>x"8800", 1731=>x"8c00", 1732=>x"8f00", 1733=>x"9100", 1734=>x"9100", 1735=>x"9300", 1736=>x"8800",
---- 1737=>x"8700", 1738=>x"8900", 1739=>x"8b00", 1740=>x"9000", 1741=>x"9000", 1742=>x"9200", 1743=>x"9000",
---- 1744=>x"8800", 1745=>x"8a00", 1746=>x"8a00", 1747=>x"8a00", 1748=>x"8d00", 1749=>x"8d00", 1750=>x"9000",
---- 1751=>x"9000", 1752=>x"8a00", 1753=>x"8c00", 1754=>x"8c00", 1755=>x"7700", 1756=>x"8e00", 1757=>x"8f00",
---- 1758=>x"9000", 1759=>x"9000", 1760=>x"8900", 1761=>x"8800", 1762=>x"8a00", 1763=>x"8a00", 1764=>x"8c00",
---- 1765=>x"8c00", 1766=>x"8d00", 1767=>x"8d00", 1768=>x"8100", 1769=>x"8700", 1770=>x"8700", 1771=>x"8900",
---- 1772=>x"8a00", 1773=>x"8c00", 1774=>x"8d00", 1775=>x"8f00", 1776=>x"8400", 1777=>x"8600", 1778=>x"8600",
---- 1779=>x"8900", 1780=>x"8b00", 1781=>x"8a00", 1782=>x"8e00", 1783=>x"9000", 1784=>x"8700", 1785=>x"8600",
---- 1786=>x"8500", 1787=>x"8700", 1788=>x"8a00", 1789=>x"8800", 1790=>x"8c00", 1791=>x"8f00", 1792=>x"8500",
---- 1793=>x"8600", 1794=>x"8600", 1795=>x"8800", 1796=>x"8a00", 1797=>x"8b00", 1798=>x"8c00", 1799=>x"8c00",
---- 1800=>x"8700", 1801=>x"8800", 1802=>x"8700", 1803=>x"8900", 1804=>x"8a00", 1805=>x"8c00", 1806=>x"8a00",
---- 1807=>x"8b00", 1808=>x"8700", 1809=>x"8a00", 1810=>x"8500", 1811=>x"8800", 1812=>x"8c00", 1813=>x"8b00",
---- 1814=>x"8800", 1815=>x"8c00", 1816=>x"8b00", 1817=>x"8800", 1818=>x"8900", 1819=>x"8800", 1820=>x"8700",
---- 1821=>x"8800", 1822=>x"8800", 1823=>x"8a00", 1824=>x"8a00", 1825=>x"8600", 1826=>x"8900", 1827=>x"8700",
---- 1828=>x"8700", 1829=>x"8900", 1830=>x"8500", 1831=>x"8b00", 1832=>x"8c00", 1833=>x"7500", 1834=>x"8900",
---- 1835=>x"8600", 1836=>x"8a00", 1837=>x"8c00", 1838=>x"8900", 1839=>x"8c00", 1840=>x"8e00", 1841=>x"8c00",
---- 1842=>x"8900", 1843=>x"8700", 1844=>x"8900", 1845=>x"8b00", 1846=>x"8b00", 1847=>x"8c00", 1848=>x"8c00",
---- 1849=>x"8c00", 1850=>x"8700", 1851=>x"8a00", 1852=>x"8b00", 1853=>x"8700", 1854=>x"8700", 1855=>x"8800",
---- 1856=>x"8e00", 1857=>x"8c00", 1858=>x"8700", 1859=>x"8700", 1860=>x"8a00", 1861=>x"8700", 1862=>x"8800",
---- 1863=>x"8900", 1864=>x"8c00", 1865=>x"7300", 1866=>x"8800", 1867=>x"8a00", 1868=>x"8a00", 1869=>x"8700",
---- 1870=>x"8800", 1871=>x"8600", 1872=>x"8b00", 1873=>x"8e00", 1874=>x"8900", 1875=>x"8700", 1876=>x"8a00",
---- 1877=>x"8600", 1878=>x"8500", 1879=>x"8800", 1880=>x"8d00", 1881=>x"8900", 1882=>x"8b00", 1883=>x"8c00",
---- 1884=>x"8900", 1885=>x"8800", 1886=>x"8700", 1887=>x"8800", 1888=>x"9200", 1889=>x"8d00", 1890=>x"8b00",
---- 1891=>x"8d00", 1892=>x"8900", 1893=>x"8900", 1894=>x"8a00", 1895=>x"8700", 1896=>x"8e00", 1897=>x"8d00",
---- 1898=>x"7400", 1899=>x"8c00", 1900=>x"8900", 1901=>x"8800", 1902=>x"8a00", 1903=>x"8600", 1904=>x"8e00",
---- 1905=>x"8e00", 1906=>x"8e00", 1907=>x"7300", 1908=>x"8a00", 1909=>x"7500", 1910=>x"8a00", 1911=>x"8b00",
---- 1912=>x"8e00", 1913=>x"9000", 1914=>x"8e00", 1915=>x"8b00", 1916=>x"8a00", 1917=>x"8c00", 1918=>x"8b00",
---- 1919=>x"8a00", 1920=>x"9000", 1921=>x"9000", 1922=>x"8c00", 1923=>x"8c00", 1924=>x"8d00", 1925=>x"8b00",
---- 1926=>x"8a00", 1927=>x"8900", 1928=>x"8f00", 1929=>x"9200", 1930=>x"8d00", 1931=>x"8d00", 1932=>x"8f00",
---- 1933=>x"8e00", 1934=>x"7400", 1935=>x"8a00", 1936=>x"8d00", 1937=>x"9000", 1938=>x"9000", 1939=>x"8e00",
---- 1940=>x"8c00", 1941=>x"8d00", 1942=>x"8e00", 1943=>x"8a00", 1944=>x"8f00", 1945=>x"9100", 1946=>x"9100",
---- 1947=>x"8f00", 1948=>x"8f00", 1949=>x"8e00", 1950=>x"8f00", 1951=>x"8d00", 1952=>x"9100", 1953=>x"9300",
---- 1954=>x"6d00", 1955=>x"9100", 1956=>x"9100", 1957=>x"8f00", 1958=>x"9100", 1959=>x"8e00", 1960=>x"9200",
---- 1961=>x"9100", 1962=>x"9000", 1963=>x"9400", 1964=>x"9100", 1965=>x"9100", 1966=>x"8e00", 1967=>x"8d00",
---- 1968=>x"8f00", 1969=>x"9100", 1970=>x"9100", 1971=>x"9200", 1972=>x"9100", 1973=>x"9100", 1974=>x"8f00",
---- 1975=>x"8d00", 1976=>x"9100", 1977=>x"9300", 1978=>x"9200", 1979=>x"9500", 1980=>x"9100", 1981=>x"9000",
---- 1982=>x"9200", 1983=>x"8f00", 1984=>x"9100", 1985=>x"6d00", 1986=>x"9100", 1987=>x"9200", 1988=>x"9000",
---- 1989=>x"8d00", 1990=>x"9300", 1991=>x"9000", 1992=>x"8e00", 1993=>x"9200", 1994=>x"9000", 1995=>x"9100",
---- 1996=>x"9100", 1997=>x"9100", 1998=>x"9200", 1999=>x"9300", 2000=>x"8f00", 2001=>x"9100", 2002=>x"9200",
---- 2003=>x"6e00", 2004=>x"9100", 2005=>x"9000", 2006=>x"9400", 2007=>x"9200", 2008=>x"8f00", 2009=>x"9200",
---- 2010=>x"8e00", 2011=>x"8f00", 2012=>x"9500", 2013=>x"9300", 2014=>x"9400", 2015=>x"9400", 2016=>x"8f00",
---- 2017=>x"9000", 2018=>x"8f00", 2019=>x"9200", 2020=>x"9000", 2021=>x"9000", 2022=>x"9500", 2023=>x"9300",
---- 2024=>x"8f00", 2025=>x"9100", 2026=>x"9000", 2027=>x"9400", 2028=>x"9200", 2029=>x"9300", 2030=>x"8f00",
---- 2031=>x"9000", 2032=>x"9100", 2033=>x"9000", 2034=>x"9200", 2035=>x"9100", 2036=>x"9200", 2037=>x"9400",
---- 2038=>x"8c00", 2039=>x"9100", 2040=>x"8f00", 2041=>x"9100", 2042=>x"9100", 2043=>x"8f00", 2044=>x"8f00",
---- 2045=>x"9000", 2046=>x"8e00", 2047=>x"9100"),
---- 18 => (0=>x"8000", 1=>x"8200", 2=>x"8100", 3=>x"8100", 4=>x"7f00", 5=>x"7f00", 6=>x"7f00", 7=>x"8000",
---- 8=>x"8000", 9=>x"8300", 10=>x"8000", 11=>x"8000", 12=>x"7f00", 13=>x"7f00", 14=>x"7f00",
---- 15=>x"8000", 16=>x"7f00", 17=>x"8100", 18=>x"8200", 19=>x"8000", 20=>x"8000", 21=>x"7f00",
---- 22=>x"8000", 23=>x"8000", 24=>x"7f00", 25=>x"8100", 26=>x"8200", 27=>x"7f00", 28=>x"8000",
---- 29=>x"8100", 30=>x"7e00", 31=>x"7c00", 32=>x"8000", 33=>x"8300", 34=>x"7f00", 35=>x"7f00",
---- 36=>x"8100", 37=>x"7e00", 38=>x"7d00", 39=>x"7e00", 40=>x"7d00", 41=>x"8000", 42=>x"8200",
---- 43=>x"7f00", 44=>x"8000", 45=>x"7e00", 46=>x"7f00", 47=>x"7f00", 48=>x"7f00", 49=>x"7c00",
---- 50=>x"8000", 51=>x"8100", 52=>x"7e00", 53=>x"7f00", 54=>x"8100", 55=>x"7f00", 56=>x"7f00",
---- 57=>x"7e00", 58=>x"8000", 59=>x"8300", 60=>x"7f00", 61=>x"8100", 62=>x"8200", 63=>x"7f00",
---- 64=>x"8100", 65=>x"8200", 66=>x"8000", 67=>x"8100", 68=>x"8000", 69=>x"8000", 70=>x"8100",
---- 71=>x"8200", 72=>x"8000", 73=>x"8200", 74=>x"8300", 75=>x"8100", 76=>x"8200", 77=>x"7d00",
---- 78=>x"7e00", 79=>x"8200", 80=>x"7f00", 81=>x"7e00", 82=>x"8300", 83=>x"8200", 84=>x"7e00",
---- 85=>x"7e00", 86=>x"8000", 87=>x"7f00", 88=>x"7f00", 89=>x"7c00", 90=>x"7f00", 91=>x"7f00",
---- 92=>x"7e00", 93=>x"7d00", 94=>x"8300", 95=>x"7f00", 96=>x"7e00", 97=>x"8000", 98=>x"7f00",
---- 99=>x"7d00", 100=>x"7d00", 101=>x"7b00", 102=>x"8000", 103=>x"8100", 104=>x"7f00", 105=>x"7f00",
---- 106=>x"7f00", 107=>x"7e00", 108=>x"7e00", 109=>x"8000", 110=>x"8000", 111=>x"7e00", 112=>x"7d00",
---- 113=>x"7e00", 114=>x"7e00", 115=>x"7e00", 116=>x"7c00", 117=>x"8000", 118=>x"8100", 119=>x"7d00",
---- 120=>x"7c00", 121=>x"7d00", 122=>x"7c00", 123=>x"7f00", 124=>x"7e00", 125=>x"7f00", 126=>x"8000",
---- 127=>x"8200", 128=>x"7f00", 129=>x"7d00", 130=>x"7e00", 131=>x"7e00", 132=>x"7f00", 133=>x"8000",
---- 134=>x"7f00", 135=>x"8000", 136=>x"8000", 137=>x"7f00", 138=>x"7b00", 139=>x"7d00", 140=>x"8000",
---- 141=>x"7f00", 142=>x"8000", 143=>x"7f00", 144=>x"7a00", 145=>x"7f00", 146=>x"7f00", 147=>x"7d00",
---- 148=>x"7c00", 149=>x"7d00", 150=>x"7e00", 151=>x"7e00", 152=>x"7d00", 153=>x"7c00", 154=>x"7e00",
---- 155=>x"7d00", 156=>x"8000", 157=>x"7d00", 158=>x"7d00", 159=>x"7f00", 160=>x"8000", 161=>x"7e00",
---- 162=>x"7d00", 163=>x"7f00", 164=>x"7d00", 165=>x"7c00", 166=>x"8000", 167=>x"7e00", 168=>x"7c00",
---- 169=>x"7f00", 170=>x"7d00", 171=>x"7e00", 172=>x"7e00", 173=>x"7e00", 174=>x"8000", 175=>x"7e00",
---- 176=>x"7e00", 177=>x"8000", 178=>x"8200", 179=>x"7f00", 180=>x"7f00", 181=>x"7d00", 182=>x"7e00",
---- 183=>x"8000", 184=>x"7d00", 185=>x"7e00", 186=>x"8100", 187=>x"7e00", 188=>x"7f00", 189=>x"8000",
---- 190=>x"8100", 191=>x"7f00", 192=>x"8000", 193=>x"7d00", 194=>x"7e00", 195=>x"7f00", 196=>x"7e00",
---- 197=>x"8000", 198=>x"7d00", 199=>x"7d00", 200=>x"8000", 201=>x"7e00", 202=>x"7c00", 203=>x"8100",
---- 204=>x"7f00", 205=>x"7d00", 206=>x"8000", 207=>x"7c00", 208=>x"7e00", 209=>x"8000", 210=>x"7d00",
---- 211=>x"8000", 212=>x"7c00", 213=>x"7c00", 214=>x"7d00", 215=>x"7e00", 216=>x"7e00", 217=>x"7e00",
---- 218=>x"7a00", 219=>x"7e00", 220=>x"7e00", 221=>x"7b00", 222=>x"7b00", 223=>x"7a00", 224=>x"7e00",
---- 225=>x"7b00", 226=>x"7d00", 227=>x"8000", 228=>x"7c00", 229=>x"7a00", 230=>x"7b00", 231=>x"7900",
---- 232=>x"7800", 233=>x"7900", 234=>x"7e00", 235=>x"7d00", 236=>x"7900", 237=>x"7d00", 238=>x"7b00",
---- 239=>x"7a00", 240=>x"7900", 241=>x"7900", 242=>x"7700", 243=>x"7a00", 244=>x"7600", 245=>x"7900",
---- 246=>x"7a00", 247=>x"7800", 248=>x"7700", 249=>x"7600", 250=>x"7a00", 251=>x"7900", 252=>x"7800",
---- 253=>x"7600", 254=>x"7700", 255=>x"7800", 256=>x"7400", 257=>x"7700", 258=>x"7800", 259=>x"7800",
---- 260=>x"7700", 261=>x"7800", 262=>x"7700", 263=>x"7700", 264=>x"6e00", 265=>x"7500", 266=>x"7400",
---- 267=>x"7100", 268=>x"7300", 269=>x"7300", 270=>x"7300", 271=>x"7700", 272=>x"6c00", 273=>x"6c00",
---- 274=>x"6a00", 275=>x"6c00", 276=>x"6e00", 277=>x"7100", 278=>x"7100", 279=>x"7300", 280=>x"6200",
---- 281=>x"6500", 282=>x"6800", 283=>x"6900", 284=>x"6a00", 285=>x"6c00", 286=>x"6e00", 287=>x"7200",
---- 288=>x"7500", 289=>x"5900", 290=>x"5d00", 291=>x"6000", 292=>x"6400", 293=>x"6700", 294=>x"6b00",
---- 295=>x"6c00", 296=>x"bb00", 297=>x"7b00", 298=>x"7200", 299=>x"6400", 300=>x"a700", 301=>x"6100",
---- 302=>x"6300", 303=>x"6900", 304=>x"da00", 305=>x"d500", 306=>x"cf00", 307=>x"b900", 308=>x"7600",
---- 309=>x"5500", 310=>x"5e00", 311=>x"6500", 312=>x"dc00", 313=>x"e400", 314=>x"e600", 315=>x"e900",
---- 316=>x"c400", 317=>x"6500", 318=>x"5500", 319=>x"5a00", 320=>x"d600", 321=>x"da00", 322=>x"e100",
---- 323=>x"e300", 324=>x"e600", 325=>x"9d00", 326=>x"4e00", 327=>x"5200", 328=>x"d800", 329=>x"d700",
---- 330=>x"dd00", 331=>x"e200", 332=>x"e300", 333=>x"d000", 334=>x"7700", 335=>x"4b00", 336=>x"d000",
---- 337=>x"d600", 338=>x"d800", 339=>x"df00", 340=>x"e000", 341=>x"e300", 342=>x"c400", 343=>x"6000",
---- 344=>x"cd00", 345=>x"d000", 346=>x"d800", 347=>x"da00", 348=>x"e000", 349=>x"de00", 350=>x"e200",
---- 351=>x"a500", 352=>x"d300", 353=>x"ce00", 354=>x"d000", 355=>x"d400", 356=>x"d500", 357=>x"df00",
---- 358=>x"df00", 359=>x"da00", 360=>x"cd00", 361=>x"d200", 362=>x"d200", 363=>x"d600", 364=>x"d500",
---- 365=>x"de00", 366=>x"e100", 367=>x"de00", 368=>x"d100", 369=>x"d400", 370=>x"2600", 371=>x"d900",
---- 372=>x"da00", 373=>x"df00", 374=>x"e500", 375=>x"e000", 376=>x"d700", 377=>x"d200", 378=>x"d500",
---- 379=>x"d200", 380=>x"d400", 381=>x"d800", 382=>x"dc00", 383=>x"e100", 384=>x"cb00", 385=>x"ca00",
---- 386=>x"cc00", 387=>x"ce00", 388=>x"ce00", 389=>x"d100", 390=>x"d400", 391=>x"d600", 392=>x"c700",
---- 393=>x"ce00", 394=>x"d100", 395=>x"d100", 396=>x"d400", 397=>x"d300", 398=>x"d400", 399=>x"d400",
---- 400=>x"ce00", 401=>x"cf00", 402=>x"d100", 403=>x"d300", 404=>x"d000", 405=>x"d300", 406=>x"d200",
---- 407=>x"d400", 408=>x"d000", 409=>x"d000", 410=>x"ce00", 411=>x"d200", 412=>x"d100", 413=>x"d100",
---- 414=>x"d400", 415=>x"ce00", 416=>x"cf00", 417=>x"d000", 418=>x"cd00", 419=>x"cb00", 420=>x"cf00",
---- 421=>x"d000", 422=>x"d100", 423=>x"cc00", 424=>x"ce00", 425=>x"d100", 426=>x"cf00", 427=>x"ce00",
---- 428=>x"d200", 429=>x"d100", 430=>x"d300", 431=>x"d100", 432=>x"ce00", 433=>x"d200", 434=>x"cf00",
---- 435=>x"cf00", 436=>x"cf00", 437=>x"cc00", 438=>x"ca00", 439=>x"cd00", 440=>x"cd00", 441=>x"cb00",
---- 442=>x"cc00", 443=>x"cb00", 444=>x"ca00", 445=>x"cd00", 446=>x"cb00", 447=>x"cd00", 448=>x"cb00",
---- 449=>x"c300", 450=>x"c400", 451=>x"c900", 452=>x"ca00", 453=>x"d100", 454=>x"d400", 455=>x"d100",
---- 456=>x"c800", 457=>x"cb00", 458=>x"c800", 459=>x"cb00", 460=>x"ce00", 461=>x"cf00", 462=>x"d000",
---- 463=>x"d400", 464=>x"cb00", 465=>x"d400", 466=>x"cd00", 467=>x"c400", 468=>x"ca00", 469=>x"ce00",
---- 470=>x"cf00", 471=>x"d000", 472=>x"cc00", 473=>x"ca00", 474=>x"d200", 475=>x"cd00", 476=>x"c800",
---- 477=>x"cb00", 478=>x"ce00", 479=>x"cf00", 480=>x"ce00", 481=>x"c900", 482=>x"c900", 483=>x"cd00",
---- 484=>x"cf00", 485=>x"c700", 486=>x"ca00", 487=>x"d000", 488=>x"cb00", 489=>x"c800", 490=>x"c600",
---- 491=>x"c300", 492=>x"c900", 493=>x"c700", 494=>x"c400", 495=>x"3300", 496=>x"c500", 497=>x"c600",
---- 498=>x"ca00", 499=>x"c700", 500=>x"c200", 501=>x"c900", 502=>x"c700", 503=>x"c900", 504=>x"ca00",
---- 505=>x"c600", 506=>x"c800", 507=>x"3400", 508=>x"cb00", 509=>x"c800", 510=>x"cb00", 511=>x"cb00",
---- 512=>x"cb00", 513=>x"c900", 514=>x"c600", 515=>x"c800", 516=>x"ca00", 517=>x"d000", 518=>x"cf00",
---- 519=>x"cb00", 520=>x"c600", 521=>x"cc00", 522=>x"c900", 523=>x"c300", 524=>x"c200", 525=>x"ca00",
---- 526=>x"bf00", 527=>x"ba00", 528=>x"c000", 529=>x"c900", 530=>x"cc00", 531=>x"c900", 532=>x"b100",
---- 533=>x"a200", 534=>x"b200", 535=>x"c600", 536=>x"c700", 537=>x"c600", 538=>x"cb00", 539=>x"bc00",
---- 540=>x"9e00", 541=>x"a800", 542=>x"c200", 543=>x"c600", 544=>x"ca00", 545=>x"ca00", 546=>x"af00",
---- 547=>x"9900", 548=>x"b300", 549=>x"c200", 550=>x"bd00", 551=>x"c000", 552=>x"c400", 553=>x"b100",
---- 554=>x"a800", 555=>x"b100", 556=>x"bd00", 557=>x"be00", 558=>x"c100", 559=>x"c600", 560=>x"aa00",
---- 561=>x"ab00", 562=>x"c000", 563=>x"c300", 564=>x"be00", 565=>x"bd00", 566=>x"ba00", 567=>x"bd00",
---- 568=>x"b200", 569=>x"bf00", 570=>x"bb00", 571=>x"b600", 572=>x"b200", 573=>x"b500", 574=>x"b500",
---- 575=>x"b900", 576=>x"bc00", 577=>x"bc00", 578=>x"af00", 579=>x"ab00", 580=>x"bb00", 581=>x"bc00",
---- 582=>x"c200", 583=>x"be00", 584=>x"c100", 585=>x"bd00", 586=>x"bb00", 587=>x"b600", 588=>x"bc00",
---- 589=>x"bf00", 590=>x"c200", 591=>x"c000", 592=>x"b500", 593=>x"bc00", 594=>x"bd00", 595=>x"c000",
---- 596=>x"ba00", 597=>x"bb00", 598=>x"c000", 599=>x"bd00", 600=>x"b200", 601=>x"b900", 602=>x"4600",
---- 603=>x"c100", 604=>x"bf00", 605=>x"b800", 606=>x"bb00", 607=>x"bf00", 608=>x"af00", 609=>x"b500",
---- 610=>x"b900", 611=>x"bd00", 612=>x"c000", 613=>x"bd00", 614=>x"b600", 615=>x"b500", 616=>x"b600",
---- 617=>x"ae00", 618=>x"b700", 619=>x"be00", 620=>x"bd00", 621=>x"bc00", 622=>x"b400", 623=>x"af00",
---- 624=>x"bc00", 625=>x"b700", 626=>x"b000", 627=>x"b500", 628=>x"b700", 629=>x"b200", 630=>x"b200",
---- 631=>x"b100", 632=>x"ba00", 633=>x"bb00", 634=>x"b400", 635=>x"ae00", 636=>x"af00", 637=>x"b200",
---- 638=>x"af00", 639=>x"ae00", 640=>x"af00", 641=>x"ba00", 642=>x"b400", 643=>x"af00", 644=>x"5600",
---- 645=>x"aa00", 646=>x"ae00", 647=>x"5000", 648=>x"a700", 649=>x"ac00", 650=>x"b200", 651=>x"ac00",
---- 652=>x"ab00", 653=>x"a600", 654=>x"aa00", 655=>x"af00", 656=>x"a900", 657=>x"a300", 658=>x"a100",
---- 659=>x"a400", 660=>x"ad00", 661=>x"5500", 662=>x"a300", 663=>x"a700", 664=>x"9f00", 665=>x"a400",
---- 666=>x"a000", 667=>x"a000", 668=>x"a300", 669=>x"ab00", 670=>x"9f00", 671=>x"9f00", 672=>x"a600",
---- 673=>x"9a00", 674=>x"a300", 675=>x"a900", 676=>x"9800", 677=>x"9d00", 678=>x"9f00", 679=>x"9600",
---- 680=>x"a500", 681=>x"a200", 682=>x"9e00", 683=>x"a100", 684=>x"9c00", 685=>x"9000", 686=>x"9b00",
---- 687=>x"9400", 688=>x"9800", 689=>x"a400", 690=>x"9e00", 691=>x"9100", 692=>x"9b00", 693=>x"8a00",
---- 694=>x"9700", 695=>x"b300", 696=>x"3f00", 697=>x"7f00", 698=>x"a100", 699=>x"9100", 700=>x"8800",
---- 701=>x"a100", 702=>x"bb00", 703=>x"c100", 704=>x"2d00", 705=>x"3e00", 706=>x"9a00", 707=>x"9600",
---- 708=>x"a100", 709=>x"c300", 710=>x"b400", 711=>x"9e00", 712=>x"2900", 713=>x"2600", 714=>x"7b00",
---- 715=>x"bc00", 716=>x"c100", 717=>x"a400", 718=>x"9700", 719=>x"a100", 720=>x"2400", 721=>x"5200",
---- 722=>x"a800", 723=>x"bf00", 724=>x"9900", 725=>x"9200", 726=>x"ae00", 727=>x"c000", 728=>x"7000",
---- 729=>x"b200", 730=>x"b400", 731=>x"8b00", 732=>x"9600", 733=>x"b900", 734=>x"cb00", 735=>x"cc00",
---- 736=>x"be00", 737=>x"a100", 738=>x"8900", 739=>x"9800", 740=>x"b300", 741=>x"c600", 742=>x"c900",
---- 743=>x"cb00", 744=>x"9200", 745=>x"7300", 746=>x"9e00", 747=>x"c400", 748=>x"be00", 749=>x"bc00",
---- 750=>x"be00", 751=>x"3f00", 752=>x"6b00", 753=>x"9800", 754=>x"c300", 755=>x"c700", 756=>x"bf00",
---- 757=>x"b800", 758=>x"b800", 759=>x"b800", 760=>x"a100", 761=>x"bb00", 762=>x"c200", 763=>x"be00",
---- 764=>x"b500", 765=>x"b200", 766=>x"b400", 767=>x"b900", 768=>x"c700", 769=>x"be00", 770=>x"bf00",
---- 771=>x"b700", 772=>x"b300", 773=>x"b500", 774=>x"ba00", 775=>x"bc00", 776=>x"c300", 777=>x"bc00",
---- 778=>x"ba00", 779=>x"b700", 780=>x"b400", 781=>x"b400", 782=>x"b800", 783=>x"bb00", 784=>x"be00",
---- 785=>x"b600", 786=>x"b700", 787=>x"b200", 788=>x"b300", 789=>x"b700", 790=>x"ba00", 791=>x"b700",
---- 792=>x"bb00", 793=>x"b400", 794=>x"b000", 795=>x"b300", 796=>x"b700", 797=>x"b600", 798=>x"b800",
---- 799=>x"b600", 800=>x"bc00", 801=>x"b500", 802=>x"b300", 803=>x"b300", 804=>x"b700", 805=>x"b400",
---- 806=>x"b300", 807=>x"b600", 808=>x"bd00", 809=>x"b900", 810=>x"b600", 811=>x"b700", 812=>x"b500",
---- 813=>x"b300", 814=>x"b700", 815=>x"b300", 816=>x"ba00", 817=>x"b500", 818=>x"4a00", 819=>x"b100",
---- 820=>x"b400", 821=>x"b800", 822=>x"b800", 823=>x"b300", 824=>x"b600", 825=>x"b300", 826=>x"b200",
---- 827=>x"b200", 828=>x"b400", 829=>x"b500", 830=>x"b400", 831=>x"ad00", 832=>x"b400", 833=>x"b200",
---- 834=>x"b400", 835=>x"b100", 836=>x"b400", 837=>x"b200", 838=>x"ad00", 839=>x"ac00", 840=>x"ad00",
---- 841=>x"af00", 842=>x"b200", 843=>x"af00", 844=>x"ae00", 845=>x"ae00", 846=>x"af00", 847=>x"b000",
---- 848=>x"a500", 849=>x"ad00", 850=>x"b000", 851=>x"ab00", 852=>x"ae00", 853=>x"af00", 854=>x"b200",
---- 855=>x"ad00", 856=>x"a900", 857=>x"b100", 858=>x"ae00", 859=>x"b000", 860=>x"b100", 861=>x"b000",
---- 862=>x"ab00", 863=>x"af00", 864=>x"aa00", 865=>x"ac00", 866=>x"b200", 867=>x"b300", 868=>x"b000",
---- 869=>x"a600", 870=>x"9f00", 871=>x"ac00", 872=>x"a600", 873=>x"a900", 874=>x"b300", 875=>x"b500",
---- 876=>x"ab00", 877=>x"9d00", 878=>x"9f00", 879=>x"a800", 880=>x"a900", 881=>x"b000", 882=>x"b700",
---- 883=>x"b300", 884=>x"a400", 885=>x"a000", 886=>x"a900", 887=>x"ae00", 888=>x"ad00", 889=>x"b900",
---- 890=>x"b400", 891=>x"a100", 892=>x"9c00", 893=>x"a600", 894=>x"ab00", 895=>x"b100", 896=>x"b500",
---- 897=>x"ae00", 898=>x"9500", 899=>x"9e00", 900=>x"5a00", 901=>x"ac00", 902=>x"b100", 903=>x"b700",
---- 904=>x"a600", 905=>x"9400", 906=>x"9a00", 907=>x"a400", 908=>x"a900", 909=>x"ad00", 910=>x"b000",
---- 911=>x"bb00", 912=>x"9400", 913=>x"9700", 914=>x"a400", 915=>x"a800", 916=>x"a900", 917=>x"5100",
---- 918=>x"b500", 919=>x"be00", 920=>x"9e00", 921=>x"9f00", 922=>x"a400", 923=>x"ab00", 924=>x"a900",
---- 925=>x"ae00", 926=>x"b800", 927=>x"bb00", 928=>x"9f00", 929=>x"a600", 930=>x"a800", 931=>x"ac00",
---- 932=>x"a900", 933=>x"b100", 934=>x"b700", 935=>x"4400", 936=>x"a500", 937=>x"ab00", 938=>x"ac00",
---- 939=>x"ad00", 940=>x"af00", 941=>x"af00", 942=>x"b500", 943=>x"b900", 944=>x"a800", 945=>x"ad00",
---- 946=>x"ab00", 947=>x"ae00", 948=>x"b100", 949=>x"b200", 950=>x"b400", 951=>x"b800", 952=>x"aa00",
---- 953=>x"ae00", 954=>x"ac00", 955=>x"ae00", 956=>x"af00", 957=>x"b400", 958=>x"b400", 959=>x"b600",
---- 960=>x"ab00", 961=>x"b000", 962=>x"b000", 963=>x"af00", 964=>x"b000", 965=>x"b200", 966=>x"b000",
---- 967=>x"b200", 968=>x"af00", 969=>x"af00", 970=>x"b200", 971=>x"b200", 972=>x"b200", 973=>x"b100",
---- 974=>x"b200", 975=>x"b700", 976=>x"af00", 977=>x"b100", 978=>x"b300", 979=>x"b500", 980=>x"b100",
---- 981=>x"af00", 982=>x"b000", 983=>x"b100", 984=>x"ab00", 985=>x"b200", 986=>x"b600", 987=>x"b500",
---- 988=>x"b100", 989=>x"b100", 990=>x"b200", 991=>x"af00", 992=>x"8d00", 993=>x"a600", 994=>x"b100",
---- 995=>x"b200", 996=>x"af00", 997=>x"b400", 998=>x"b200", 999=>x"ad00", 1000=>x"4e00", 1001=>x"6a00",
---- 1002=>x"8f00", 1003=>x"5700", 1004=>x"ac00", 1005=>x"ad00", 1006=>x"ab00", 1007=>x"ab00", 1008=>x"4800",
---- 1009=>x"4800", 1010=>x"6300", 1011=>x"8700", 1012=>x"a300", 1013=>x"a700", 1014=>x"a700", 1015=>x"a900",
---- 1016=>x"6600", 1017=>x"6100", 1018=>x"6500", 1019=>x"7700", 1020=>x"9400", 1021=>x"9d00", 1022=>x"9e00",
---- 1023=>x"a400", 1024=>x"7800", 1025=>x"7500", 1026=>x"7300", 1027=>x"7900", 1028=>x"8600", 1029=>x"9400",
---- 1030=>x"9b00", 1031=>x"a100", 1032=>x"8100", 1033=>x"7d00", 1034=>x"7e00", 1035=>x"7e00", 1036=>x"8900",
---- 1037=>x"8c00", 1038=>x"9400", 1039=>x"9d00", 1040=>x"8800", 1041=>x"8400", 1042=>x"8000", 1043=>x"7f00",
---- 1044=>x"8800", 1045=>x"8d00", 1046=>x"6e00", 1047=>x"9600", 1048=>x"7700", 1049=>x"7700", 1050=>x"8000",
---- 1051=>x"7e00", 1052=>x"8500", 1053=>x"8900", 1054=>x"9100", 1055=>x"9500", 1056=>x"6600", 1057=>x"8200",
---- 1058=>x"7800", 1059=>x"7c00", 1060=>x"8600", 1061=>x"8800", 1062=>x"8f00", 1063=>x"9200", 1064=>x"5c00",
---- 1065=>x"7b00", 1066=>x"7200", 1067=>x"7800", 1068=>x"8300", 1069=>x"8600", 1070=>x"8b00", 1071=>x"8e00",
---- 1072=>x"6000", 1073=>x"6c00", 1074=>x"6f00", 1075=>x"7300", 1076=>x"7a00", 1077=>x"8200", 1078=>x"8700",
---- 1079=>x"8d00", 1080=>x"7300", 1081=>x"6a00", 1082=>x"7800", 1083=>x"7500", 1084=>x"7800", 1085=>x"8100",
---- 1086=>x"8800", 1087=>x"8e00", 1088=>x"8000", 1089=>x"7600", 1090=>x"7600", 1091=>x"7900", 1092=>x"7d00",
---- 1093=>x"8100", 1094=>x"8500", 1095=>x"8900", 1096=>x"8400", 1097=>x"8000", 1098=>x"7700", 1099=>x"8800",
---- 1100=>x"7f00", 1101=>x"8000", 1102=>x"8000", 1103=>x"8c00", 1104=>x"8200", 1105=>x"7d00", 1106=>x"7a00",
---- 1107=>x"7a00", 1108=>x"7d00", 1109=>x"8000", 1110=>x"8000", 1111=>x"8b00", 1112=>x"7c00", 1113=>x"7700",
---- 1114=>x"7f00", 1115=>x"8400", 1116=>x"8000", 1117=>x"8100", 1118=>x"7f00", 1119=>x"8900", 1120=>x"8000",
---- 1121=>x"7800", 1122=>x"8400", 1123=>x"8500", 1124=>x"8200", 1125=>x"8100", 1126=>x"7d00", 1127=>x"8400",
---- 1128=>x"8300", 1129=>x"8100", 1130=>x"8600", 1131=>x"8800", 1132=>x"8400", 1133=>x"8000", 1134=>x"7f00",
---- 1135=>x"8000", 1136=>x"8200", 1137=>x"8400", 1138=>x"8a00", 1139=>x"8900", 1140=>x"8100", 1141=>x"7f00",
---- 1142=>x"8100", 1143=>x"8000", 1144=>x"8800", 1145=>x"8d00", 1146=>x"8f00", 1147=>x"8800", 1148=>x"8400",
---- 1149=>x"8100", 1150=>x"8300", 1151=>x"7f00", 1152=>x"8900", 1153=>x"8f00", 1154=>x"8b00", 1155=>x"8500",
---- 1156=>x"8300", 1157=>x"8200", 1158=>x"8100", 1159=>x"8000", 1160=>x"8b00", 1161=>x"8f00", 1162=>x"9000",
---- 1163=>x"8800", 1164=>x"8100", 1165=>x"8200", 1166=>x"7f00", 1167=>x"7c00", 1168=>x"9400", 1169=>x"9200",
---- 1170=>x"8f00", 1171=>x"8a00", 1172=>x"8300", 1173=>x"8600", 1174=>x"8100", 1175=>x"8100", 1176=>x"9200",
---- 1177=>x"9200", 1178=>x"8f00", 1179=>x"8a00", 1180=>x"8300", 1181=>x"8500", 1182=>x"8300", 1183=>x"8000",
---- 1184=>x"9400", 1185=>x"9200", 1186=>x"9200", 1187=>x"8c00", 1188=>x"8700", 1189=>x"8400", 1190=>x"8000",
---- 1191=>x"8100", 1192=>x"9300", 1193=>x"9300", 1194=>x"9000", 1195=>x"8b00", 1196=>x"8700", 1197=>x"8100",
---- 1198=>x"7e00", 1199=>x"8500", 1200=>x"8d00", 1201=>x"9000", 1202=>x"8f00", 1203=>x"8900", 1204=>x"8500",
---- 1205=>x"7d00", 1206=>x"7e00", 1207=>x"8200", 1208=>x"8900", 1209=>x"8b00", 1210=>x"8c00", 1211=>x"8800",
---- 1212=>x"8100", 1213=>x"7d00", 1214=>x"7d00", 1215=>x"8000", 1216=>x"8700", 1217=>x"8600", 1218=>x"7600",
---- 1219=>x"8700", 1220=>x"7d00", 1221=>x"7f00", 1222=>x"7c00", 1223=>x"7e00", 1224=>x"7a00", 1225=>x"8500",
---- 1226=>x"8600", 1227=>x"8300", 1228=>x"8000", 1229=>x"7c00", 1230=>x"7900", 1231=>x"7c00", 1232=>x"8400",
---- 1233=>x"8400", 1234=>x"8500", 1235=>x"8100", 1236=>x"8000", 1237=>x"7b00", 1238=>x"7800", 1239=>x"7c00",
---- 1240=>x"8400", 1241=>x"8200", 1242=>x"8400", 1243=>x"7f00", 1244=>x"7c00", 1245=>x"7b00", 1246=>x"7800",
---- 1247=>x"7a00", 1248=>x"7f00", 1249=>x"7d00", 1250=>x"8000", 1251=>x"8500", 1252=>x"7e00", 1253=>x"7b00",
---- 1254=>x"7b00", 1255=>x"7600", 1256=>x"7500", 1257=>x"7c00", 1258=>x"8400", 1259=>x"8900", 1260=>x"8200",
---- 1261=>x"7d00", 1262=>x"7c00", 1263=>x"7900", 1264=>x"7100", 1265=>x"8000", 1266=>x"8700", 1267=>x"8800",
---- 1268=>x"8900", 1269=>x"8900", 1270=>x"8300", 1271=>x"7c00", 1272=>x"7500", 1273=>x"8500", 1274=>x"8c00",
---- 1275=>x"8b00", 1276=>x"8c00", 1277=>x"8e00", 1278=>x"8d00", 1279=>x"8200", 1280=>x"7900", 1281=>x"8600",
---- 1282=>x"8900", 1283=>x"8800", 1284=>x"8500", 1285=>x"8b00", 1286=>x"8900", 1287=>x"8700", 1288=>x"8000",
---- 1289=>x"8500", 1290=>x"8400", 1291=>x"5b00", 1292=>x"3e00", 1293=>x"4f00", 1294=>x"6900", 1295=>x"7200",
---- 1296=>x"7a00", 1297=>x"8500", 1298=>x"7c00", 1299=>x"5400", 1300=>x"3c00", 1301=>x"5000", 1302=>x"6000",
---- 1303=>x"a700", 1304=>x"7700", 1305=>x"7c00", 1306=>x"7d00", 1307=>x"7e00", 1308=>x"7c00", 1309=>x"8000",
---- 1310=>x"8100", 1311=>x"7600", 1312=>x"8600", 1313=>x"8200", 1314=>x"7c00", 1315=>x"7f00", 1316=>x"8300",
---- 1317=>x"8400", 1318=>x"8600", 1319=>x"7d00", 1320=>x"9100", 1321=>x"8f00", 1322=>x"7a00", 1323=>x"8300",
---- 1324=>x"8100", 1325=>x"8600", 1326=>x"9100", 1327=>x"8e00", 1328=>x"9300", 1329=>x"9200", 1330=>x"8f00",
---- 1331=>x"8a00", 1332=>x"8b00", 1333=>x"9300", 1334=>x"a700", 1335=>x"b300", 1336=>x"9400", 1337=>x"9400",
---- 1338=>x"9000", 1339=>x"8f00", 1340=>x"9500", 1341=>x"a000", 1342=>x"b900", 1343=>x"c500", 1344=>x"9300",
---- 1345=>x"9300", 1346=>x"9200", 1347=>x"9400", 1348=>x"9900", 1349=>x"a700", 1350=>x"c400", 1351=>x"cc00",
---- 1352=>x"9700", 1353=>x"9400", 1354=>x"9700", 1355=>x"9900", 1356=>x"9f00", 1357=>x"ae00", 1358=>x"cc00",
---- 1359=>x"ce00", 1360=>x"9500", 1361=>x"9900", 1362=>x"9a00", 1363=>x"9b00", 1364=>x"a200", 1365=>x"b200",
---- 1366=>x"d100", 1367=>x"cf00", 1368=>x"9400", 1369=>x"9500", 1370=>x"9900", 1371=>x"9c00", 1372=>x"a200",
---- 1373=>x"b500", 1374=>x"cd00", 1375=>x"d400", 1376=>x"9400", 1377=>x"9a00", 1378=>x"9d00", 1379=>x"a000",
---- 1380=>x"a400", 1381=>x"a900", 1382=>x"b400", 1383=>x"bb00", 1384=>x"9400", 1385=>x"9200", 1386=>x"9300",
---- 1387=>x"8d00", 1388=>x"8b00", 1389=>x"8600", 1390=>x"8e00", 1391=>x"9000", 1392=>x"7b00", 1393=>x"7a00",
---- 1394=>x"7d00", 1395=>x"7900", 1396=>x"7800", 1397=>x"7400", 1398=>x"7c00", 1399=>x"8500", 1400=>x"6300",
---- 1401=>x"6100", 1402=>x"5d00", 1403=>x"5800", 1404=>x"5e00", 1405=>x"6400", 1406=>x"8f00", 1407=>x"7600",
---- 1408=>x"7000", 1409=>x"6e00", 1410=>x"6a00", 1411=>x"6600", 1412=>x"6a00", 1413=>x"6c00", 1414=>x"7500",
---- 1415=>x"7d00", 1416=>x"8400", 1417=>x"8c00", 1418=>x"9400", 1419=>x"9300", 1420=>x"9700", 1421=>x"9900",
---- 1422=>x"9f00", 1423=>x"ae00", 1424=>x"8900", 1425=>x"9900", 1426=>x"a900", 1427=>x"b400", 1428=>x"b800",
---- 1429=>x"b900", 1430=>x"b800", 1431=>x"c800", 1432=>x"8500", 1433=>x"9500", 1434=>x"9600", 1435=>x"9d00",
---- 1436=>x"a500", 1437=>x"a300", 1438=>x"9a00", 1439=>x"9e00", 1440=>x"8000", 1441=>x"8900", 1442=>x"8e00",
---- 1443=>x"9000", 1444=>x"9200", 1445=>x"9600", 1446=>x"9100", 1447=>x"8b00", 1448=>x"7b00", 1449=>x"8100",
---- 1450=>x"8700", 1451=>x"7900", 1452=>x"8e00", 1453=>x"8d00", 1454=>x"8900", 1455=>x"8700", 1456=>x"7600",
---- 1457=>x"7600", 1458=>x"7700", 1459=>x"7800", 1460=>x"7d00", 1461=>x"7800", 1462=>x"7600", 1463=>x"7700",
---- 1464=>x"7e00", 1465=>x"7b00", 1466=>x"7600", 1467=>x"7700", 1468=>x"7900", 1469=>x"7d00", 1470=>x"8100",
---- 1471=>x"7300", 1472=>x"8f00", 1473=>x"9000", 1474=>x"9000", 1475=>x"9200", 1476=>x"9000", 1477=>x"6a00",
---- 1478=>x"9a00", 1479=>x"9b00", 1480=>x"9900", 1481=>x"9f00", 1482=>x"a400", 1483=>x"a300", 1484=>x"9e00",
---- 1485=>x"9b00", 1486=>x"9c00", 1487=>x"9e00", 1488=>x"a400", 1489=>x"a600", 1490=>x"a900", 1491=>x"ac00",
---- 1492=>x"a400", 1493=>x"9e00", 1494=>x"9c00", 1495=>x"9d00", 1496=>x"a600", 1497=>x"a900", 1498=>x"ab00",
---- 1499=>x"a900", 1500=>x"a900", 1501=>x"a300", 1502=>x"a300", 1503=>x"a200", 1504=>x"a400", 1505=>x"aa00",
---- 1506=>x"a600", 1507=>x"a200", 1508=>x"a900", 1509=>x"a800", 1510=>x"a700", 1511=>x"a400", 1512=>x"a700",
---- 1513=>x"a800", 1514=>x"a600", 1515=>x"a500", 1516=>x"a900", 1517=>x"ad00", 1518=>x"af00", 1519=>x"a400",
---- 1520=>x"aa00", 1521=>x"ab00", 1522=>x"a800", 1523=>x"a600", 1524=>x"a900", 1525=>x"aa00", 1526=>x"a800",
---- 1527=>x"9f00", 1528=>x"a800", 1529=>x"ac00", 1530=>x"a800", 1531=>x"a200", 1532=>x"a300", 1533=>x"a300",
---- 1534=>x"9e00", 1535=>x"9b00", 1536=>x"a400", 1537=>x"a400", 1538=>x"5d00", 1539=>x"9a00", 1540=>x"9a00",
---- 1541=>x"9a00", 1542=>x"9b00", 1543=>x"9400", 1544=>x"a200", 1545=>x"a400", 1546=>x"5f00", 1547=>x"9800",
---- 1548=>x"9800", 1549=>x"9900", 1550=>x"9200", 1551=>x"8500", 1552=>x"a200", 1553=>x"a700", 1554=>x"a600",
---- 1555=>x"a800", 1556=>x"ad00", 1557=>x"aa00", 1558=>x"a200", 1559=>x"9d00", 1560=>x"9a00", 1561=>x"9d00",
---- 1562=>x"9e00", 1563=>x"a000", 1564=>x"a100", 1565=>x"a000", 1566=>x"a900", 1567=>x"b200", 1568=>x"9700",
---- 1569=>x"9500", 1570=>x"9400", 1571=>x"9600", 1572=>x"9900", 1573=>x"9c00", 1574=>x"a600", 1575=>x"ad00",
---- 1576=>x"8f00", 1577=>x"9000", 1578=>x"9100", 1579=>x"9200", 1580=>x"6700", 1581=>x"a100", 1582=>x"aa00",
---- 1583=>x"ae00", 1584=>x"8e00", 1585=>x"9000", 1586=>x"8f00", 1587=>x"9500", 1588=>x"9800", 1589=>x"a400",
---- 1590=>x"ac00", 1591=>x"b000", 1592=>x"8e00", 1593=>x"8f00", 1594=>x"9000", 1595=>x"9500", 1596=>x"9a00",
---- 1597=>x"a600", 1598=>x"ab00", 1599=>x"b300", 1600=>x"8f00", 1601=>x"9000", 1602=>x"9400", 1603=>x"9800",
---- 1604=>x"9f00", 1605=>x"a700", 1606=>x"ae00", 1607=>x"b700", 1608=>x"8e00", 1609=>x"9500", 1610=>x"9700",
---- 1611=>x"9d00", 1612=>x"a200", 1613=>x"a900", 1614=>x"ae00", 1615=>x"b500", 1616=>x"9100", 1617=>x"9300",
---- 1618=>x"9900", 1619=>x"9d00", 1620=>x"a600", 1621=>x"ad00", 1622=>x"b100", 1623=>x"b500", 1624=>x"9200",
---- 1625=>x"9700", 1626=>x"9c00", 1627=>x"a200", 1628=>x"a400", 1629=>x"a900", 1630=>x"ac00", 1631=>x"b300",
---- 1632=>x"9500", 1633=>x"9b00", 1634=>x"9e00", 1635=>x"a100", 1636=>x"a400", 1637=>x"a700", 1638=>x"a800",
---- 1639=>x"b000", 1640=>x"9800", 1641=>x"9b00", 1642=>x"9f00", 1643=>x"a100", 1644=>x"a300", 1645=>x"a600",
---- 1646=>x"a900", 1647=>x"4f00", 1648=>x"9800", 1649=>x"9c00", 1650=>x"a200", 1651=>x"a200", 1652=>x"a400",
---- 1653=>x"a800", 1654=>x"a700", 1655=>x"aa00", 1656=>x"9900", 1657=>x"9d00", 1658=>x"a100", 1659=>x"a000",
---- 1660=>x"a200", 1661=>x"a500", 1662=>x"a500", 1663=>x"a900", 1664=>x"6800", 1665=>x"9900", 1666=>x"a000",
---- 1667=>x"a100", 1668=>x"a100", 1669=>x"a200", 1670=>x"a500", 1671=>x"a800", 1672=>x"9700", 1673=>x"9800",
---- 1674=>x"9c00", 1675=>x"a000", 1676=>x"a100", 1677=>x"a100", 1678=>x"a400", 1679=>x"a500", 1680=>x"9700",
---- 1681=>x"9800", 1682=>x"9b00", 1683=>x"9e00", 1684=>x"9f00", 1685=>x"a200", 1686=>x"a200", 1687=>x"a500",
---- 1688=>x"9500", 1689=>x"9800", 1690=>x"9a00", 1691=>x"9d00", 1692=>x"a100", 1693=>x"a000", 1694=>x"a300",
---- 1695=>x"a500", 1696=>x"9400", 1697=>x"9600", 1698=>x"9900", 1699=>x"9b00", 1700=>x"9e00", 1701=>x"9f00",
---- 1702=>x"a200", 1703=>x"a400", 1704=>x"9500", 1705=>x"9600", 1706=>x"9700", 1707=>x"9a00", 1708=>x"9b00",
---- 1709=>x"9e00", 1710=>x"9f00", 1711=>x"a200", 1712=>x"9300", 1713=>x"9600", 1714=>x"9900", 1715=>x"9e00",
---- 1716=>x"9c00", 1717=>x"9d00", 1718=>x"a000", 1719=>x"9f00", 1720=>x"9000", 1721=>x"9500", 1722=>x"9900",
---- 1723=>x"6600", 1724=>x"9a00", 1725=>x"9c00", 1726=>x"9b00", 1727=>x"a000", 1728=>x"9200", 1729=>x"9300",
---- 1730=>x"9700", 1731=>x"9900", 1732=>x"9a00", 1733=>x"9b00", 1734=>x"9e00", 1735=>x"a000", 1736=>x"9200",
---- 1737=>x"9200", 1738=>x"9500", 1739=>x"9700", 1740=>x"9900", 1741=>x"9a00", 1742=>x"9d00", 1743=>x"a100",
---- 1744=>x"9300", 1745=>x"9400", 1746=>x"9500", 1747=>x"9600", 1748=>x"9c00", 1749=>x"9c00", 1750=>x"9f00",
---- 1751=>x"9f00", 1752=>x"9100", 1753=>x"9300", 1754=>x"9500", 1755=>x"9400", 1756=>x"9b00", 1757=>x"9b00",
---- 1758=>x"9d00", 1759=>x"9e00", 1760=>x"8f00", 1761=>x"9200", 1762=>x"9300", 1763=>x"9200", 1764=>x"9700",
---- 1765=>x"9a00", 1766=>x"9b00", 1767=>x"9d00", 1768=>x"8d00", 1769=>x"9000", 1770=>x"9300", 1771=>x"9400",
---- 1772=>x"9500", 1773=>x"9900", 1774=>x"9b00", 1775=>x"9e00", 1776=>x"8c00", 1777=>x"8e00", 1778=>x"9400",
---- 1779=>x"9700", 1780=>x"9600", 1781=>x"9a00", 1782=>x"9c00", 1783=>x"9b00", 1784=>x"8f00", 1785=>x"8e00",
---- 1786=>x"9300", 1787=>x"9300", 1788=>x"9600", 1789=>x"9800", 1790=>x"9700", 1791=>x"9a00", 1792=>x"8e00",
---- 1793=>x"8e00", 1794=>x"9100", 1795=>x"9200", 1796=>x"9400", 1797=>x"9400", 1798=>x"9600", 1799=>x"9d00",
---- 1800=>x"8e00", 1801=>x"8e00", 1802=>x"9100", 1803=>x"9000", 1804=>x"9300", 1805=>x"9500", 1806=>x"9800",
---- 1807=>x"9b00", 1808=>x"8b00", 1809=>x"8e00", 1810=>x"9200", 1811=>x"9200", 1812=>x"9400", 1813=>x"6b00",
---- 1814=>x"9600", 1815=>x"9a00", 1816=>x"8e00", 1817=>x"8e00", 1818=>x"8f00", 1819=>x"9200", 1820=>x"9400",
---- 1821=>x"9600", 1822=>x"9700", 1823=>x"9800", 1824=>x"9000", 1825=>x"8d00", 1826=>x"8f00", 1827=>x"9200",
---- 1828=>x"9200", 1829=>x"9400", 1830=>x"9300", 1831=>x"9800", 1832=>x"8e00", 1833=>x"8d00", 1834=>x"8f00",
---- 1835=>x"9000", 1836=>x"9400", 1837=>x"9400", 1838=>x"9400", 1839=>x"9700", 1840=>x"8c00", 1841=>x"8f00",
---- 1842=>x"8e00", 1843=>x"9000", 1844=>x"9400", 1845=>x"9500", 1846=>x"9400", 1847=>x"9700", 1848=>x"8b00",
---- 1849=>x"8d00", 1850=>x"9100", 1851=>x"9100", 1852=>x"9400", 1853=>x"9500", 1854=>x"9600", 1855=>x"9700",
---- 1856=>x"8c00", 1857=>x"8a00", 1858=>x"8e00", 1859=>x"9100", 1860=>x"9000", 1861=>x"9100", 1862=>x"9500",
---- 1863=>x"6900", 1864=>x"7500", 1865=>x"8a00", 1866=>x"8e00", 1867=>x"8e00", 1868=>x"8f00", 1869=>x"9200",
---- 1870=>x"9100", 1871=>x"9500", 1872=>x"8600", 1873=>x"8900", 1874=>x"8e00", 1875=>x"8c00", 1876=>x"8f00",
---- 1877=>x"8e00", 1878=>x"9000", 1879=>x"9300", 1880=>x"8800", 1881=>x"7400", 1882=>x"8c00", 1883=>x"8b00",
---- 1884=>x"8f00", 1885=>x"9200", 1886=>x"8f00", 1887=>x"9200", 1888=>x"8a00", 1889=>x"8a00", 1890=>x"8a00",
---- 1891=>x"8700", 1892=>x"8c00", 1893=>x"8f00", 1894=>x"8f00", 1895=>x"9100", 1896=>x"8600", 1897=>x"8d00",
---- 1898=>x"8900", 1899=>x"8900", 1900=>x"8b00", 1901=>x"8d00", 1902=>x"7200", 1903=>x"8f00", 1904=>x"8900",
---- 1905=>x"8c00", 1906=>x"8a00", 1907=>x"8b00", 1908=>x"8c00", 1909=>x"8b00", 1910=>x"8b00", 1911=>x"8e00",
---- 1912=>x"8800", 1913=>x"8800", 1914=>x"8900", 1915=>x"8c00", 1916=>x"8c00", 1917=>x"8800", 1918=>x"8b00",
---- 1919=>x"8e00", 1920=>x"8700", 1921=>x"8900", 1922=>x"8b00", 1923=>x"8b00", 1924=>x"8c00", 1925=>x"8a00",
---- 1926=>x"8b00", 1927=>x"8c00", 1928=>x"7800", 1929=>x"8b00", 1930=>x"8b00", 1931=>x"7200", 1932=>x"8c00",
---- 1933=>x"8e00", 1934=>x"7300", 1935=>x"8c00", 1936=>x"8a00", 1937=>x"8d00", 1938=>x"8a00", 1939=>x"8e00",
---- 1940=>x"8900", 1941=>x"8a00", 1942=>x"8900", 1943=>x"8a00", 1944=>x"8b00", 1945=>x"8e00", 1946=>x"8b00",
---- 1947=>x"8e00", 1948=>x"8b00", 1949=>x"8a00", 1950=>x"8b00", 1951=>x"8a00", 1952=>x"8e00", 1953=>x"8d00",
---- 1954=>x"8b00", 1955=>x"8c00", 1956=>x"8b00", 1957=>x"8b00", 1958=>x"8c00", 1959=>x"8b00", 1960=>x"8f00",
---- 1961=>x"9000", 1962=>x"8b00", 1963=>x"8900", 1964=>x"8c00", 1965=>x"8f00", 1966=>x"8d00", 1967=>x"8d00",
---- 1968=>x"8e00", 1969=>x"8e00", 1970=>x"8c00", 1971=>x"8900", 1972=>x"8900", 1973=>x"8c00", 1974=>x"8f00",
---- 1975=>x"8e00", 1976=>x"9000", 1977=>x"8d00", 1978=>x"9000", 1979=>x"8e00", 1980=>x"8b00", 1981=>x"8e00",
---- 1982=>x"8f00", 1983=>x"8e00", 1984=>x"9000", 1985=>x"8f00", 1986=>x"9200", 1987=>x"8e00", 1988=>x"8d00",
---- 1989=>x"8f00", 1990=>x"8b00", 1991=>x"8d00", 1992=>x"9100", 1993=>x"8f00", 1994=>x"9500", 1995=>x"9300",
---- 1996=>x"8e00", 1997=>x"8f00", 1998=>x"8f00", 1999=>x"9200", 2000=>x"9100", 2001=>x"6f00", 2002=>x"9400",
---- 2003=>x"9200", 2004=>x"9100", 2005=>x"9000", 2006=>x"8f00", 2007=>x"9100", 2008=>x"9100", 2009=>x"9200",
---- 2010=>x"9700", 2011=>x"9100", 2012=>x"6a00", 2013=>x"9400", 2014=>x"9000", 2015=>x"9400", 2016=>x"9300",
---- 2017=>x"9200", 2018=>x"9200", 2019=>x"9300", 2020=>x"9500", 2021=>x"9100", 2022=>x"9100", 2023=>x"9700",
---- 2024=>x"9400", 2025=>x"9100", 2026=>x"9100", 2027=>x"9100", 2028=>x"9700", 2029=>x"9500", 2030=>x"6a00",
---- 2031=>x"9600", 2032=>x"9200", 2033=>x"9200", 2034=>x"9300", 2035=>x"9200", 2036=>x"9500", 2037=>x"9500",
---- 2038=>x"9400", 2039=>x"9100", 2040=>x"9300", 2041=>x"9000", 2042=>x"9200", 2043=>x"9000", 2044=>x"9400",
---- 2045=>x"9400", 2046=>x"9700", 2047=>x"9600"),
---- 19 => (0=>x"7d00", 1=>x"7c00", 2=>x"7800", 3=>x"7a00", 4=>x"7500", 5=>x"7100", 6=>x"7000", 7=>x"6600",
---- 8=>x"8300", 9=>x"7b00", 10=>x"7800", 11=>x"7900", 12=>x"7600", 13=>x"7100", 14=>x"7000",
---- 15=>x"6600", 16=>x"7a00", 17=>x"7a00", 18=>x"7a00", 19=>x"7800", 20=>x"7300", 21=>x"7200",
---- 22=>x"6f00", 23=>x"6600", 24=>x"7c00", 25=>x"7900", 26=>x"7b00", 27=>x"7800", 28=>x"7300",
---- 29=>x"7100", 30=>x"6c00", 31=>x"6700", 32=>x"7c00", 33=>x"7c00", 34=>x"7800", 35=>x"7700",
---- 36=>x"7400", 37=>x"7000", 38=>x"6f00", 39=>x"6d00", 40=>x"7c00", 41=>x"7b00", 42=>x"7600",
---- 43=>x"7700", 44=>x"7500", 45=>x"7200", 46=>x"6f00", 47=>x"6b00", 48=>x"7c00", 49=>x"7b00",
---- 50=>x"7a00", 51=>x"7a00", 52=>x"7500", 53=>x"7100", 54=>x"6f00", 55=>x"6e00", 56=>x"7b00",
---- 57=>x"8300", 58=>x"7c00", 59=>x"7900", 60=>x"7600", 61=>x"7200", 62=>x"6e00", 63=>x"7300",
---- 64=>x"8000", 65=>x"7c00", 66=>x"7900", 67=>x"7900", 68=>x"7600", 69=>x"7500", 70=>x"7200",
---- 71=>x"7700", 72=>x"7e00", 73=>x"7d00", 74=>x"7d00", 75=>x"7a00", 76=>x"7400", 77=>x"7200",
---- 78=>x"7100", 79=>x"7200", 80=>x"7e00", 81=>x"7c00", 82=>x"7b00", 83=>x"7b00", 84=>x"8000",
---- 85=>x"7900", 86=>x"7100", 87=>x"7100", 88=>x"7e00", 89=>x"7b00", 90=>x"7b00", 91=>x"7a00",
---- 92=>x"7900", 93=>x"7800", 94=>x"7200", 95=>x"7100", 96=>x"7d00", 97=>x"7c00", 98=>x"7e00",
---- 99=>x"7900", 100=>x"7900", 101=>x"7800", 102=>x"7300", 103=>x"6e00", 104=>x"7e00", 105=>x"7c00",
---- 106=>x"7a00", 107=>x"7a00", 108=>x"7e00", 109=>x"7d00", 110=>x"7400", 111=>x"6e00", 112=>x"7d00",
---- 113=>x"7b00", 114=>x"7b00", 115=>x"7900", 116=>x"7900", 117=>x"7900", 118=>x"7700", 119=>x"7100",
---- 120=>x"8000", 121=>x"8100", 122=>x"7d00", 123=>x"7700", 124=>x"7400", 125=>x"7700", 126=>x"7600",
---- 127=>x"7400", 128=>x"7c00", 129=>x"8000", 130=>x"7c00", 131=>x"7900", 132=>x"7700", 133=>x"7800",
---- 134=>x"7300", 135=>x"7000", 136=>x"7d00", 137=>x"7e00", 138=>x"7d00", 139=>x"7a00", 140=>x"7a00",
---- 141=>x"7700", 142=>x"7400", 143=>x"6f00", 144=>x"8000", 145=>x"7c00", 146=>x"7b00", 147=>x"7900",
---- 148=>x"7800", 149=>x"7500", 150=>x"7700", 151=>x"7400", 152=>x"8100", 153=>x"7d00", 154=>x"7c00",
---- 155=>x"7a00", 156=>x"7800", 157=>x"7500", 158=>x"7800", 159=>x"7900", 160=>x"7d00", 161=>x"7c00",
---- 162=>x"7c00", 163=>x"7800", 164=>x"7500", 165=>x"8c00", 166=>x"7400", 167=>x"7300", 168=>x"7d00",
---- 169=>x"7900", 170=>x"7a00", 171=>x"7a00", 172=>x"7500", 173=>x"7600", 174=>x"7300", 175=>x"7300",
---- 176=>x"7d00", 177=>x"7a00", 178=>x"7c00", 179=>x"7a00", 180=>x"7600", 181=>x"7700", 182=>x"6f00",
---- 183=>x"7300", 184=>x"7b00", 185=>x"7e00", 186=>x"7d00", 187=>x"7800", 188=>x"7500", 189=>x"7300",
---- 190=>x"7300", 191=>x"7100", 192=>x"8100", 193=>x"7d00", 194=>x"7a00", 195=>x"7700", 196=>x"7900",
---- 197=>x"7700", 198=>x"7200", 199=>x"7100", 200=>x"7d00", 201=>x"7c00", 202=>x"7900", 203=>x"7700",
---- 204=>x"7800", 205=>x"7800", 206=>x"7500", 207=>x"6f00", 208=>x"7c00", 209=>x"7600", 210=>x"7700",
---- 211=>x"7900", 212=>x"7500", 213=>x"7500", 214=>x"7600", 215=>x"7100", 216=>x"7b00", 217=>x"7800",
---- 218=>x"7900", 219=>x"7800", 220=>x"8a00", 221=>x"7000", 222=>x"7400", 223=>x"7000", 224=>x"7b00",
---- 225=>x"7700", 226=>x"7600", 227=>x"7500", 228=>x"7400", 229=>x"7100", 230=>x"7300", 231=>x"6f00",
---- 232=>x"7700", 233=>x"7400", 234=>x"7100", 235=>x"7300", 236=>x"7100", 237=>x"7000", 238=>x"7000",
---- 239=>x"6f00", 240=>x"7800", 241=>x"7500", 242=>x"7300", 243=>x"7400", 244=>x"7300", 245=>x"7200",
---- 246=>x"7000", 247=>x"6d00", 248=>x"7700", 249=>x"7600", 250=>x"7500", 251=>x"7300", 252=>x"7100",
---- 253=>x"7100", 254=>x"6d00", 255=>x"6b00", 256=>x"7500", 257=>x"7400", 258=>x"7500", 259=>x"7200",
---- 260=>x"8f00", 261=>x"7100", 262=>x"7000", 263=>x"6f00", 264=>x"7400", 265=>x"7500", 266=>x"7400",
---- 267=>x"7100", 268=>x"7100", 269=>x"6f00", 270=>x"6e00", 271=>x"6f00", 272=>x"7300", 273=>x"7200",
---- 274=>x"7200", 275=>x"7100", 276=>x"6d00", 277=>x"6d00", 278=>x"6e00", 279=>x"6a00", 280=>x"7200",
---- 281=>x"7100", 282=>x"8d00", 283=>x"6f00", 284=>x"6f00", 285=>x"6f00", 286=>x"6e00", 287=>x"6a00",
---- 288=>x"7200", 289=>x"6e00", 290=>x"7000", 291=>x"6f00", 292=>x"6c00", 293=>x"6a00", 294=>x"6a00",
---- 295=>x"6c00", 296=>x"6e00", 297=>x"6c00", 298=>x"6e00", 299=>x"6d00", 300=>x"6b00", 301=>x"6a00",
---- 302=>x"6b00", 303=>x"6900", 304=>x"6c00", 305=>x"6c00", 306=>x"6c00", 307=>x"6b00", 308=>x"6a00",
---- 309=>x"6800", 310=>x"6700", 311=>x"6800", 312=>x"6600", 313=>x"9700", 314=>x"9600", 315=>x"6a00",
---- 316=>x"6500", 317=>x"6400", 318=>x"6500", 319=>x"6800", 320=>x"5d00", 321=>x"6200", 322=>x"6700",
---- 323=>x"6500", 324=>x"6400", 325=>x"6600", 326=>x"6400", 327=>x"6600", 328=>x"5900", 329=>x"5b00",
---- 330=>x"6400", 331=>x"6500", 332=>x"6700", 333=>x"6500", 334=>x"6500", 335=>x"6400", 336=>x"b000",
---- 337=>x"5700", 338=>x"5c00", 339=>x"6000", 340=>x"6000", 341=>x"6400", 342=>x"6200", 343=>x"6100",
---- 344=>x"5400", 345=>x"4e00", 346=>x"5400", 347=>x"5c00", 348=>x"5d00", 349=>x"6300", 350=>x"6100",
---- 351=>x"6100", 352=>x"9a00", 353=>x"4f00", 354=>x"4e00", 355=>x"5400", 356=>x"5900", 357=>x"5e00",
---- 358=>x"6200", 359=>x"6000", 360=>x"d500", 361=>x"7900", 362=>x"4800", 363=>x"5100", 364=>x"5500",
---- 365=>x"5800", 366=>x"5900", 367=>x"5c00", 368=>x"de00", 369=>x"bf00", 370=>x"6100", 371=>x"4800",
---- 372=>x"5000", 373=>x"5100", 374=>x"5400", 375=>x"5700", 376=>x"df00", 377=>x"e400", 378=>x"a200",
---- 379=>x"4d00", 380=>x"4b00", 381=>x"4a00", 382=>x"5000", 383=>x"5300", 384=>x"d900", 385=>x"de00",
---- 386=>x"d300", 387=>x"9b00", 388=>x"6700", 389=>x"5000", 390=>x"4d00", 391=>x"4c00", 392=>x"d600",
---- 393=>x"da00", 394=>x"e000", 395=>x"e200", 396=>x"cb00", 397=>x"9000", 398=>x"4b00", 399=>x"4600",
---- 400=>x"d600", 401=>x"d900", 402=>x"da00", 403=>x"de00", 404=>x"e600", 405=>x"db00", 406=>x"9400",
---- 407=>x"5f00", 408=>x"d300", 409=>x"d600", 410=>x"d500", 411=>x"d500", 412=>x"da00", 413=>x"e200",
---- 414=>x"df00", 415=>x"9600", 416=>x"d200", 417=>x"d600", 418=>x"d300", 419=>x"d300", 420=>x"d400",
---- 421=>x"da00", 422=>x"e100", 423=>x"d600", 424=>x"cd00", 425=>x"d600", 426=>x"d900", 427=>x"d700",
---- 428=>x"d800", 429=>x"da00", 430=>x"d600", 431=>x"e000", 432=>x"c900", 433=>x"cf00", 434=>x"d300",
---- 435=>x"d700", 436=>x"d700", 437=>x"dd00", 438=>x"dc00", 439=>x"dd00", 440=>x"cc00", 441=>x"d000",
---- 442=>x"d400", 443=>x"d700", 444=>x"d800", 445=>x"d800", 446=>x"df00", 447=>x"e100", 448=>x"cd00",
---- 449=>x"ce00", 450=>x"d200", 451=>x"d400", 452=>x"d500", 453=>x"d300", 454=>x"d900", 455=>x"df00",
---- 456=>x"d000", 457=>x"ca00", 458=>x"cf00", 459=>x"d300", 460=>x"d100", 461=>x"d500", 462=>x"d700",
---- 463=>x"df00", 464=>x"d300", 465=>x"cb00", 466=>x"cd00", 467=>x"d400", 468=>x"d100", 469=>x"d200",
---- 470=>x"d600", 471=>x"d800", 472=>x"cf00", 473=>x"d100", 474=>x"d100", 475=>x"d000", 476=>x"d000",
---- 477=>x"d200", 478=>x"d200", 479=>x"d400", 480=>x"ce00", 481=>x"ce00", 482=>x"cf00", 483=>x"cd00",
---- 484=>x"ca00", 485=>x"cc00", 486=>x"cd00", 487=>x"d200", 488=>x"cf00", 489=>x"cc00", 490=>x"ca00",
---- 491=>x"cc00", 492=>x"cd00", 493=>x"cb00", 494=>x"d000", 495=>x"cf00", 496=>x"ce00", 497=>x"d000",
---- 498=>x"cb00", 499=>x"d000", 500=>x"d100", 501=>x"d200", 502=>x"d100", 503=>x"d100", 504=>x"d100",
---- 505=>x"d100", 506=>x"cd00", 507=>x"ce00", 508=>x"cd00", 509=>x"cc00", 510=>x"cb00", 511=>x"cc00",
---- 512=>x"ca00", 513=>x"c600", 514=>x"c300", 515=>x"c700", 516=>x"c900", 517=>x"cb00", 518=>x"cc00",
---- 519=>x"ce00", 520=>x"c400", 521=>x"3f00", 522=>x"c500", 523=>x"cc00", 524=>x"cd00", 525=>x"ce00",
---- 526=>x"c900", 527=>x"cc00", 528=>x"cb00", 529=>x"c700", 530=>x"c600", 531=>x"cc00", 532=>x"ca00",
---- 533=>x"c900", 534=>x"c900", 535=>x"c800", 536=>x"c700", 537=>x"c800", 538=>x"c800", 539=>x"cd00",
---- 540=>x"c900", 541=>x"c800", 542=>x"cb00", 543=>x"c900", 544=>x"c400", 545=>x"c900", 546=>x"c900",
---- 547=>x"c900", 548=>x"c800", 549=>x"ca00", 550=>x"c900", 551=>x"c900", 552=>x"c600", 553=>x"c700",
---- 554=>x"c500", 555=>x"c600", 556=>x"c300", 557=>x"c800", 558=>x"c600", 559=>x"c700", 560=>x"c000",
---- 561=>x"c100", 562=>x"c000", 563=>x"c400", 564=>x"c300", 565=>x"c100", 566=>x"c500", 567=>x"c100",
---- 568=>x"c000", 569=>x"bf00", 570=>x"c000", 571=>x"c700", 572=>x"c700", 573=>x"c000", 574=>x"ba00",
---- 575=>x"c100", 576=>x"c400", 577=>x"c500", 578=>x"bf00", 579=>x"c400", 580=>x"c300", 581=>x"bc00",
---- 582=>x"b600", 583=>x"bb00", 584=>x"bc00", 585=>x"c300", 586=>x"bf00", 587=>x"b700", 588=>x"bb00",
---- 589=>x"b800", 590=>x"b600", 591=>x"b900", 592=>x"bd00", 593=>x"b900", 594=>x"bc00", 595=>x"b500",
---- 596=>x"af00", 597=>x"b100", 598=>x"b800", 599=>x"ba00", 600=>x"b900", 601=>x"b500", 602=>x"b100",
---- 603=>x"b100", 604=>x"b000", 605=>x"ab00", 606=>x"b300", 607=>x"ba00", 608=>x"b300", 609=>x"b700",
---- 610=>x"b900", 611=>x"ae00", 612=>x"aa00", 613=>x"b000", 614=>x"ac00", 615=>x"b500", 616=>x"b200",
---- 617=>x"b400", 618=>x"b400", 619=>x"b900", 620=>x"b500", 621=>x"ac00", 622=>x"b100", 623=>x"a800",
---- 624=>x"aa00", 625=>x"b400", 626=>x"b700", 627=>x"b600", 628=>x"b800", 629=>x"ac00", 630=>x"aa00",
---- 631=>x"a400", 632=>x"a700", 633=>x"a700", 634=>x"b200", 635=>x"b700", 636=>x"b100", 637=>x"ac00",
---- 638=>x"6100", 639=>x"a000", 640=>x"a700", 641=>x"a900", 642=>x"a700", 643=>x"b600", 644=>x"af00",
---- 645=>x"a500", 646=>x"9700", 647=>x"9800", 648=>x"a300", 649=>x"a600", 650=>x"a700", 651=>x"a500",
---- 652=>x"a600", 653=>x"9d00", 654=>x"a500", 655=>x"bc00", 656=>x"a900", 657=>x"9b00", 658=>x"9e00",
---- 659=>x"6a00", 660=>x"9900", 661=>x"b400", 662=>x"c600", 663=>x"be00", 664=>x"a500", 665=>x"9600",
---- 666=>x"9500", 667=>x"5300", 668=>x"bc00", 669=>x"c400", 670=>x"b300", 671=>x"aa00", 672=>x"9600",
---- 673=>x"a300", 674=>x"b500", 675=>x"c500", 676=>x"b800", 677=>x"aa00", 678=>x"b600", 679=>x"b500",
---- 680=>x"a600", 681=>x"c700", 682=>x"bf00", 683=>x"af00", 684=>x"a800", 685=>x"b100", 686=>x"c200",
---- 687=>x"c300", 688=>x"c600", 689=>x"b900", 690=>x"a800", 691=>x"aa00", 692=>x"bb00", 693=>x"c100",
---- 694=>x"c400", 695=>x"c900", 696=>x"ab00", 697=>x"a500", 698=>x"ab00", 699=>x"c000", 700=>x"ca00",
---- 701=>x"cd00", 702=>x"ca00", 703=>x"c600", 704=>x"a000", 705=>x"ac00", 706=>x"bd00", 707=>x"bd00",
---- 708=>x"c400", 709=>x"c900", 710=>x"c700", 711=>x"c100", 712=>x"b200", 713=>x"c500", 714=>x"c900",
---- 715=>x"c200", 716=>x"c400", 717=>x"c600", 718=>x"c300", 719=>x"be00", 720=>x"c500", 721=>x"c900",
---- 722=>x"c800", 723=>x"c300", 724=>x"c600", 725=>x"c400", 726=>x"c100", 727=>x"c100", 728=>x"ca00",
---- 729=>x"c500", 730=>x"c400", 731=>x"c100", 732=>x"c100", 733=>x"c000", 734=>x"c000", 735=>x"c100",
---- 736=>x"c600", 737=>x"c500", 738=>x"c500", 739=>x"c200", 740=>x"c000", 741=>x"c200", 742=>x"c000",
---- 743=>x"c000", 744=>x"3e00", 745=>x"c400", 746=>x"c400", 747=>x"c000", 748=>x"c100", 749=>x"c200",
---- 750=>x"be00", 751=>x"c000", 752=>x"bf00", 753=>x"c200", 754=>x"c100", 755=>x"be00", 756=>x"be00",
---- 757=>x"3c00", 758=>x"bb00", 759=>x"b900", 760=>x"bf00", 761=>x"bf00", 762=>x"bc00", 763=>x"be00",
---- 764=>x"bf00", 765=>x"bc00", 766=>x"ba00", 767=>x"bc00", 768=>x"bc00", 769=>x"bc00", 770=>x"bc00",
---- 771=>x"bd00", 772=>x"bd00", 773=>x"b900", 774=>x"bb00", 775=>x"bb00", 776=>x"b800", 777=>x"4600",
---- 778=>x"b800", 779=>x"b900", 780=>x"bb00", 781=>x"b600", 782=>x"b800", 783=>x"bc00", 784=>x"b500",
---- 785=>x"b400", 786=>x"b300", 787=>x"b500", 788=>x"b500", 789=>x"b700", 790=>x"b800", 791=>x"b900",
---- 792=>x"b500", 793=>x"b300", 794=>x"b300", 795=>x"b300", 796=>x"af00", 797=>x"b200", 798=>x"b900",
---- 799=>x"bc00", 800=>x"b500", 801=>x"af00", 802=>x"b000", 803=>x"b300", 804=>x"ae00", 805=>x"af00",
---- 806=>x"b700", 807=>x"bf00", 808=>x"b000", 809=>x"ad00", 810=>x"ac00", 811=>x"b400", 812=>x"b700",
---- 813=>x"af00", 814=>x"b600", 815=>x"bd00", 816=>x"aa00", 817=>x"a700", 818=>x"ae00", 819=>x"b700",
---- 820=>x"b400", 821=>x"b400", 822=>x"b600", 823=>x"bd00", 824=>x"aa00", 825=>x"ab00", 826=>x"b300",
---- 827=>x"b800", 828=>x"b600", 829=>x"b600", 830=>x"ba00", 831=>x"ba00", 832=>x"b000", 833=>x"5200",
---- 834=>x"b500", 835=>x"b900", 836=>x"4700", 837=>x"b600", 838=>x"b800", 839=>x"b600", 840=>x"b000",
---- 841=>x"ac00", 842=>x"b300", 843=>x"b300", 844=>x"b300", 845=>x"b400", 846=>x"bb00", 847=>x"bf00",
---- 848=>x"ae00", 849=>x"b100", 850=>x"ab00", 851=>x"ac00", 852=>x"b600", 853=>x"c000", 854=>x"c600",
---- 855=>x"c100", 856=>x"b000", 857=>x"a700", 858=>x"a600", 859=>x"b800", 860=>x"c200", 861=>x"c400",
---- 862=>x"c800", 863=>x"c300", 864=>x"a700", 865=>x"ab00", 866=>x"bb00", 867=>x"c400", 868=>x"c400",
---- 869=>x"c500", 870=>x"cb00", 871=>x"c500", 872=>x"b200", 873=>x"bb00", 874=>x"bd00", 875=>x"c300",
---- 876=>x"c500", 877=>x"c400", 878=>x"cc00", 879=>x"c800", 880=>x"b800", 881=>x"b900", 882=>x"bc00",
---- 883=>x"c500", 884=>x"c200", 885=>x"3a00", 886=>x"c900", 887=>x"c800", 888=>x"b800", 889=>x"bd00",
---- 890=>x"c000", 891=>x"c400", 892=>x"c300", 893=>x"c500", 894=>x"ca00", 895=>x"ca00", 896=>x"b800",
---- 897=>x"c100", 898=>x"c300", 899=>x"c800", 900=>x"c600", 901=>x"c700", 902=>x"cb00", 903=>x"ca00",
---- 904=>x"ba00", 905=>x"bf00", 906=>x"c000", 907=>x"c500", 908=>x"c500", 909=>x"c700", 910=>x"c900",
---- 911=>x"c900", 912=>x"bc00", 913=>x"be00", 914=>x"c300", 915=>x"c600", 916=>x"c800", 917=>x"c600",
---- 918=>x"c900", 919=>x"cb00", 920=>x"c000", 921=>x"c300", 922=>x"c300", 923=>x"c400", 924=>x"c800",
---- 925=>x"c900", 926=>x"c900", 927=>x"cd00", 928=>x"c100", 929=>x"c300", 930=>x"c400", 931=>x"c500",
---- 932=>x"c400", 933=>x"c900", 934=>x"cb00", 935=>x"cc00", 936=>x"c000", 937=>x"c100", 938=>x"3d00",
---- 939=>x"c600", 940=>x"c600", 941=>x"c600", 942=>x"cc00", 943=>x"cc00", 944=>x"bf00", 945=>x"c300",
---- 946=>x"c400", 947=>x"c400", 948=>x"c800", 949=>x"c700", 950=>x"c800", 951=>x"ca00", 952=>x"be00",
---- 953=>x"bf00", 954=>x"c400", 955=>x"c600", 956=>x"c500", 957=>x"c600", 958=>x"c500", 959=>x"c500",
---- 960=>x"bb00", 961=>x"bd00", 962=>x"c100", 963=>x"c500", 964=>x"c600", 965=>x"c400", 966=>x"c200",
---- 967=>x"c500", 968=>x"b700", 969=>x"ba00", 970=>x"be00", 971=>x"c200", 972=>x"c500", 973=>x"c300",
---- 974=>x"c300", 975=>x"c400", 976=>x"b500", 977=>x"b800", 978=>x"bc00", 979=>x"c300", 980=>x"c400",
---- 981=>x"c400", 982=>x"c200", 983=>x"bf00", 984=>x"af00", 985=>x"b700", 986=>x"b900", 987=>x"be00",
---- 988=>x"c200", 989=>x"c200", 990=>x"bd00", 991=>x"be00", 992=>x"ad00", 993=>x"b000", 994=>x"b900",
---- 995=>x"bf00", 996=>x"c200", 997=>x"c200", 998=>x"be00", 999=>x"4400", 1000=>x"af00", 1001=>x"b100",
---- 1002=>x"b800", 1003=>x"bd00", 1004=>x"bf00", 1005=>x"c000", 1006=>x"be00", 1007=>x"ba00", 1008=>x"aa00",
---- 1009=>x"b000", 1010=>x"b500", 1011=>x"bb00", 1012=>x"c000", 1013=>x"bf00", 1014=>x"bf00", 1015=>x"bc00",
---- 1016=>x"a300", 1017=>x"aa00", 1018=>x"b500", 1019=>x"bb00", 1020=>x"c100", 1021=>x"c400", 1022=>x"c100",
---- 1023=>x"bc00", 1024=>x"9f00", 1025=>x"5800", 1026=>x"b200", 1027=>x"c000", 1028=>x"c200", 1029=>x"c400",
---- 1030=>x"c300", 1031=>x"be00", 1032=>x"9d00", 1033=>x"a500", 1034=>x"b200", 1035=>x"be00", 1036=>x"c200",
---- 1037=>x"c300", 1038=>x"c700", 1039=>x"c600", 1040=>x"9d00", 1041=>x"a500", 1042=>x"b300", 1043=>x"be00",
---- 1044=>x"c700", 1045=>x"ca00", 1046=>x"cb00", 1047=>x"c900", 1048=>x"9a00", 1049=>x"a400", 1050=>x"b300",
---- 1051=>x"bf00", 1052=>x"cc00", 1053=>x"cf00", 1054=>x"cf00", 1055=>x"cd00", 1056=>x"9a00", 1057=>x"a300",
---- 1058=>x"ae00", 1059=>x"c400", 1060=>x"d100", 1061=>x"d600", 1062=>x"d700", 1063=>x"af00", 1064=>x"6700",
---- 1065=>x"a500", 1066=>x"b400", 1067=>x"c800", 1068=>x"d700", 1069=>x"dc00", 1070=>x"c700", 1071=>x"7300",
---- 1072=>x"9b00", 1073=>x"a700", 1074=>x"b800", 1075=>x"ca00", 1076=>x"d700", 1077=>x"d900", 1078=>x"a700",
---- 1079=>x"5a00", 1080=>x"9d00", 1081=>x"a900", 1082=>x"bc00", 1083=>x"d400", 1084=>x"da00", 1085=>x"d500",
---- 1086=>x"8b00", 1087=>x"6400", 1088=>x"9800", 1089=>x"ab00", 1090=>x"c500", 1091=>x"da00", 1092=>x"dd00",
---- 1093=>x"cb00", 1094=>x"7f00", 1095=>x"5e00", 1096=>x"9b00", 1097=>x"ad00", 1098=>x"c400", 1099=>x"db00",
---- 1100=>x"df00", 1101=>x"c500", 1102=>x"8800", 1103=>x"6500", 1104=>x"9600", 1105=>x"a800", 1106=>x"c100",
---- 1107=>x"da00", 1108=>x"e000", 1109=>x"c700", 1110=>x"aa00", 1111=>x"a100", 1112=>x"9400", 1113=>x"a300",
---- 1114=>x"bb00", 1115=>x"d900", 1116=>x"e000", 1117=>x"cc00", 1118=>x"ab00", 1119=>x"a200", 1120=>x"9200",
---- 1121=>x"a400", 1122=>x"ba00", 1123=>x"d600", 1124=>x"e200", 1125=>x"d000", 1126=>x"b200", 1127=>x"9f00",
---- 1128=>x"8e00", 1129=>x"a500", 1130=>x"bb00", 1131=>x"d200", 1132=>x"df00", 1133=>x"d400", 1134=>x"bb00",
---- 1135=>x"b000", 1136=>x"8e00", 1137=>x"a200", 1138=>x"b600", 1139=>x"cf00", 1140=>x"de00", 1141=>x"d600",
---- 1142=>x"bf00", 1143=>x"ba00", 1144=>x"8a00", 1145=>x"a200", 1146=>x"b500", 1147=>x"3100", 1148=>x"de00",
---- 1149=>x"d700", 1150=>x"c100", 1151=>x"b800", 1152=>x"8700", 1153=>x"9a00", 1154=>x"b500", 1155=>x"cc00",
---- 1156=>x"db00", 1157=>x"db00", 1158=>x"c300", 1159=>x"b600", 1160=>x"8300", 1161=>x"9800", 1162=>x"b000",
---- 1163=>x"c900", 1164=>x"dc00", 1165=>x"de00", 1166=>x"c900", 1167=>x"b600", 1168=>x"8500", 1169=>x"9200",
---- 1170=>x"a900", 1171=>x"c900", 1172=>x"dd00", 1173=>x"dc00", 1174=>x"cd00", 1175=>x"b700", 1176=>x"8100",
---- 1177=>x"6e00", 1178=>x"ab00", 1179=>x"c800", 1180=>x"d900", 1181=>x"dc00", 1182=>x"d000", 1183=>x"ba00",
---- 1184=>x"8400", 1185=>x"9300", 1186=>x"a400", 1187=>x"c400", 1188=>x"dc00", 1189=>x"e000", 1190=>x"d400",
---- 1191=>x"b800", 1192=>x"8600", 1193=>x"8f00", 1194=>x"a300", 1195=>x"c000", 1196=>x"d900", 1197=>x"df00",
---- 1198=>x"d500", 1199=>x"b900", 1200=>x"8600", 1201=>x"9100", 1202=>x"a100", 1203=>x"bc00", 1204=>x"d600",
---- 1205=>x"df00", 1206=>x"d900", 1207=>x"bc00", 1208=>x"8400", 1209=>x"9000", 1210=>x"9d00", 1211=>x"b000",
---- 1212=>x"cd00", 1213=>x"df00", 1214=>x"dc00", 1215=>x"be00", 1216=>x"8600", 1217=>x"8c00", 1218=>x"9800",
---- 1219=>x"ac00", 1220=>x"ca00", 1221=>x"dd00", 1222=>x"dc00", 1223=>x"c400", 1224=>x"8200", 1225=>x"8600",
---- 1226=>x"9900", 1227=>x"af00", 1228=>x"c900", 1229=>x"db00", 1230=>x"df00", 1231=>x"cb00", 1232=>x"7e00",
---- 1233=>x"8800", 1234=>x"9800", 1235=>x"ac00", 1236=>x"c200", 1237=>x"d500", 1238=>x"e300", 1239=>x"d600",
---- 1240=>x"7e00", 1241=>x"8800", 1242=>x"9400", 1243=>x"a400", 1244=>x"b800", 1245=>x"d400", 1246=>x"e500",
---- 1247=>x"dd00", 1248=>x"7f00", 1249=>x"8600", 1250=>x"9300", 1251=>x"a200", 1252=>x"b200", 1253=>x"d200",
---- 1254=>x"e400", 1255=>x"df00", 1256=>x"7f00", 1257=>x"8700", 1258=>x"9000", 1259=>x"a100", 1260=>x"ae00",
---- 1261=>x"cc00", 1262=>x"e600", 1263=>x"1d00", 1264=>x"7f00", 1265=>x"8700", 1266=>x"8d00", 1267=>x"a100",
---- 1268=>x"b300", 1269=>x"cb00", 1270=>x"e700", 1271=>x"e300", 1272=>x"7900", 1273=>x"7c00", 1274=>x"8a00",
---- 1275=>x"9e00", 1276=>x"b500", 1277=>x"c800", 1278=>x"dd00", 1279=>x"e000", 1280=>x"7900", 1281=>x"7600",
---- 1282=>x"8400", 1283=>x"9600", 1284=>x"ac00", 1285=>x"c500", 1286=>x"cf00", 1287=>x"d400", 1288=>x"7a00",
---- 1289=>x"7b00", 1290=>x"7d00", 1291=>x"8500", 1292=>x"a100", 1293=>x"bc00", 1294=>x"cc00", 1295=>x"bc00",
---- 1296=>x"5c00", 1297=>x"6d00", 1298=>x"7900", 1299=>x"7e00", 1300=>x"9300", 1301=>x"b100", 1302=>x"c300",
---- 1303=>x"ac00", 1304=>x"6a00", 1305=>x"6500", 1306=>x"7300", 1307=>x"7700", 1308=>x"8900", 1309=>x"b200",
---- 1310=>x"b800", 1311=>x"aa00", 1312=>x"7600", 1313=>x"7d00", 1314=>x"8b00", 1315=>x"9c00", 1316=>x"b100",
---- 1317=>x"be00", 1318=>x"b300", 1319=>x"a600", 1320=>x"8400", 1321=>x"9a00", 1322=>x"bb00", 1323=>x"c800",
---- 1324=>x"c400", 1325=>x"be00", 1326=>x"b000", 1327=>x"a700", 1328=>x"9a00", 1329=>x"a000", 1330=>x"be00",
---- 1331=>x"c600", 1332=>x"c000", 1333=>x"bf00", 1334=>x"b300", 1335=>x"a600", 1336=>x"a900", 1337=>x"a600",
---- 1338=>x"bf00", 1339=>x"c700", 1340=>x"c000", 1341=>x"c100", 1342=>x"b200", 1343=>x"a200", 1344=>x"b500",
---- 1345=>x"aa00", 1346=>x"c200", 1347=>x"c800", 1348=>x"c500", 1349=>x"c500", 1350=>x"b100", 1351=>x"a000",
---- 1352=>x"bd00", 1353=>x"ac00", 1354=>x"c200", 1355=>x"ce00", 1356=>x"c500", 1357=>x"c000", 1358=>x"af00",
---- 1359=>x"a000", 1360=>x"c000", 1361=>x"a900", 1362=>x"b900", 1363=>x"cd00", 1364=>x"c700", 1365=>x"be00",
---- 1366=>x"b000", 1367=>x"9b00", 1368=>x"c300", 1369=>x"b200", 1370=>x"c800", 1371=>x"d200", 1372=>x"cb00",
---- 1373=>x"c300", 1374=>x"b400", 1375=>x"9800", 1376=>x"c500", 1377=>x"cc00", 1378=>x"c000", 1379=>x"b400",
---- 1380=>x"ac00", 1381=>x"b500", 1382=>x"b400", 1383=>x"9300", 1384=>x"9a00", 1385=>x"a600", 1386=>x"9b00",
---- 1387=>x"9600", 1388=>x"9200", 1389=>x"9b00", 1390=>x"9900", 1391=>x"7b00", 1392=>x"8900", 1393=>x"8d00",
---- 1394=>x"7800", 1395=>x"6600", 1396=>x"7200", 1397=>x"7900", 1398=>x"6a00", 1399=>x"6000", 1400=>x"7c00",
---- 1401=>x"7400", 1402=>x"5b00", 1403=>x"5200", 1404=>x"5f00", 1405=>x"6f00", 1406=>x"7000", 1407=>x"7300",
---- 1408=>x"8000", 1409=>x"8100", 1410=>x"8300", 1411=>x"7b00", 1412=>x"7900", 1413=>x"8700", 1414=>x"8500",
---- 1415=>x"8500", 1416=>x"b100", 1417=>x"b400", 1418=>x"a200", 1419=>x"8900", 1420=>x"8600", 1421=>x"8d00",
---- 1422=>x"9000", 1423=>x"9000", 1424=>x"c800", 1425=>x"c400", 1426=>x"a000", 1427=>x"8700", 1428=>x"8800",
---- 1429=>x"8f00", 1430=>x"9500", 1431=>x"8f00", 1432=>x"a400", 1433=>x"a600", 1434=>x"8f00", 1435=>x"8700",
---- 1436=>x"9000", 1437=>x"9300", 1438=>x"9700", 1439=>x"8e00", 1440=>x"8f00", 1441=>x"8e00", 1442=>x"8400",
---- 1443=>x"8e00", 1444=>x"9300", 1445=>x"9700", 1446=>x"8f00", 1447=>x"8b00", 1448=>x"8100", 1449=>x"8200",
---- 1450=>x"8d00", 1451=>x"9700", 1452=>x"9300", 1453=>x"9300", 1454=>x"8d00", 1455=>x"7900", 1456=>x"8000",
---- 1457=>x"9400", 1458=>x"9a00", 1459=>x"9300", 1460=>x"8f00", 1461=>x"9000", 1462=>x"8000", 1463=>x"4e00",
---- 1464=>x"9600", 1465=>x"9b00", 1466=>x"9600", 1467=>x"8c00", 1468=>x"8d00", 1469=>x"9100", 1470=>x"5c00",
---- 1471=>x"3c00", 1472=>x"9800", 1473=>x"9900", 1474=>x"8d00", 1475=>x"8b00", 1476=>x"9000", 1477=>x"8200",
---- 1478=>x"3500", 1479=>x"3f00", 1480=>x"9b00", 1481=>x"9600", 1482=>x"9000", 1483=>x"9000", 1484=>x"9200",
---- 1485=>x"5c00", 1486=>x"d700", 1487=>x"4800", 1488=>x"9b00", 1489=>x"9600", 1490=>x"9200", 1491=>x"9500",
---- 1492=>x"8600", 1493=>x"3300", 1494=>x"2800", 1495=>x"4000", 1496=>x"9c00", 1497=>x"9600", 1498=>x"9500",
---- 1499=>x"9800", 1500=>x"6c00", 1501=>x"2500", 1502=>x"3100", 1503=>x"4400", 1504=>x"9900", 1505=>x"9100",
---- 1506=>x"9800", 1507=>x"6c00", 1508=>x"4c00", 1509=>x"2500", 1510=>x"3a00", 1511=>x"4500", 1512=>x"9700",
---- 1513=>x"9100", 1514=>x"9900", 1515=>x"8000", 1516=>x"3700", 1517=>x"2700", 1518=>x"3e00", 1519=>x"3c00",
---- 1520=>x"9400", 1521=>x"9400", 1522=>x"9100", 1523=>x"6f00", 1524=>x"3200", 1525=>x"2900", 1526=>x"3f00",
---- 1527=>x"3500", 1528=>x"9400", 1529=>x"9100", 1530=>x"8a00", 1531=>x"6e00", 1532=>x"3500", 1533=>x"2b00",
---- 1534=>x"3d00", 1535=>x"3700", 1536=>x"8e00", 1537=>x"8900", 1538=>x"8600", 1539=>x"6100", 1540=>x"3300",
---- 1541=>x"2e00", 1542=>x"3700", 1543=>x"3700", 1544=>x"8200", 1545=>x"8400", 1546=>x"7d00", 1547=>x"5500",
---- 1548=>x"3200", 1549=>x"3200", 1550=>x"3400", 1551=>x"3600", 1552=>x"9e00", 1553=>x"a300", 1554=>x"9700",
---- 1555=>x"7100", 1556=>x"4400", 1557=>x"3900", 1558=>x"3300", 1559=>x"3800", 1560=>x"4600", 1561=>x"bf00",
---- 1562=>x"c400", 1563=>x"bd00", 1564=>x"a900", 1565=>x"8900", 1566=>x"a100", 1567=>x"4100", 1568=>x"b300",
---- 1569=>x"bf00", 1570=>x"c300", 1571=>x"c700", 1572=>x"cc00", 1573=>x"cb00", 1574=>x"c000", 1575=>x"a000",
---- 1576=>x"b700", 1577=>x"bf00", 1578=>x"c400", 1579=>x"c500", 1580=>x"c600", 1581=>x"c800", 1582=>x"cd00",
---- 1583=>x"d000", 1584=>x"b700", 1585=>x"bf00", 1586=>x"c300", 1587=>x"c500", 1588=>x"c800", 1589=>x"c800",
---- 1590=>x"c900", 1591=>x"c900", 1592=>x"bb00", 1593=>x"bd00", 1594=>x"c200", 1595=>x"c400", 1596=>x"c800",
---- 1597=>x"c700", 1598=>x"c900", 1599=>x"c800", 1600=>x"bc00", 1601=>x"bf00", 1602=>x"c100", 1603=>x"c200",
---- 1604=>x"c300", 1605=>x"c400", 1606=>x"c900", 1607=>x"c800", 1608=>x"ba00", 1609=>x"bd00", 1610=>x"be00",
---- 1611=>x"be00", 1612=>x"be00", 1613=>x"c100", 1614=>x"c500", 1615=>x"c500", 1616=>x"b900", 1617=>x"bd00",
---- 1618=>x"be00", 1619=>x"bd00", 1620=>x"bd00", 1621=>x"c200", 1622=>x"c300", 1623=>x"c200", 1624=>x"b900",
---- 1625=>x"bd00", 1626=>x"ba00", 1627=>x"bc00", 1628=>x"4100", 1629=>x"c000", 1630=>x"c000", 1631=>x"c100",
---- 1632=>x"b400", 1633=>x"b700", 1634=>x"b900", 1635=>x"b900", 1636=>x"be00", 1637=>x"be00", 1638=>x"be00",
---- 1639=>x"bd00", 1640=>x"b300", 1641=>x"b400", 1642=>x"b500", 1643=>x"b800", 1644=>x"ba00", 1645=>x"bb00",
---- 1646=>x"bd00", 1647=>x"bf00", 1648=>x"af00", 1649=>x"b000", 1650=>x"b400", 1651=>x"b300", 1652=>x"b400",
---- 1653=>x"bb00", 1654=>x"bd00", 1655=>x"bd00", 1656=>x"af00", 1657=>x"ac00", 1658=>x"af00", 1659=>x"b100",
---- 1660=>x"b300", 1661=>x"b500", 1662=>x"b900", 1663=>x"b800", 1664=>x"ad00", 1665=>x"b000", 1666=>x"ad00",
---- 1667=>x"b000", 1668=>x"b300", 1669=>x"b500", 1670=>x"b700", 1671=>x"b600", 1672=>x"a800", 1673=>x"ae00",
---- 1674=>x"ad00", 1675=>x"ae00", 1676=>x"b300", 1677=>x"b400", 1678=>x"b500", 1679=>x"ba00", 1680=>x"a900",
---- 1681=>x"ac00", 1682=>x"ad00", 1683=>x"ad00", 1684=>x"b200", 1685=>x"b100", 1686=>x"b500", 1687=>x"b900",
---- 1688=>x"a500", 1689=>x"a800", 1690=>x"aa00", 1691=>x"ad00", 1692=>x"b100", 1693=>x"b200", 1694=>x"b700",
---- 1695=>x"b700", 1696=>x"a500", 1697=>x"a900", 1698=>x"ab00", 1699=>x"ad00", 1700=>x"af00", 1701=>x"b200",
---- 1702=>x"b600", 1703=>x"b300", 1704=>x"a400", 1705=>x"a700", 1706=>x"ac00", 1707=>x"ac00", 1708=>x"af00",
---- 1709=>x"b200", 1710=>x"b100", 1711=>x"b500", 1712=>x"a300", 1713=>x"a700", 1714=>x"aa00", 1715=>x"aa00",
---- 1716=>x"af00", 1717=>x"af00", 1718=>x"b000", 1719=>x"b900", 1720=>x"a600", 1721=>x"a600", 1722=>x"a700",
---- 1723=>x"aa00", 1724=>x"ab00", 1725=>x"af00", 1726=>x"b200", 1727=>x"b300", 1728=>x"a300", 1729=>x"a600",
---- 1730=>x"a600", 1731=>x"a800", 1732=>x"ac00", 1733=>x"ad00", 1734=>x"4f00", 1735=>x"b400", 1736=>x"a200",
---- 1737=>x"a400", 1738=>x"a400", 1739=>x"a600", 1740=>x"ab00", 1741=>x"b000", 1742=>x"af00", 1743=>x"b100",
---- 1744=>x"a100", 1745=>x"a300", 1746=>x"a300", 1747=>x"5900", 1748=>x"ab00", 1749=>x"b000", 1750=>x"ac00",
---- 1751=>x"b100", 1752=>x"9f00", 1753=>x"a100", 1754=>x"a300", 1755=>x"a500", 1756=>x"a700", 1757=>x"ac00",
---- 1758=>x"af00", 1759=>x"b200", 1760=>x"9e00", 1761=>x"a100", 1762=>x"a300", 1763=>x"a400", 1764=>x"a800",
---- 1765=>x"ab00", 1766=>x"b100", 1767=>x"b200", 1768=>x"9f00", 1769=>x"a000", 1770=>x"a000", 1771=>x"a300",
---- 1772=>x"a500", 1773=>x"a900", 1774=>x"aa00", 1775=>x"ac00", 1776=>x"9b00", 1777=>x"9f00", 1778=>x"5f00",
---- 1779=>x"a200", 1780=>x"a600", 1781=>x"aa00", 1782=>x"a800", 1783=>x"a900", 1784=>x"9e00", 1785=>x"9c00",
---- 1786=>x"9d00", 1787=>x"a100", 1788=>x"a700", 1789=>x"a700", 1790=>x"a900", 1791=>x"aa00", 1792=>x"9f00",
---- 1793=>x"9e00", 1794=>x"9d00", 1795=>x"a100", 1796=>x"a400", 1797=>x"a700", 1798=>x"a700", 1799=>x"ad00",
---- 1800=>x"6400", 1801=>x"9c00", 1802=>x"a000", 1803=>x"a300", 1804=>x"a400", 1805=>x"a700", 1806=>x"a500",
---- 1807=>x"a900", 1808=>x"9b00", 1809=>x"9c00", 1810=>x"9f00", 1811=>x"a100", 1812=>x"a400", 1813=>x"a600",
---- 1814=>x"a700", 1815=>x"a500", 1816=>x"9a00", 1817=>x"9b00", 1818=>x"9d00", 1819=>x"9e00", 1820=>x"a100",
---- 1821=>x"a500", 1822=>x"a400", 1823=>x"a600", 1824=>x"9800", 1825=>x"9a00", 1826=>x"9b00", 1827=>x"9f00",
---- 1828=>x"9c00", 1829=>x"a200", 1830=>x"a300", 1831=>x"a500", 1832=>x"9800", 1833=>x"9800", 1834=>x"9a00",
---- 1835=>x"9c00", 1836=>x"9d00", 1837=>x"9f00", 1838=>x"a000", 1839=>x"a500", 1840=>x"9600", 1841=>x"9900",
---- 1842=>x"9900", 1843=>x"9b00", 1844=>x"9d00", 1845=>x"a100", 1846=>x"a300", 1847=>x"a500", 1848=>x"9a00",
---- 1849=>x"9a00", 1850=>x"9900", 1851=>x"9800", 1852=>x"a000", 1853=>x"a200", 1854=>x"a100", 1855=>x"a400",
---- 1856=>x"9500", 1857=>x"9700", 1858=>x"9900", 1859=>x"9d00", 1860=>x"9d00", 1861=>x"9f00", 1862=>x"a000",
---- 1863=>x"a300", 1864=>x"9300", 1865=>x"9800", 1866=>x"9900", 1867=>x"9b00", 1868=>x"6300", 1869=>x"9f00",
---- 1870=>x"6000", 1871=>x"a200", 1872=>x"9400", 1873=>x"9600", 1874=>x"9700", 1875=>x"9700", 1876=>x"9a00",
---- 1877=>x"9f00", 1878=>x"a000", 1879=>x"a100", 1880=>x"9400", 1881=>x"9500", 1882=>x"9600", 1883=>x"9600",
---- 1884=>x"9900", 1885=>x"9b00", 1886=>x"9e00", 1887=>x"9d00", 1888=>x"9500", 1889=>x"9700", 1890=>x"9600",
---- 1891=>x"9900", 1892=>x"9c00", 1893=>x"9b00", 1894=>x"9c00", 1895=>x"9f00", 1896=>x"9200", 1897=>x"9300",
---- 1898=>x"9400", 1899=>x"9900", 1900=>x"9a00", 1901=>x"6400", 1902=>x"9d00", 1903=>x"9d00", 1904=>x"9100",
---- 1905=>x"9200", 1906=>x"9200", 1907=>x"9400", 1908=>x"9a00", 1909=>x"9b00", 1910=>x"9d00", 1911=>x"9b00",
---- 1912=>x"9000", 1913=>x"9300", 1914=>x"9100", 1915=>x"9300", 1916=>x"9800", 1917=>x"6600", 1918=>x"9b00",
---- 1919=>x"9b00", 1920=>x"8f00", 1921=>x"9200", 1922=>x"9100", 1923=>x"9500", 1924=>x"9800", 1925=>x"9700",
---- 1926=>x"9800", 1927=>x"9c00", 1928=>x"9100", 1929=>x"9000", 1930=>x"9100", 1931=>x"9300", 1932=>x"9400",
---- 1933=>x"9500", 1934=>x"9700", 1935=>x"9a00", 1936=>x"9000", 1937=>x"9100", 1938=>x"9000", 1939=>x"9200",
---- 1940=>x"9400", 1941=>x"9300", 1942=>x"9800", 1943=>x"9a00", 1944=>x"8d00", 1945=>x"8e00", 1946=>x"8f00",
---- 1947=>x"9500", 1948=>x"9400", 1949=>x"9200", 1950=>x"9500", 1951=>x"9a00", 1952=>x"8a00", 1953=>x"8e00",
---- 1954=>x"9000", 1955=>x"9000", 1956=>x"9400", 1957=>x"9300", 1958=>x"9600", 1959=>x"9700", 1960=>x"8c00",
---- 1961=>x"8d00", 1962=>x"9100", 1963=>x"8e00", 1964=>x"9100", 1965=>x"9600", 1966=>x"9500", 1967=>x"9700",
---- 1968=>x"8d00", 1969=>x"8d00", 1970=>x"8e00", 1971=>x"9000", 1972=>x"9100", 1973=>x"9300", 1974=>x"9500",
---- 1975=>x"9600", 1976=>x"8e00", 1977=>x"8c00", 1978=>x"8f00", 1979=>x"8d00", 1980=>x"9100", 1981=>x"9500",
---- 1982=>x"9700", 1983=>x"9700", 1984=>x"8d00", 1985=>x"8f00", 1986=>x"9000", 1987=>x"8e00", 1988=>x"9100",
---- 1989=>x"9300", 1990=>x"9400", 1991=>x"9400", 1992=>x"8e00", 1993=>x"9100", 1994=>x"9100", 1995=>x"9200",
---- 1996=>x"9300", 1997=>x"9400", 1998=>x"9200", 1999=>x"9700", 2000=>x"8f00", 2001=>x"9200", 2002=>x"9200",
---- 2003=>x"9200", 2004=>x"9300", 2005=>x"9400", 2006=>x"9400", 2007=>x"6900", 2008=>x"9200", 2009=>x"9300",
---- 2010=>x"9200", 2011=>x"9000", 2012=>x"9500", 2013=>x"9500", 2014=>x"9400", 2015=>x"9600", 2016=>x"9300",
---- 2017=>x"9300", 2018=>x"9200", 2019=>x"9200", 2020=>x"9300", 2021=>x"9700", 2022=>x"9600", 2023=>x"9b00",
---- 2024=>x"9400", 2025=>x"9400", 2026=>x"9100", 2027=>x"9200", 2028=>x"9300", 2029=>x"9600", 2030=>x"9600",
---- 2031=>x"9b00", 2032=>x"9300", 2033=>x"9500", 2034=>x"9600", 2035=>x"9100", 2036=>x"9400", 2037=>x"9600",
---- 2038=>x"9500", 2039=>x"9500", 2040=>x"9500", 2041=>x"9600", 2042=>x"9700", 2043=>x"9300", 2044=>x"9700",
---- 2045=>x"9600", 2046=>x"9700", 2047=>x"9600"),
---- 20 => (0=>x"6900", 1=>x"7400", 2=>x"7b00", 3=>x"8800", 4=>x"8e00", 5=>x"9200", 6=>x"9800", 7=>x"9a00",
---- 8=>x"6900", 9=>x"7400", 10=>x"7b00", 11=>x"8800", 12=>x"8d00", 13=>x"9200", 14=>x"9800",
---- 15=>x"9a00", 16=>x"6900", 17=>x"7300", 18=>x"7c00", 19=>x"8600", 20=>x"8c00", 21=>x"9300",
---- 22=>x"9700", 23=>x"9900", 24=>x"6500", 25=>x"6f00", 26=>x"7b00", 27=>x"8000", 28=>x"8900",
---- 29=>x"9100", 30=>x"9400", 31=>x"9900", 32=>x"6500", 33=>x"6a00", 34=>x"7200", 35=>x"7b00",
---- 36=>x"8500", 37=>x"8c00", 38=>x"9300", 39=>x"9800", 40=>x"6b00", 41=>x"6700", 42=>x"6c00",
---- 43=>x"7400", 44=>x"7f00", 45=>x"8800", 46=>x"8e00", 47=>x"9600", 48=>x"6d00", 49=>x"6a00",
---- 50=>x"6600", 51=>x"9000", 52=>x"7c00", 53=>x"8700", 54=>x"8d00", 55=>x"9300", 56=>x"6e00",
---- 57=>x"6b00", 58=>x"6600", 59=>x"6c00", 60=>x"7400", 61=>x"8100", 62=>x"8d00", 63=>x"9200",
---- 64=>x"6e00", 65=>x"6b00", 66=>x"6a00", 67=>x"6900", 68=>x"6f00", 69=>x"7b00", 70=>x"8a00",
---- 71=>x"9200", 72=>x"6f00", 73=>x"6f00", 74=>x"6800", 75=>x"6500", 76=>x"6d00", 77=>x"7900",
---- 78=>x"8400", 79=>x"8c00", 80=>x"6e00", 81=>x"6b00", 82=>x"6c00", 83=>x"6700", 84=>x"6c00",
---- 85=>x"7300", 86=>x"7f00", 87=>x"8a00", 88=>x"6e00", 89=>x"6f00", 90=>x"6a00", 91=>x"6800",
---- 92=>x"6a00", 93=>x"6d00", 94=>x"8400", 95=>x"8800", 96=>x"6e00", 97=>x"6d00", 98=>x"6a00",
---- 99=>x"6a00", 100=>x"6f00", 101=>x"7200", 102=>x"7c00", 103=>x"8500", 104=>x"6e00", 105=>x"6d00",
---- 106=>x"6a00", 107=>x"6900", 108=>x"6e00", 109=>x"7500", 110=>x"7900", 111=>x"8500", 112=>x"7000",
---- 113=>x"6f00", 114=>x"6b00", 115=>x"6a00", 116=>x"6e00", 117=>x"7500", 118=>x"7d00", 119=>x"8400",
---- 120=>x"7000", 121=>x"7000", 122=>x"6e00", 123=>x"6c00", 124=>x"6d00", 125=>x"7600", 126=>x"7e00",
---- 127=>x"8600", 128=>x"9200", 129=>x"6e00", 130=>x"6c00", 131=>x"6b00", 132=>x"6c00", 133=>x"7400",
---- 134=>x"8000", 135=>x"8400", 136=>x"6f00", 137=>x"7200", 138=>x"6c00", 139=>x"6b00", 140=>x"7100",
---- 141=>x"7500", 142=>x"7900", 143=>x"8100", 144=>x"7200", 145=>x"7200", 146=>x"6e00", 147=>x"6b00",
---- 148=>x"6e00", 149=>x"7500", 150=>x"7900", 151=>x"8100", 152=>x"7400", 153=>x"6f00", 154=>x"6c00",
---- 155=>x"6900", 156=>x"6b00", 157=>x"7000", 158=>x"7a00", 159=>x"8200", 160=>x"7100", 161=>x"7300",
---- 162=>x"7000", 163=>x"6e00", 164=>x"6f00", 165=>x"7500", 166=>x"7c00", 167=>x"8100", 168=>x"8d00",
---- 169=>x"7300", 170=>x"6f00", 171=>x"6d00", 172=>x"6d00", 173=>x"7300", 174=>x"7900", 175=>x"7c00",
---- 176=>x"7400", 177=>x"7000", 178=>x"6d00", 179=>x"6a00", 180=>x"6e00", 181=>x"7000", 182=>x"7300",
---- 183=>x"7d00", 184=>x"7500", 185=>x"6f00", 186=>x"6e00", 187=>x"6900", 188=>x"6d00", 189=>x"7300",
---- 190=>x"7500", 191=>x"7e00", 192=>x"7200", 193=>x"7200", 194=>x"6e00", 195=>x"6c00", 196=>x"6c00",
---- 197=>x"6f00", 198=>x"7700", 199=>x"7c00", 200=>x"7000", 201=>x"9100", 202=>x"6d00", 203=>x"6b00",
---- 204=>x"6c00", 205=>x"6f00", 206=>x"7600", 207=>x"7c00", 208=>x"7100", 209=>x"6f00", 210=>x"6c00",
---- 211=>x"6900", 212=>x"6a00", 213=>x"6e00", 214=>x"7300", 215=>x"7e00", 216=>x"7000", 217=>x"7400",
---- 218=>x"6e00", 219=>x"6700", 220=>x"6c00", 221=>x"7000", 222=>x"7700", 223=>x"8000", 224=>x"7200",
---- 225=>x"6d00", 226=>x"6f00", 227=>x"6a00", 228=>x"6f00", 229=>x"7200", 230=>x"7700", 231=>x"7f00",
---- 232=>x"6d00", 233=>x"6b00", 234=>x"6900", 235=>x"6b00", 236=>x"6c00", 237=>x"7000", 238=>x"7500",
---- 239=>x"7d00", 240=>x"6c00", 241=>x"6b00", 242=>x"6700", 243=>x"6600", 244=>x"6c00", 245=>x"6f00",
---- 246=>x"7400", 247=>x"7c00", 248=>x"6c00", 249=>x"6900", 250=>x"6900", 251=>x"6300", 252=>x"6b00",
---- 253=>x"6f00", 254=>x"7400", 255=>x"8000", 256=>x"6a00", 257=>x"6a00", 258=>x"6900", 259=>x"6500",
---- 260=>x"6800", 261=>x"6d00", 262=>x"7200", 263=>x"7e00", 264=>x"9400", 265=>x"6a00", 266=>x"6500",
---- 267=>x"6500", 268=>x"6500", 269=>x"6e00", 270=>x"7400", 271=>x"8000", 272=>x"6b00", 273=>x"6a00",
---- 274=>x"6900", 275=>x"6500", 276=>x"6800", 277=>x"6d00", 278=>x"7400", 279=>x"7e00", 280=>x"6a00",
---- 281=>x"6c00", 282=>x"6900", 283=>x"6400", 284=>x"6600", 285=>x"6d00", 286=>x"7200", 287=>x"7d00",
---- 288=>x"6f00", 289=>x"6d00", 290=>x"9600", 291=>x"9800", 292=>x"6500", 293=>x"6a00", 294=>x"7300",
---- 295=>x"7e00", 296=>x"6b00", 297=>x"6a00", 298=>x"6600", 299=>x"6400", 300=>x"6400", 301=>x"9500",
---- 302=>x"7100", 303=>x"7c00", 304=>x"6a00", 305=>x"6900", 306=>x"6700", 307=>x"6300", 308=>x"6400",
---- 309=>x"6f00", 310=>x"7200", 311=>x"7f00", 312=>x"6800", 313=>x"9900", 314=>x"6700", 315=>x"6200",
---- 316=>x"6600", 317=>x"6a00", 318=>x"7000", 319=>x"7f00", 320=>x"6500", 321=>x"6600", 322=>x"6400",
---- 323=>x"6100", 324=>x"6500", 325=>x"6c00", 326=>x"7000", 327=>x"7e00", 328=>x"6500", 329=>x"6400",
---- 330=>x"6500", 331=>x"5e00", 332=>x"6000", 333=>x"6b00", 334=>x"6f00", 335=>x"7d00", 336=>x"6200",
---- 337=>x"6100", 338=>x"6200", 339=>x"6000", 340=>x"5f00", 341=>x"6b00", 342=>x"7000", 343=>x"7c00",
---- 344=>x"6700", 345=>x"6000", 346=>x"6000", 347=>x"5e00", 348=>x"6000", 349=>x"6800", 350=>x"6f00",
---- 351=>x"7b00", 352=>x"6000", 353=>x"5e00", 354=>x"6000", 355=>x"5e00", 356=>x"6000", 357=>x"9800",
---- 358=>x"7200", 359=>x"7a00", 360=>x"6000", 361=>x"a000", 362=>x"5f00", 363=>x"5e00", 364=>x"5f00",
---- 365=>x"6500", 366=>x"6e00", 367=>x"7b00", 368=>x"5800", 369=>x"5800", 370=>x"5b00", 371=>x"5a00",
---- 372=>x"5d00", 373=>x"6600", 374=>x"6f00", 375=>x"7c00", 376=>x"5400", 377=>x"5800", 378=>x"5a00",
---- 379=>x"5800", 380=>x"5e00", 381=>x"6500", 382=>x"7000", 383=>x"7d00", 384=>x"4f00", 385=>x"5400",
---- 386=>x"5700", 387=>x"5700", 388=>x"5900", 389=>x"6300", 390=>x"7000", 391=>x"7c00", 392=>x"4900",
---- 393=>x"4d00", 394=>x"5500", 395=>x"5400", 396=>x"5900", 397=>x"6100", 398=>x"6e00", 399=>x"7d00",
---- 400=>x"4500", 401=>x"4900", 402=>x"4f00", 403=>x"5100", 404=>x"5600", 405=>x"6200", 406=>x"6c00",
---- 407=>x"7900", 408=>x"4300", 409=>x"4200", 410=>x"4700", 411=>x"4d00", 412=>x"5300", 413=>x"5c00",
---- 414=>x"6c00", 415=>x"7d00", 416=>x"7500", 417=>x"3200", 418=>x"4000", 419=>x"4800", 420=>x"5200",
---- 421=>x"5d00", 422=>x"6b00", 423=>x"7b00", 424=>x"c200", 425=>x"4d00", 426=>x"3900", 427=>x"4500",
---- 428=>x"4e00", 429=>x"5900", 430=>x"6800", 431=>x"7900", 432=>x"dc00", 433=>x"8000", 434=>x"4d00",
---- 435=>x"4600", 436=>x"4700", 437=>x"5600", 438=>x"6400", 439=>x"7500", 440=>x"e300", 441=>x"cb00",
---- 442=>x"8900", 443=>x"3900", 444=>x"4700", 445=>x"4f00", 446=>x"6300", 447=>x"7700", 448=>x"e200",
---- 449=>x"e600", 450=>x"c100", 451=>x"4a00", 452=>x"3a00", 453=>x"4c00", 454=>x"6000", 455=>x"7600",
---- 456=>x"1e00", 457=>x"1d00", 458=>x"e200", 459=>x"7500", 460=>x"3100", 461=>x"4d00", 462=>x"5f00",
---- 463=>x"7200", 464=>x"e100", 465=>x"de00", 466=>x"e300", 467=>x"a400", 468=>x"3900", 469=>x"4700",
---- 470=>x"5a00", 471=>x"7200", 472=>x"da00", 473=>x"e100", 474=>x"e100", 475=>x"cc00", 476=>x"a500",
---- 477=>x"3d00", 478=>x"5700", 479=>x"6b00", 480=>x"d600", 481=>x"dd00", 482=>x"e100", 483=>x"df00",
---- 484=>x"9b00", 485=>x"4000", 486=>x"5100", 487=>x"6a00", 488=>x"d000", 489=>x"d900", 490=>x"e000",
---- 491=>x"e000", 492=>x"d100", 493=>x"7100", 494=>x"4600", 495=>x"6600", 496=>x"cd00", 497=>x"d300",
---- 498=>x"da00", 499=>x"de00", 500=>x"e000", 501=>x"b400", 502=>x"5400", 503=>x"5d00", 504=>x"cd00",
---- 505=>x"d000", 506=>x"d100", 507=>x"d600", 508=>x"da00", 509=>x"db00", 510=>x"8800", 511=>x"5400",
---- 512=>x"ce00", 513=>x"cf00", 514=>x"cf00", 515=>x"d300", 516=>x"d500", 517=>x"db00", 518=>x"c000",
---- 519=>x"7800", 520=>x"ce00", 521=>x"ce00", 522=>x"cf00", 523=>x"cf00", 524=>x"d200", 525=>x"d700",
---- 526=>x"d900", 527=>x"c400", 528=>x"ca00", 529=>x"cd00", 530=>x"cb00", 531=>x"cb00", 532=>x"ce00",
---- 533=>x"d400", 534=>x"d500", 535=>x"d800", 536=>x"c800", 537=>x"c600", 538=>x"c400", 539=>x"c700",
---- 540=>x"cb00", 541=>x"cd00", 542=>x"d200", 543=>x"d400", 544=>x"c800", 545=>x"c600", 546=>x"c500",
---- 547=>x"c200", 548=>x"c600", 549=>x"c800", 550=>x"cb00", 551=>x"cf00", 552=>x"c800", 553=>x"c900",
---- 554=>x"c600", 555=>x"c400", 556=>x"c100", 557=>x"c400", 558=>x"c600", 559=>x"c500", 560=>x"c000",
---- 561=>x"c400", 562=>x"c400", 563=>x"c500", 564=>x"c000", 565=>x"bc00", 566=>x"c300", 567=>x"bf00",
---- 568=>x"bd00", 569=>x"bc00", 570=>x"c100", 571=>x"c200", 572=>x"c000", 573=>x"b800", 574=>x"bc00",
---- 575=>x"bc00", 576=>x"be00", 577=>x"bf00", 578=>x"bb00", 579=>x"be00", 580=>x"bb00", 581=>x"b800",
---- 582=>x"b800", 583=>x"bf00", 584=>x"bb00", 585=>x"bc00", 586=>x"b700", 587=>x"4600", 588=>x"bb00",
---- 589=>x"b600", 590=>x"b200", 591=>x"ba00", 592=>x"ba00", 593=>x"b300", 594=>x"b900", 595=>x"4900",
---- 596=>x"b900", 597=>x"b300", 598=>x"ac00", 599=>x"aa00", 600=>x"b900", 601=>x"b600", 602=>x"b000",
---- 603=>x"b300", 604=>x"b000", 605=>x"ae00", 606=>x"a200", 607=>x"a200", 608=>x"b900", 609=>x"b800",
---- 610=>x"aa00", 611=>x"ae00", 612=>x"a200", 613=>x"9f00", 614=>x"a000", 615=>x"ba00", 616=>x"b500",
---- 617=>x"b300", 618=>x"a700", 619=>x"a000", 620=>x"9b00", 621=>x"b000", 622=>x"c900", 623=>x"cc00",
---- 624=>x"ab00", 625=>x"a800", 626=>x"9c00", 627=>x"a400", 628=>x"c200", 629=>x"d000", 630=>x"c100",
---- 631=>x"b400", 632=>x"9800", 633=>x"a600", 634=>x"b700", 635=>x"c700", 636=>x"c200", 637=>x"b700",
---- 638=>x"b600", 639=>x"ba00", 640=>x"aa00", 641=>x"c600", 642=>x"c500", 643=>x"b500", 644=>x"b100",
---- 645=>x"b300", 646=>x"bc00", 647=>x"c500", 648=>x"c800", 649=>x"b700", 650=>x"a900", 651=>x"b200",
---- 652=>x"bc00", 653=>x"c100", 654=>x"c400", 655=>x"cd00", 656=>x"af00", 657=>x"af00", 658=>x"b500",
---- 659=>x"bf00", 660=>x"c400", 661=>x"cc00", 662=>x"cb00", 663=>x"cb00", 664=>x"b200", 665=>x"bc00",
---- 666=>x"c200", 667=>x"c600", 668=>x"c700", 669=>x"c700", 670=>x"c400", 671=>x"c200", 672=>x"ba00",
---- 673=>x"ca00", 674=>x"cd00", 675=>x"c800", 676=>x"c000", 677=>x"bd00", 678=>x"b900", 679=>x"b700",
---- 680=>x"c100", 681=>x"cc00", 682=>x"c800", 683=>x"bf00", 684=>x"bb00", 685=>x"bb00", 686=>x"bb00",
---- 687=>x"bc00", 688=>x"c500", 689=>x"c600", 690=>x"c200", 691=>x"bc00", 692=>x"bd00", 693=>x"c000",
---- 694=>x"c100", 695=>x"c000", 696=>x"c100", 697=>x"c500", 698=>x"c200", 699=>x"c100", 700=>x"bf00",
---- 701=>x"c000", 702=>x"c000", 703=>x"c000", 704=>x"3f00", 705=>x"c300", 706=>x"c300", 707=>x"c300",
---- 708=>x"c300", 709=>x"c300", 710=>x"be00", 711=>x"bf00", 712=>x"c200", 713=>x"c500", 714=>x"c500",
---- 715=>x"c100", 716=>x"c000", 717=>x"c200", 718=>x"bf00", 719=>x"c000", 720=>x"c300", 721=>x"c500",
---- 722=>x"c300", 723=>x"c100", 724=>x"be00", 725=>x"be00", 726=>x"c100", 727=>x"c300", 728=>x"c200",
---- 729=>x"c100", 730=>x"c300", 731=>x"c300", 732=>x"be00", 733=>x"c000", 734=>x"c100", 735=>x"c400",
---- 736=>x"c300", 737=>x"c500", 738=>x"c200", 739=>x"c200", 740=>x"c200", 741=>x"c000", 742=>x"c200",
---- 743=>x"c200", 744=>x"4000", 745=>x"c100", 746=>x"c300", 747=>x"c300", 748=>x"c000", 749=>x"bf00",
---- 750=>x"c000", 751=>x"c000", 752=>x"be00", 753=>x"3e00", 754=>x"be00", 755=>x"be00", 756=>x"bd00",
---- 757=>x"c100", 758=>x"c100", 759=>x"c200", 760=>x"be00", 761=>x"bd00", 762=>x"bf00", 763=>x"be00",
---- 764=>x"bf00", 765=>x"c100", 766=>x"c000", 767=>x"c100", 768=>x"bb00", 769=>x"be00", 770=>x"c000",
---- 771=>x"be00", 772=>x"bf00", 773=>x"be00", 774=>x"c200", 775=>x"c200", 776=>x"4400", 777=>x"be00",
---- 778=>x"bf00", 779=>x"be00", 780=>x"bf00", 781=>x"c000", 782=>x"c200", 783=>x"c300", 784=>x"bd00",
---- 785=>x"bf00", 786=>x"c100", 787=>x"bf00", 788=>x"bd00", 789=>x"c200", 790=>x"c300", 791=>x"c300",
---- 792=>x"bd00", 793=>x"bd00", 794=>x"be00", 795=>x"bd00", 796=>x"c200", 797=>x"c200", 798=>x"c400",
---- 799=>x"c800", 800=>x"bd00", 801=>x"c100", 802=>x"c000", 803=>x"bd00", 804=>x"c100", 805=>x"c300",
---- 806=>x"4100", 807=>x"a100", 808=>x"c000", 809=>x"c000", 810=>x"c100", 811=>x"bf00", 812=>x"bc00",
---- 813=>x"b900", 814=>x"ac00", 815=>x"7600", 816=>x"bc00", 817=>x"bc00", 818=>x"b900", 819=>x"b600",
---- 820=>x"b900", 821=>x"c000", 822=>x"b800", 823=>x"a200", 824=>x"b700", 825=>x"b600", 826=>x"b300",
---- 827=>x"b900", 828=>x"c000", 829=>x"c200", 830=>x"bf00", 831=>x"ae00", 832=>x"ba00", 833=>x"ba00",
---- 834=>x"bc00", 835=>x"c100", 836=>x"c600", 837=>x"c400", 838=>x"bf00", 839=>x"b400", 840=>x"c000",
---- 841=>x"c100", 842=>x"c200", 843=>x"c300", 844=>x"c400", 845=>x"ca00", 846=>x"c500", 847=>x"c000",
---- 848=>x"c100", 849=>x"3f00", 850=>x"c300", 851=>x"c500", 852=>x"c300", 853=>x"c600", 854=>x"c600",
---- 855=>x"c400", 856=>x"c300", 857=>x"3b00", 858=>x"c500", 859=>x"c600", 860=>x"c500", 861=>x"c500",
---- 862=>x"c800", 863=>x"c500", 864=>x"c500", 865=>x"c400", 866=>x"c600", 867=>x"c400", 868=>x"c600",
---- 869=>x"c600", 870=>x"c500", 871=>x"c500", 872=>x"c700", 873=>x"c400", 874=>x"c400", 875=>x"c700",
---- 876=>x"ca00", 877=>x"c800", 878=>x"c900", 879=>x"c400", 880=>x"c800", 881=>x"c700", 882=>x"c900",
---- 883=>x"c900", 884=>x"cb00", 885=>x"cc00", 886=>x"cc00", 887=>x"ca00", 888=>x"c800", 889=>x"3600",
---- 890=>x"cc00", 891=>x"cc00", 892=>x"d100", 893=>x"d200", 894=>x"cf00", 895=>x"d100", 896=>x"c700",
---- 897=>x"c800", 898=>x"cb00", 899=>x"ce00", 900=>x"d100", 901=>x"d300", 902=>x"d100", 903=>x"d200",
---- 904=>x"c900", 905=>x"c900", 906=>x"ce00", 907=>x"d000", 908=>x"cf00", 909=>x"d200", 910=>x"d100",
---- 911=>x"d300", 912=>x"ca00", 913=>x"cb00", 914=>x"d000", 915=>x"d200", 916=>x"2c00", 917=>x"d200",
---- 918=>x"d400", 919=>x"d400", 920=>x"cb00", 921=>x"cb00", 922=>x"ce00", 923=>x"d100", 924=>x"d200",
---- 925=>x"d200", 926=>x"d300", 927=>x"d400", 928=>x"cc00", 929=>x"cc00", 930=>x"d000", 931=>x"cf00",
---- 932=>x"d100", 933=>x"d300", 934=>x"d500", 935=>x"d500", 936=>x"cb00", 937=>x"cd00", 938=>x"ce00",
---- 939=>x"d000", 940=>x"d100", 941=>x"d200", 942=>x"d500", 943=>x"d600", 944=>x"cb00", 945=>x"cc00",
---- 946=>x"cc00", 947=>x"cf00", 948=>x"d200", 949=>x"d100", 950=>x"d400", 951=>x"d500", 952=>x"c900",
---- 953=>x"ca00", 954=>x"cd00", 955=>x"cc00", 956=>x"cf00", 957=>x"d100", 958=>x"d200", 959=>x"d300",
---- 960=>x"c800", 961=>x"c900", 962=>x"ca00", 963=>x"cb00", 964=>x"cd00", 965=>x"d100", 966=>x"d200",
---- 967=>x"d300", 968=>x"c600", 969=>x"c600", 970=>x"c900", 971=>x"cc00", 972=>x"ca00", 973=>x"ce00",
---- 974=>x"d100", 975=>x"d400", 976=>x"c300", 977=>x"c500", 978=>x"c800", 979=>x"c900", 980=>x"c900",
---- 981=>x"cb00", 982=>x"ce00", 983=>x"d200", 984=>x"c000", 985=>x"c100", 986=>x"c400", 987=>x"c800",
---- 988=>x"c800", 989=>x"ca00", 990=>x"ce00", 991=>x"ce00", 992=>x"bd00", 993=>x"c000", 994=>x"c300",
---- 995=>x"c700", 996=>x"c900", 997=>x"c800", 998=>x"cd00", 999=>x"ca00", 1000=>x"c300", 1001=>x"c100",
---- 1002=>x"be00", 1003=>x"c200", 1004=>x"c200", 1005=>x"b900", 1006=>x"a900", 1007=>x"8d00", 1008=>x"c100",
---- 1009=>x"bf00", 1010=>x"b900", 1011=>x"bb00", 1012=>x"aa00", 1013=>x"8700", 1014=>x"6200", 1015=>x"5200",
---- 1016=>x"be00", 1017=>x"ba00", 1018=>x"b000", 1019=>x"a700", 1020=>x"8400", 1021=>x"9200", 1022=>x"6800",
---- 1023=>x"7000", 1024=>x"bf00", 1025=>x"bd00", 1026=>x"aa00", 1027=>x"9300", 1028=>x"8400", 1029=>x"8000",
---- 1030=>x"6f00", 1031=>x"5500", 1032=>x"bf00", 1033=>x"b800", 1034=>x"9b00", 1035=>x"7500", 1036=>x"5900",
---- 1037=>x"4600", 1038=>x"3600", 1039=>x"3100", 1040=>x"be00", 1041=>x"9900", 1042=>x"6000", 1043=>x"4000",
---- 1044=>x"3300", 1045=>x"3200", 1046=>x"3200", 1047=>x"3900", 1048=>x"9a00", 1049=>x"4500", 1050=>x"3200",
---- 1051=>x"3000", 1052=>x"3500", 1053=>x"3a00", 1054=>x"3e00", 1055=>x"5600", 1056=>x"5000", 1057=>x"2c00",
---- 1058=>x"3100", 1059=>x"2c00", 1060=>x"2e00", 1061=>x"3e00", 1062=>x"7d00", 1063=>x"6e00", 1064=>x"4000",
---- 1065=>x"3600", 1066=>x"4400", 1067=>x"3400", 1068=>x"2b00", 1069=>x"4100", 1070=>x"6100", 1071=>x"6100",
---- 1072=>x"6200", 1073=>x"4500", 1074=>x"5300", 1075=>x"5800", 1076=>x"4600", 1077=>x"5f00", 1078=>x"3f00",
---- 1079=>x"6000", 1080=>x"8400", 1081=>x"7500", 1082=>x"4900", 1083=>x"5d00", 1084=>x"5f00", 1085=>x"4d00",
---- 1086=>x"4f00", 1087=>x"9a00", 1088=>x"7800", 1089=>x"9100", 1090=>x"7400", 1091=>x"5900", 1092=>x"5900",
---- 1093=>x"6500", 1094=>x"9a00", 1095=>x"ba00", 1096=>x"6100", 1097=>x"7700", 1098=>x"8c00", 1099=>x"8c00",
---- 1100=>x"7100", 1101=>x"a100", 1102=>x"b000", 1103=>x"5300", 1104=>x"9500", 1105=>x"8600", 1106=>x"9100",
---- 1107=>x"8f00", 1108=>x"8600", 1109=>x"9000", 1110=>x"9400", 1111=>x"8100", 1112=>x"9800", 1113=>x"9000",
---- 1114=>x"8f00", 1115=>x"7d00", 1116=>x"6d00", 1117=>x"8f00", 1118=>x"6f00", 1119=>x"5b00", 1120=>x"9500",
---- 1121=>x"8d00", 1122=>x"8500", 1123=>x"8000", 1124=>x"7e00", 1125=>x"7d00", 1126=>x"7d00", 1127=>x"7500",
---- 1128=>x"a300", 1129=>x"9d00", 1130=>x"9100", 1131=>x"8c00", 1132=>x"8a00", 1133=>x"8400", 1134=>x"7e00",
---- 1135=>x"7c00", 1136=>x"aa00", 1137=>x"a000", 1138=>x"9c00", 1139=>x"9700", 1140=>x"9200", 1141=>x"8500",
---- 1142=>x"8000", 1143=>x"8000", 1144=>x"b000", 1145=>x"a100", 1146=>x"9e00", 1147=>x"9a00", 1148=>x"9800",
---- 1149=>x"8c00", 1150=>x"7900", 1151=>x"8300", 1152=>x"b500", 1153=>x"5500", 1154=>x"9f00", 1155=>x"9900",
---- 1156=>x"9500", 1157=>x"8e00", 1158=>x"8900", 1159=>x"8600", 1160=>x"af00", 1161=>x"ad00", 1162=>x"a400",
---- 1163=>x"9700", 1164=>x"9200", 1165=>x"8d00", 1166=>x"8800", 1167=>x"8800", 1168=>x"aa00", 1169=>x"a800",
---- 1170=>x"a500", 1171=>x"9e00", 1172=>x"9700", 1173=>x"8d00", 1174=>x"8900", 1175=>x"8500", 1176=>x"aa00",
---- 1177=>x"a400", 1178=>x"a200", 1179=>x"a000", 1180=>x"9700", 1181=>x"8f00", 1182=>x"8800", 1183=>x"8600",
---- 1184=>x"a900", 1185=>x"a300", 1186=>x"a100", 1187=>x"9f00", 1188=>x"9b00", 1189=>x"9100", 1190=>x"8d00",
---- 1191=>x"8700", 1192=>x"a900", 1193=>x"a400", 1194=>x"a400", 1195=>x"9e00", 1196=>x"9800", 1197=>x"9400",
---- 1198=>x"8f00", 1199=>x"8900", 1200=>x"a700", 1201=>x"a800", 1202=>x"a300", 1203=>x"9e00", 1204=>x"9900",
---- 1205=>x"9200", 1206=>x"9000", 1207=>x"8a00", 1208=>x"a500", 1209=>x"a400", 1210=>x"9f00", 1211=>x"9a00",
---- 1212=>x"9500", 1213=>x"9500", 1214=>x"9200", 1215=>x"8a00", 1216=>x"a100", 1217=>x"a000", 1218=>x"a000",
---- 1219=>x"9b00", 1220=>x"9400", 1221=>x"9600", 1222=>x"8f00", 1223=>x"8b00", 1224=>x"a400", 1225=>x"a400",
---- 1226=>x"9e00", 1227=>x"9b00", 1228=>x"9400", 1229=>x"9300", 1230=>x"8c00", 1231=>x"8800", 1232=>x"a500",
---- 1233=>x"9f00", 1234=>x"9c00", 1235=>x"9800", 1236=>x"9500", 1237=>x"9100", 1238=>x"8e00", 1239=>x"8a00",
---- 1240=>x"ab00", 1241=>x"9b00", 1242=>x"9b00", 1243=>x"9800", 1244=>x"9400", 1245=>x"9000", 1246=>x"8e00",
---- 1247=>x"8900", 1248=>x"b300", 1249=>x"9900", 1250=>x"9d00", 1251=>x"9600", 1252=>x"9600", 1253=>x"9400",
---- 1254=>x"7400", 1255=>x"8900", 1256=>x"ba00", 1257=>x"9300", 1258=>x"6800", 1259=>x"9700", 1260=>x"9800",
---- 1261=>x"9300", 1262=>x"8a00", 1263=>x"8700", 1264=>x"bb00", 1265=>x"8e00", 1266=>x"9300", 1267=>x"9500",
---- 1268=>x"9600", 1269=>x"9000", 1270=>x"8b00", 1271=>x"8400", 1272=>x"b700", 1273=>x"8d00", 1274=>x"9700",
---- 1275=>x"6c00", 1276=>x"9100", 1277=>x"8b00", 1278=>x"8800", 1279=>x"8200", 1280=>x"a800", 1281=>x"8f00",
---- 1282=>x"9400", 1283=>x"9400", 1284=>x"9100", 1285=>x"8e00", 1286=>x"8a00", 1287=>x"8300", 1288=>x"9900",
---- 1289=>x"9400", 1290=>x"9300", 1291=>x"9600", 1292=>x"9000", 1293=>x"8d00", 1294=>x"8600", 1295=>x"7f00",
---- 1296=>x"a100", 1297=>x"9700", 1298=>x"9200", 1299=>x"9200", 1300=>x"8d00", 1301=>x"8c00", 1302=>x"8700",
---- 1303=>x"8100", 1304=>x"a200", 1305=>x"9900", 1306=>x"9400", 1307=>x"8e00", 1308=>x"8c00", 1309=>x"8a00",
---- 1310=>x"8300", 1311=>x"8400", 1312=>x"9e00", 1313=>x"9900", 1314=>x"9500", 1315=>x"8f00", 1316=>x"8a00",
---- 1317=>x"8500", 1318=>x"8400", 1319=>x"8100", 1320=>x"9b00", 1321=>x"9600", 1322=>x"9500", 1323=>x"8f00",
---- 1324=>x"8b00", 1325=>x"8500", 1326=>x"8200", 1327=>x"7800", 1328=>x"9a00", 1329=>x"9700", 1330=>x"9100",
---- 1331=>x"8d00", 1332=>x"7800", 1333=>x"8300", 1334=>x"8300", 1335=>x"6b00", 1336=>x"9900", 1337=>x"9100",
---- 1338=>x"9200", 1339=>x"8e00", 1340=>x"8600", 1341=>x"8600", 1342=>x"7f00", 1343=>x"4b00", 1344=>x"9700",
---- 1345=>x"9000", 1346=>x"9200", 1347=>x"8c00", 1348=>x"8700", 1349=>x"8a00", 1350=>x"6c00", 1351=>x"3100",
---- 1352=>x"9400", 1353=>x"9000", 1354=>x"9000", 1355=>x"8a00", 1356=>x"8800", 1357=>x"8400", 1358=>x"4d00",
---- 1359=>x"2a00", 1360=>x"8d00", 1361=>x"9200", 1362=>x"8d00", 1363=>x"8800", 1364=>x"8a00", 1365=>x"7300",
---- 1366=>x"3600", 1367=>x"2e00", 1368=>x"8d00", 1369=>x"8e00", 1370=>x"8b00", 1371=>x"8a00", 1372=>x"8800",
---- 1373=>x"5500", 1374=>x"2900", 1375=>x"2e00", 1376=>x"8300", 1377=>x"8600", 1378=>x"8a00", 1379=>x"8d00",
---- 1380=>x"7a00", 1381=>x"3a00", 1382=>x"2a00", 1383=>x"2d00", 1384=>x"7700", 1385=>x"7900", 1386=>x"8c00",
---- 1387=>x"8c00", 1388=>x"5700", 1389=>x"2b00", 1390=>x"2f00", 1391=>x"2f00", 1392=>x"7800", 1393=>x"8e00",
---- 1394=>x"9000", 1395=>x"7e00", 1396=>x"3900", 1397=>x"2e00", 1398=>x"2e00", 1399=>x"2f00", 1400=>x"8700",
---- 1401=>x"9000", 1402=>x"9300", 1403=>x"5d00", 1404=>x"2a00", 1405=>x"2f00", 1406=>x"2b00", 1407=>x"cf00",
---- 1408=>x"9100", 1409=>x"9200", 1410=>x"8100", 1411=>x"3700", 1412=>x"2a00", 1413=>x"2d00", 1414=>x"2e00",
---- 1415=>x"3300", 1416=>x"9000", 1417=>x"8c00", 1418=>x"ad00", 1419=>x"2800", 1420=>x"2f00", 1421=>x"2f00",
---- 1422=>x"2f00", 1423=>x"3700", 1424=>x"8c00", 1425=>x"7000", 1426=>x"3100", 1427=>x"2c00", 1428=>x"2a00",
---- 1429=>x"2e00", 1430=>x"3300", 1431=>x"3500", 1432=>x"8800", 1433=>x"4400", 1434=>x"2800", 1435=>x"2d00",
---- 1436=>x"2b00", 1437=>x"2d00", 1438=>x"3500", 1439=>x"3200", 1440=>x"6900", 1441=>x"2e00", 1442=>x"2e00",
---- 1443=>x"2f00", 1444=>x"2d00", 1445=>x"2f00", 1446=>x"3800", 1447=>x"3000", 1448=>x"4d00", 1449=>x"2900",
---- 1450=>x"2f00", 1451=>x"3000", 1452=>x"2f00", 1453=>x"3300", 1454=>x"3700", 1455=>x"3000", 1456=>x"4100",
---- 1457=>x"2a00", 1458=>x"2c00", 1459=>x"2900", 1460=>x"2a00", 1461=>x"2f00", 1462=>x"2d00", 1463=>x"3000",
---- 1464=>x"4100", 1465=>x"2900", 1466=>x"2e00", 1467=>x"2b00", 1468=>x"2b00", 1469=>x"2f00", 1470=>x"3500",
---- 1471=>x"3500", 1472=>x"3e00", 1473=>x"2e00", 1474=>x"2c00", 1475=>x"2d00", 1476=>x"2d00", 1477=>x"3400",
---- 1478=>x"3a00", 1479=>x"3400", 1480=>x"3800", 1481=>x"2a00", 1482=>x"2b00", 1483=>x"2e00", 1484=>x"3100",
---- 1485=>x"3200", 1486=>x"3300", 1487=>x"3c00", 1488=>x"3000", 1489=>x"2b00", 1490=>x"2e00", 1491=>x"3100",
---- 1492=>x"2f00", 1493=>x"3300", 1494=>x"3a00", 1495=>x"3f00", 1496=>x"2d00", 1497=>x"2c00", 1498=>x"3000",
---- 1499=>x"3000", 1500=>x"3200", 1501=>x"3900", 1502=>x"3f00", 1503=>x"3900", 1504=>x"2b00", 1505=>x"3100",
---- 1506=>x"3400", 1507=>x"2f00", 1508=>x"3200", 1509=>x"3800", 1510=>x"4000", 1511=>x"3800", 1512=>x"3000",
---- 1513=>x"3500", 1514=>x"3500", 1515=>x"3200", 1516=>x"3500", 1517=>x"3600", 1518=>x"c200", 1519=>x"4200",
---- 1520=>x"3500", 1521=>x"3900", 1522=>x"3800", 1523=>x"3600", 1524=>x"3500", 1525=>x"3700", 1526=>x"3c00",
---- 1527=>x"4600", 1528=>x"3800", 1529=>x"3b00", 1530=>x"3a00", 1531=>x"3900", 1532=>x"3800", 1533=>x"3700",
---- 1534=>x"3c00", 1535=>x"4a00", 1536=>x"3800", 1537=>x"3500", 1538=>x"3700", 1539=>x"3900", 1540=>x"3900",
---- 1541=>x"3600", 1542=>x"4000", 1543=>x"4300", 1544=>x"3900", 1545=>x"3800", 1546=>x"3700", 1547=>x"3a00",
---- 1548=>x"3900", 1549=>x"3400", 1550=>x"4000", 1551=>x"4300", 1552=>x"3f00", 1553=>x"3c00", 1554=>x"3900",
---- 1555=>x"3700", 1556=>x"3a00", 1557=>x"3400", 1558=>x"3d00", 1559=>x"4200", 1560=>x"3300", 1561=>x"3200",
---- 1562=>x"3600", 1563=>x"3800", 1564=>x"3500", 1565=>x"3300", 1566=>x"3600", 1567=>x"3a00", 1568=>x"6a00",
---- 1569=>x"4400", 1570=>x"3500", 1571=>x"3700", 1572=>x"3500", 1573=>x"3300", 1574=>x"3500", 1575=>x"3700",
---- 1576=>x"c900", 1577=>x"a700", 1578=>x"7700", 1579=>x"4b00", 1580=>x"3700", 1581=>x"3400", 1582=>x"3600",
---- 1583=>x"3a00", 1584=>x"cb00", 1585=>x"cf00", 1586=>x"c900", 1587=>x"ae00", 1588=>x"7d00", 1589=>x"4600",
---- 1590=>x"2f00", 1591=>x"2c00", 1592=>x"ca00", 1593=>x"c800", 1594=>x"cb00", 1595=>x"d300", 1596=>x"cf00",
---- 1597=>x"b000", 1598=>x"7800", 1599=>x"3e00", 1600=>x"ca00", 1601=>x"cb00", 1602=>x"3500", 1603=>x"cb00",
---- 1604=>x"cf00", 1605=>x"d500", 1606=>x"d000", 1607=>x"a600", 1608=>x"c800", 1609=>x"cb00", 1610=>x"cb00",
---- 1611=>x"cc00", 1612=>x"cc00", 1613=>x"ce00", 1614=>x"d300", 1615=>x"d800", 1616=>x"c600", 1617=>x"c700",
---- 1618=>x"ca00", 1619=>x"cc00", 1620=>x"cc00", 1621=>x"ce00", 1622=>x"cf00", 1623=>x"d100", 1624=>x"c300",
---- 1625=>x"c700", 1626=>x"c900", 1627=>x"cc00", 1628=>x"cc00", 1629=>x"cd00", 1630=>x"d000", 1631=>x"d000",
---- 1632=>x"c200", 1633=>x"c500", 1634=>x"c600", 1635=>x"c900", 1636=>x"cb00", 1637=>x"cd00", 1638=>x"cf00",
---- 1639=>x"d100", 1640=>x"c200", 1641=>x"c400", 1642=>x"3a00", 1643=>x"c700", 1644=>x"ca00", 1645=>x"3200",
---- 1646=>x"cf00", 1647=>x"cf00", 1648=>x"c000", 1649=>x"c100", 1650=>x"c100", 1651=>x"c700", 1652=>x"c900",
---- 1653=>x"ca00", 1654=>x"ce00", 1655=>x"d000", 1656=>x"bc00", 1657=>x"c000", 1658=>x"c400", 1659=>x"c700",
---- 1660=>x"c900", 1661=>x"ca00", 1662=>x"cb00", 1663=>x"cf00", 1664=>x"b900", 1665=>x"c000", 1666=>x"c200",
---- 1667=>x"c400", 1668=>x"c800", 1669=>x"c900", 1670=>x"cd00", 1671=>x"cf00", 1672=>x"ba00", 1673=>x"bf00",
---- 1674=>x"bf00", 1675=>x"c400", 1676=>x"c400", 1677=>x"c400", 1678=>x"cc00", 1679=>x"3200", 1680=>x"b900",
---- 1681=>x"be00", 1682=>x"bf00", 1683=>x"c400", 1684=>x"c500", 1685=>x"c700", 1686=>x"ca00", 1687=>x"cb00",
---- 1688=>x"b700", 1689=>x"c000", 1690=>x"c000", 1691=>x"c000", 1692=>x"c400", 1693=>x"c600", 1694=>x"ca00",
---- 1695=>x"cc00", 1696=>x"b800", 1697=>x"ba00", 1698=>x"bd00", 1699=>x"c000", 1700=>x"c500", 1701=>x"c500",
---- 1702=>x"c900", 1703=>x"cc00", 1704=>x"b900", 1705=>x"bb00", 1706=>x"bd00", 1707=>x"be00", 1708=>x"c400",
---- 1709=>x"c600", 1710=>x"c800", 1711=>x"cc00", 1712=>x"ba00", 1713=>x"ba00", 1714=>x"bb00", 1715=>x"bb00",
---- 1716=>x"c200", 1717=>x"c600", 1718=>x"ca00", 1719=>x"cc00", 1720=>x"b700", 1721=>x"bb00", 1722=>x"bc00",
---- 1723=>x"bd00", 1724=>x"c100", 1725=>x"c400", 1726=>x"c800", 1727=>x"cc00", 1728=>x"b400", 1729=>x"bb00",
---- 1730=>x"bc00", 1731=>x"bd00", 1732=>x"c300", 1733=>x"c400", 1734=>x"c700", 1735=>x"ca00", 1736=>x"b300",
---- 1737=>x"ba00", 1738=>x"bb00", 1739=>x"bc00", 1740=>x"c200", 1741=>x"c300", 1742=>x"c600", 1743=>x"cc00",
---- 1744=>x"b500", 1745=>x"ba00", 1746=>x"bc00", 1747=>x"bc00", 1748=>x"bf00", 1749=>x"c200", 1750=>x"c400",
---- 1751=>x"ca00", 1752=>x"b500", 1753=>x"b600", 1754=>x"ba00", 1755=>x"be00", 1756=>x"c100", 1757=>x"c300",
---- 1758=>x"c500", 1759=>x"c800", 1760=>x"b000", 1761=>x"4a00", 1762=>x"ba00", 1763=>x"bf00", 1764=>x"c000",
---- 1765=>x"c100", 1766=>x"c600", 1767=>x"c700", 1768=>x"b000", 1769=>x"b700", 1770=>x"ba00", 1771=>x"bd00",
---- 1772=>x"c000", 1773=>x"c000", 1774=>x"c500", 1775=>x"c800", 1776=>x"b200", 1777=>x"b600", 1778=>x"b900",
---- 1779=>x"bc00", 1780=>x"bd00", 1781=>x"3f00", 1782=>x"c400", 1783=>x"c700", 1784=>x"b000", 1785=>x"b200",
---- 1786=>x"b600", 1787=>x"b800", 1788=>x"bd00", 1789=>x"c000", 1790=>x"c300", 1791=>x"c500", 1792=>x"5000",
---- 1793=>x"af00", 1794=>x"b400", 1795=>x"b800", 1796=>x"bf00", 1797=>x"c000", 1798=>x"c000", 1799=>x"c500",
---- 1800=>x"ab00", 1801=>x"ae00", 1802=>x"b500", 1803=>x"b800", 1804=>x"ba00", 1805=>x"bf00", 1806=>x"c100",
---- 1807=>x"c500", 1808=>x"a900", 1809=>x"af00", 1810=>x"b400", 1811=>x"b700", 1812=>x"b900", 1813=>x"be00",
---- 1814=>x"c300", 1815=>x"c200", 1816=>x"aa00", 1817=>x"aa00", 1818=>x"af00", 1819=>x"b300", 1820=>x"ba00",
---- 1821=>x"ba00", 1822=>x"c000", 1823=>x"c100", 1824=>x"aa00", 1825=>x"ae00", 1826=>x"ad00", 1827=>x"b300",
---- 1828=>x"b700", 1829=>x"b900", 1830=>x"bf00", 1831=>x"c000", 1832=>x"a700", 1833=>x"ae00", 1834=>x"af00",
---- 1835=>x"b300", 1836=>x"b500", 1837=>x"b700", 1838=>x"bb00", 1839=>x"c000", 1840=>x"a800", 1841=>x"ab00",
---- 1842=>x"ab00", 1843=>x"b000", 1844=>x"b300", 1845=>x"b800", 1846=>x"bc00", 1847=>x"be00", 1848=>x"a600",
---- 1849=>x"a900", 1850=>x"a900", 1851=>x"ab00", 1852=>x"b100", 1853=>x"b700", 1854=>x"bb00", 1855=>x"bd00",
---- 1856=>x"a600", 1857=>x"aa00", 1858=>x"a800", 1859=>x"ac00", 1860=>x"ac00", 1861=>x"b200", 1862=>x"b900",
---- 1863=>x"bd00", 1864=>x"a700", 1865=>x"a900", 1866=>x"aa00", 1867=>x"ab00", 1868=>x"ad00", 1869=>x"b100",
---- 1870=>x"ba00", 1871=>x"b900", 1872=>x"a500", 1873=>x"a800", 1874=>x"a900", 1875=>x"a900", 1876=>x"a900",
---- 1877=>x"b100", 1878=>x"b600", 1879=>x"b800", 1880=>x"a200", 1881=>x"a400", 1882=>x"a700", 1883=>x"a800",
---- 1884=>x"ad00", 1885=>x"b100", 1886=>x"b300", 1887=>x"b900", 1888=>x"a000", 1889=>x"a300", 1890=>x"a600",
---- 1891=>x"a700", 1892=>x"ac00", 1893=>x"b200", 1894=>x"b000", 1895=>x"b600", 1896=>x"9e00", 1897=>x"a100",
---- 1898=>x"a500", 1899=>x"a600", 1900=>x"ac00", 1901=>x"b300", 1902=>x"af00", 1903=>x"b500", 1904=>x"9c00",
---- 1905=>x"9f00", 1906=>x"a400", 1907=>x"a600", 1908=>x"ab00", 1909=>x"ae00", 1910=>x"ae00", 1911=>x"b400",
---- 1912=>x"9b00", 1913=>x"a100", 1914=>x"9f00", 1915=>x"a700", 1916=>x"ab00", 1917=>x"a800", 1918=>x"ab00",
---- 1919=>x"b200", 1920=>x"6200", 1921=>x"a100", 1922=>x"a000", 1923=>x"a400", 1924=>x"a400", 1925=>x"a700",
---- 1926=>x"ab00", 1927=>x"ad00", 1928=>x"9c00", 1929=>x"9f00", 1930=>x"a200", 1931=>x"a600", 1932=>x"a200",
---- 1933=>x"a400", 1934=>x"ac00", 1935=>x"b100", 1936=>x"9900", 1937=>x"9e00", 1938=>x"a200", 1939=>x"a200",
---- 1940=>x"a300", 1941=>x"a600", 1942=>x"a900", 1943=>x"aa00", 1944=>x"9a00", 1945=>x"9e00", 1946=>x"a100",
---- 1947=>x"a100", 1948=>x"a200", 1949=>x"a800", 1950=>x"a800", 1951=>x"a700", 1952=>x"9a00", 1953=>x"9b00",
---- 1954=>x"6100", 1955=>x"9f00", 1956=>x"a100", 1957=>x"a800", 1958=>x"a800", 1959=>x"aa00", 1960=>x"9800",
---- 1961=>x"9b00", 1962=>x"9d00", 1963=>x"9f00", 1964=>x"a100", 1965=>x"a400", 1966=>x"a800", 1967=>x"aa00",
---- 1968=>x"9900", 1969=>x"9d00", 1970=>x"9f00", 1971=>x"9f00", 1972=>x"a000", 1973=>x"a300", 1974=>x"a600",
---- 1975=>x"a900", 1976=>x"9700", 1977=>x"9a00", 1978=>x"9f00", 1979=>x"9e00", 1980=>x"9d00", 1981=>x"a400",
---- 1982=>x"a500", 1983=>x"a600", 1984=>x"9400", 1985=>x"9a00", 1986=>x"9b00", 1987=>x"9b00", 1988=>x"9d00",
---- 1989=>x"a200", 1990=>x"a400", 1991=>x"aa00", 1992=>x"9600", 1993=>x"9900", 1994=>x"9b00", 1995=>x"9a00",
---- 1996=>x"9d00", 1997=>x"a000", 1998=>x"a400", 1999=>x"a600", 2000=>x"9600", 2001=>x"9500", 2002=>x"9900",
---- 2003=>x"9b00", 2004=>x"9d00", 2005=>x"a200", 2006=>x"a300", 2007=>x"a600", 2008=>x"9700", 2009=>x"9700",
---- 2010=>x"9700", 2011=>x"9c00", 2012=>x"9e00", 2013=>x"a000", 2014=>x"a500", 2015=>x"a500", 2016=>x"9900",
---- 2017=>x"9800", 2018=>x"9700", 2019=>x"9d00", 2020=>x"a000", 2021=>x"a200", 2022=>x"a600", 2023=>x"a700",
---- 2024=>x"9900", 2025=>x"9b00", 2026=>x"9900", 2027=>x"9c00", 2028=>x"a000", 2029=>x"a000", 2030=>x"a400",
---- 2031=>x"a300", 2032=>x"9a00", 2033=>x"9a00", 2034=>x"9a00", 2035=>x"9d00", 2036=>x"9c00", 2037=>x"5e00",
---- 2038=>x"a500", 2039=>x"a400", 2040=>x"9d00", 2041=>x"6100", 2042=>x"9d00", 2043=>x"9e00", 2044=>x"9e00",
---- 2045=>x"a100", 2046=>x"a300", 2047=>x"a800"),
---- 21 => (0=>x"9f00", 1=>x"a100", 2=>x"a000", 3=>x"9e00", 4=>x"9600", 5=>x"9700", 6=>x"9800", 7=>x"9800",
---- 8=>x"9f00", 9=>x"a000", 10=>x"a100", 11=>x"9d00", 12=>x"9600", 13=>x"9700", 14=>x"9700",
---- 15=>x"9800", 16=>x"9f00", 17=>x"a100", 18=>x"a200", 19=>x"9e00", 20=>x"9600", 21=>x"9800",
---- 22=>x"9800", 23=>x"9800", 24=>x"9d00", 25=>x"a000", 26=>x"a100", 27=>x"9d00", 28=>x"9a00",
---- 29=>x"9800", 30=>x"9800", 31=>x"9900", 32=>x"9a00", 33=>x"9d00", 34=>x"a100", 35=>x"a000",
---- 36=>x"9c00", 37=>x"9900", 38=>x"9900", 39=>x"9800", 40=>x"9800", 41=>x"9c00", 42=>x"a100",
---- 43=>x"a000", 44=>x"9c00", 45=>x"9b00", 46=>x"9a00", 47=>x"9b00", 48=>x"9800", 49=>x"9a00",
---- 50=>x"a100", 51=>x"a000", 52=>x"9f00", 53=>x"9d00", 54=>x"9a00", 55=>x"9d00", 56=>x"9700",
---- 57=>x"9900", 58=>x"9d00", 59=>x"a100", 60=>x"a200", 61=>x"a100", 62=>x"a000", 63=>x"9f00",
---- 64=>x"9300", 65=>x"9700", 66=>x"9b00", 67=>x"9d00", 68=>x"a000", 69=>x"a300", 70=>x"a200",
---- 71=>x"a100", 72=>x"8f00", 73=>x"9800", 74=>x"6500", 75=>x"9e00", 76=>x"a100", 77=>x"a400",
---- 78=>x"a100", 79=>x"a200", 80=>x"9200", 81=>x"9500", 82=>x"6500", 83=>x"6300", 84=>x"a000",
---- 85=>x"a400", 86=>x"a300", 87=>x"a300", 88=>x"9100", 89=>x"9700", 90=>x"9900", 91=>x"9b00",
---- 92=>x"a000", 93=>x"a100", 94=>x"a300", 95=>x"a400", 96=>x"8d00", 97=>x"9500", 98=>x"9900",
---- 99=>x"9e00", 100=>x"9f00", 101=>x"5c00", 102=>x"a300", 103=>x"a200", 104=>x"8d00", 105=>x"9100",
---- 106=>x"9900", 107=>x"9e00", 108=>x"a100", 109=>x"a100", 110=>x"a200", 111=>x"a200", 112=>x"8b00",
---- 113=>x"9300", 114=>x"9900", 115=>x"9c00", 116=>x"9f00", 117=>x"a000", 118=>x"a200", 119=>x"a100",
---- 120=>x"8a00", 121=>x"9200", 122=>x"9600", 123=>x"9a00", 124=>x"9e00", 125=>x"9c00", 126=>x"9e00",
---- 127=>x"a300", 128=>x"8800", 129=>x"8d00", 130=>x"9300", 131=>x"9900", 132=>x"9c00", 133=>x"9d00",
---- 134=>x"9e00", 135=>x"a000", 136=>x"8900", 137=>x"8d00", 138=>x"9300", 139=>x"9800", 140=>x"9900",
---- 141=>x"9b00", 142=>x"9e00", 143=>x"9f00", 144=>x"8900", 145=>x"8c00", 146=>x"8f00", 147=>x"9500",
---- 148=>x"9800", 149=>x"9a00", 150=>x"9c00", 151=>x"9c00", 152=>x"8700", 153=>x"8b00", 154=>x"8f00",
---- 155=>x"9400", 156=>x"9600", 157=>x"9800", 158=>x"9b00", 159=>x"9900", 160=>x"8500", 161=>x"8c00",
---- 162=>x"9000", 163=>x"9300", 164=>x"9400", 165=>x"9600", 166=>x"9a00", 167=>x"9b00", 168=>x"8600",
---- 169=>x"8a00", 170=>x"8f00", 171=>x"9000", 172=>x"9300", 173=>x"9500", 174=>x"9700", 175=>x"9900",
---- 176=>x"8200", 177=>x"8b00", 178=>x"8c00", 179=>x"9000", 180=>x"9200", 181=>x"9300", 182=>x"9400",
---- 183=>x"9700", 184=>x"8500", 185=>x"8a00", 186=>x"8d00", 187=>x"9100", 188=>x"9100", 189=>x"9200",
---- 190=>x"9200", 191=>x"9600", 192=>x"8200", 193=>x"8a00", 194=>x"8f00", 195=>x"9000", 196=>x"9000",
---- 197=>x"8e00", 198=>x"9100", 199=>x"9200", 200=>x"8500", 201=>x"8a00", 202=>x"8c00", 203=>x"9100",
---- 204=>x"9100", 205=>x"7000", 206=>x"9000", 207=>x"9100", 208=>x"8600", 209=>x"8b00", 210=>x"8d00",
---- 211=>x"9500", 212=>x"9000", 213=>x"9000", 214=>x"8f00", 215=>x"9200", 216=>x"8500", 217=>x"8a00",
---- 218=>x"8f00", 219=>x"9100", 220=>x"9200", 221=>x"8f00", 222=>x"9100", 223=>x"9000", 224=>x"8800",
---- 225=>x"8e00", 226=>x"8f00", 227=>x"9000", 228=>x"9200", 229=>x"9100", 230=>x"8f00", 231=>x"9000",
---- 232=>x"8400", 233=>x"8b00", 234=>x"8e00", 235=>x"9200", 236=>x"9200", 237=>x"9200", 238=>x"9000",
---- 239=>x"9200", 240=>x"8500", 241=>x"8c00", 242=>x"8f00", 243=>x"9200", 244=>x"9200", 245=>x"9200",
---- 246=>x"9000", 247=>x"9100", 248=>x"8900", 249=>x"7300", 250=>x"8f00", 251=>x"9200", 252=>x"9500",
---- 253=>x"9200", 254=>x"9100", 255=>x"9100", 256=>x"8600", 257=>x"8c00", 258=>x"9000", 259=>x"9400",
---- 260=>x"9700", 261=>x"9300", 262=>x"9200", 263=>x"9100", 264=>x"8700", 265=>x"8c00", 266=>x"9100",
---- 267=>x"9300", 268=>x"9700", 269=>x"9700", 270=>x"9500", 271=>x"9200", 272=>x"8900", 273=>x"8f00",
---- 274=>x"9300", 275=>x"9600", 276=>x"9900", 277=>x"9600", 278=>x"9600", 279=>x"9400", 280=>x"8700",
---- 281=>x"8e00", 282=>x"9300", 283=>x"9700", 284=>x"9900", 285=>x"9800", 286=>x"9600", 287=>x"9700",
---- 288=>x"8700", 289=>x"8f00", 290=>x"9200", 291=>x"9800", 292=>x"9900", 293=>x"9900", 294=>x"9900",
---- 295=>x"9600", 296=>x"8a00", 297=>x"9600", 298=>x"9500", 299=>x"9900", 300=>x"9700", 301=>x"9c00",
---- 302=>x"9d00", 303=>x"9b00", 304=>x"8b00", 305=>x"9300", 306=>x"9700", 307=>x"9a00", 308=>x"9b00",
---- 309=>x"9b00", 310=>x"9f00", 311=>x"9c00", 312=>x"8900", 313=>x"9100", 314=>x"9500", 315=>x"9800",
---- 316=>x"9e00", 317=>x"9b00", 318=>x"9d00", 319=>x"9b00", 320=>x"8700", 321=>x"9000", 322=>x"9500",
---- 323=>x"9900", 324=>x"9b00", 325=>x"9a00", 326=>x"9c00", 327=>x"9a00", 328=>x"8900", 329=>x"8f00",
---- 330=>x"9400", 331=>x"9600", 332=>x"9b00", 333=>x"9900", 334=>x"9b00", 335=>x"9a00", 336=>x"8500",
---- 337=>x"8e00", 338=>x"9300", 339=>x"9900", 340=>x"9d00", 341=>x"9900", 342=>x"9800", 343=>x"9900",
---- 344=>x"8500", 345=>x"8d00", 346=>x"9500", 347=>x"9b00", 348=>x"9d00", 349=>x"9900", 350=>x"9800",
---- 351=>x"9900", 352=>x"8500", 353=>x"8d00", 354=>x"9600", 355=>x"9900", 356=>x"9a00", 357=>x"9a00",
---- 358=>x"9900", 359=>x"9900", 360=>x"8500", 361=>x"8c00", 362=>x"9500", 363=>x"9a00", 364=>x"9c00",
---- 365=>x"9c00", 366=>x"9d00", 367=>x"9a00", 368=>x"8600", 369=>x"8d00", 370=>x"9500", 371=>x"9b00",
---- 372=>x"9d00", 373=>x"9b00", 374=>x"9a00", 375=>x"9b00", 376=>x"8700", 377=>x"8f00", 378=>x"9500",
---- 379=>x"9900", 380=>x"9d00", 381=>x"9a00", 382=>x"9b00", 383=>x"9800", 384=>x"8600", 385=>x"8d00",
---- 386=>x"9400", 387=>x"9b00", 388=>x"9b00", 389=>x"9a00", 390=>x"9c00", 391=>x"9800", 392=>x"8600",
---- 393=>x"8e00", 394=>x"9300", 395=>x"9a00", 396=>x"9b00", 397=>x"9a00", 398=>x"9b00", 399=>x"9c00",
---- 400=>x"8600", 401=>x"8f00", 402=>x"9600", 403=>x"9800", 404=>x"9c00", 405=>x"9a00", 406=>x"9a00",
---- 407=>x"9900", 408=>x"8600", 409=>x"8d00", 410=>x"9500", 411=>x"9b00", 412=>x"9c00", 413=>x"9a00",
---- 414=>x"9b00", 415=>x"9900", 416=>x"8200", 417=>x"8a00", 418=>x"9500", 419=>x"9800", 420=>x"9a00",
---- 421=>x"9900", 422=>x"9900", 423=>x"9a00", 424=>x"8400", 425=>x"8b00", 426=>x"9400", 427=>x"9700",
---- 428=>x"9a00", 429=>x"9a00", 430=>x"9900", 431=>x"9b00", 432=>x"8000", 433=>x"8c00", 434=>x"9300",
---- 435=>x"9700", 436=>x"9a00", 437=>x"9a00", 438=>x"9b00", 439=>x"9a00", 440=>x"8200", 441=>x"8c00",
---- 442=>x"9100", 443=>x"9700", 444=>x"9900", 445=>x"9800", 446=>x"9b00", 447=>x"9c00", 448=>x"8200",
---- 449=>x"8900", 450=>x"9400", 451=>x"9800", 452=>x"9700", 453=>x"9800", 454=>x"9900", 455=>x"9800",
---- 456=>x"8300", 457=>x"8b00", 458=>x"9300", 459=>x"9700", 460=>x"6900", 461=>x"9700", 462=>x"9900",
---- 463=>x"9900", 464=>x"8100", 465=>x"8b00", 466=>x"9300", 467=>x"9600", 468=>x"9800", 469=>x"9a00",
---- 470=>x"9a00", 471=>x"9900", 472=>x"7e00", 473=>x"8900", 474=>x"9200", 475=>x"9500", 476=>x"9700",
---- 477=>x"9900", 478=>x"9c00", 479=>x"9a00", 480=>x"7d00", 481=>x"8800", 482=>x"9700", 483=>x"9600",
---- 484=>x"9900", 485=>x"9800", 486=>x"9900", 487=>x"9b00", 488=>x"7b00", 489=>x"8900", 490=>x"8f00",
---- 491=>x"9b00", 492=>x"9c00", 493=>x"9a00", 494=>x"9d00", 495=>x"9c00", 496=>x"7b00", 497=>x"8600",
---- 498=>x"8d00", 499=>x"9c00", 500=>x"a000", 501=>x"9a00", 502=>x"9e00", 503=>x"9d00", 504=>x"7900",
---- 505=>x"8600", 506=>x"9000", 507=>x"9800", 508=>x"9b00", 509=>x"9900", 510=>x"9d00", 511=>x"9d00",
---- 512=>x"7100", 513=>x"8200", 514=>x"8f00", 515=>x"9600", 516=>x"9900", 517=>x"9b00", 518=>x"9c00",
---- 519=>x"9c00", 520=>x"9300", 521=>x"7f00", 522=>x"8c00", 523=>x"9600", 524=>x"9800", 525=>x"9900",
---- 526=>x"9b00", 527=>x"9c00", 528=>x"d500", 529=>x"a200", 530=>x"8500", 531=>x"9400", 532=>x"9600",
---- 533=>x"9700", 534=>x"9900", 535=>x"9900", 536=>x"da00", 537=>x"cf00", 538=>x"9a00", 539=>x"8f00",
---- 540=>x"9a00", 541=>x"9a00", 542=>x"9800", 543=>x"9700", 544=>x"cf00", 545=>x"d500", 546=>x"ba00",
---- 547=>x"8f00", 548=>x"9a00", 549=>x"9a00", 550=>x"9700", 551=>x"9500", 552=>x"cd00", 553=>x"d100",
---- 554=>x"cd00", 555=>x"9c00", 556=>x"9600", 557=>x"9a00", 558=>x"9600", 559=>x"9400", 560=>x"c200",
---- 561=>x"ca00", 562=>x"d000", 563=>x"a600", 564=>x"9200", 565=>x"9900", 566=>x"9700", 567=>x"9100",
---- 568=>x"b900", 569=>x"c100", 570=>x"ca00", 571=>x"bb00", 572=>x"9200", 573=>x"9200", 574=>x"9600",
---- 575=>x"a900", 576=>x"ba00", 577=>x"bb00", 578=>x"be00", 579=>x"cb00", 580=>x"a800", 581=>x"9800",
---- 582=>x"b800", 583=>x"d300", 584=>x"b900", 585=>x"b800", 586=>x"ba00", 587=>x"c100", 588=>x"c000",
---- 589=>x"c500", 590=>x"d300", 591=>x"cb00", 592=>x"b400", 593=>x"b200", 594=>x"ba00", 595=>x"c300",
---- 596=>x"cb00", 597=>x"c500", 598=>x"be00", 599=>x"c000", 600=>x"af00", 601=>x"c300", 602=>x"cc00",
---- 603=>x"c300", 604=>x"b900", 605=>x"ad00", 606=>x"b700", 607=>x"c700", 608=>x"cb00", 609=>x"c800",
---- 610=>x"b700", 611=>x"aa00", 612=>x"b900", 613=>x"c100", 614=>x"c700", 615=>x"c800", 616=>x"bd00",
---- 617=>x"b200", 618=>x"b700", 619=>x"bb00", 620=>x"c200", 621=>x"c800", 622=>x"ca00", 623=>x"d000",
---- 624=>x"b900", 625=>x"c000", 626=>x"c200", 627=>x"c600", 628=>x"ca00", 629=>x"ca00", 630=>x"cd00",
---- 631=>x"cb00", 632=>x"c200", 633=>x"c300", 634=>x"c800", 635=>x"ce00", 636=>x"cd00", 637=>x"c700",
---- 638=>x"c700", 639=>x"c700", 640=>x"c800", 641=>x"cc00", 642=>x"ce00", 643=>x"cb00", 644=>x"c900",
---- 645=>x"c600", 646=>x"be00", 647=>x"bf00", 648=>x"d100", 649=>x"cc00", 650=>x"c900", 651=>x"c500",
---- 652=>x"c200", 653=>x"c000", 654=>x"bf00", 655=>x"c200", 656=>x"c800", 657=>x"c500", 658=>x"c300",
---- 659=>x"c100", 660=>x"bd00", 661=>x"c100", 662=>x"c300", 663=>x"c300", 664=>x"bb00", 665=>x"b800",
---- 666=>x"be00", 667=>x"c000", 668=>x"be00", 669=>x"c200", 670=>x"c300", 671=>x"c600", 672=>x"b600",
---- 673=>x"b900", 674=>x"bd00", 675=>x"c100", 676=>x"c200", 677=>x"c300", 678=>x"c200", 679=>x"c700",
---- 680=>x"bd00", 681=>x"c000", 682=>x"c300", 683=>x"c400", 684=>x"c300", 685=>x"c300", 686=>x"c600",
---- 687=>x"c700", 688=>x"c000", 689=>x"c100", 690=>x"c300", 691=>x"c600", 692=>x"c600", 693=>x"c600",
---- 694=>x"c800", 695=>x"c600", 696=>x"c300", 697=>x"c000", 698=>x"c500", 699=>x"c800", 700=>x"c800",
---- 701=>x"c900", 702=>x"c900", 703=>x"c900", 704=>x"c300", 705=>x"c400", 706=>x"c600", 707=>x"c900",
---- 708=>x"c700", 709=>x"c900", 710=>x"c900", 711=>x"ca00", 712=>x"c400", 713=>x"c400", 714=>x"c700",
---- 715=>x"ca00", 716=>x"c700", 717=>x"c800", 718=>x"c800", 719=>x"c900", 720=>x"c400", 721=>x"c600",
---- 722=>x"c700", 723=>x"c800", 724=>x"c900", 725=>x"c900", 726=>x"c700", 727=>x"c800", 728=>x"c300",
---- 729=>x"c600", 730=>x"c600", 731=>x"c700", 732=>x"c800", 733=>x"c800", 734=>x"c800", 735=>x"c300",
---- 736=>x"c200", 737=>x"c600", 738=>x"c400", 739=>x"c300", 740=>x"c700", 741=>x"c900", 742=>x"cb00",
---- 743=>x"c800", 744=>x"c200", 745=>x"c400", 746=>x"c400", 747=>x"c600", 748=>x"c800", 749=>x"cc00",
---- 750=>x"ca00", 751=>x"c900", 752=>x"c400", 753=>x"c400", 754=>x"c400", 755=>x"c600", 756=>x"c600",
---- 757=>x"c600", 758=>x"c400", 759=>x"cd00", 760=>x"c300", 761=>x"c500", 762=>x"c400", 763=>x"c500",
---- 764=>x"c700", 765=>x"cb00", 766=>x"c900", 767=>x"af00", 768=>x"c200", 769=>x"c500", 770=>x"c600",
---- 771=>x"c600", 772=>x"ce00", 773=>x"bc00", 774=>x"8100", 775=>x"5500", 776=>x"c500", 777=>x"c700",
---- 778=>x"cf00", 779=>x"bd00", 780=>x"8100", 781=>x"5900", 782=>x"5500", 783=>x"5000", 784=>x"c800",
---- 785=>x"ca00", 786=>x"6e00", 787=>x"5e00", 788=>x"2d00", 789=>x"bf00", 790=>x"7900", 791=>x"6700",
---- 792=>x"b700", 793=>x"6200", 794=>x"2c00", 795=>x"5600", 796=>x"5b00", 797=>x"3f00", 798=>x"8100",
---- 799=>x"8400", 800=>x"5f00", 801=>x"2b00", 802=>x"2c00", 803=>x"5900", 804=>x"7700", 805=>x"4d00",
---- 806=>x"5c00", 807=>x"9300", 808=>x"4d00", 809=>x"5000", 810=>x"5100", 811=>x"4400", 812=>x"6000",
---- 813=>x"7100", 814=>x"5600", 815=>x"7100", 816=>x"6900", 817=>x"4a00", 818=>x"a500", 819=>x"6400",
---- 820=>x"4f00", 821=>x"5b00", 822=>x"6300", 823=>x"5600", 824=>x"8400", 825=>x"5d00", 826=>x"4c00",
---- 827=>x"5200", 828=>x"7300", 829=>x"6300", 830=>x"6400", 831=>x"6400", 832=>x"9600", 833=>x"6e00",
---- 834=>x"5d00", 835=>x"5000", 836=>x"5800", 837=>x"8400", 838=>x"6c00", 839=>x"5f00", 840=>x"ab00",
---- 841=>x"8600", 842=>x"6000", 843=>x"5800", 844=>x"4800", 845=>x"4b00", 846=>x"7400", 847=>x"5500",
---- 848=>x"b700", 849=>x"6800", 850=>x"7000", 851=>x"5800", 852=>x"4d00", 853=>x"3700", 854=>x"4a00",
---- 855=>x"6f00", 856=>x"b900", 857=>x"9f00", 858=>x"7700", 859=>x"6100", 860=>x"5400", 861=>x"4200",
---- 862=>x"2700", 863=>x"4500", 864=>x"b700", 865=>x"a500", 866=>x"8500", 867=>x"6300", 868=>x"5200",
---- 869=>x"4300", 870=>x"3000", 871=>x"2b00", 872=>x"be00", 873=>x"aa00", 874=>x"8800", 875=>x"6700",
---- 876=>x"5500", 877=>x"4000", 878=>x"2f00", 879=>x"2c00", 880=>x"c300", 881=>x"b100", 882=>x"9200",
---- 883=>x"6b00", 884=>x"5a00", 885=>x"4600", 886=>x"2800", 887=>x"2b00", 888=>x"c800", 889=>x"b900",
---- 890=>x"a000", 891=>x"7500", 892=>x"5e00", 893=>x"4d00", 894=>x"2c00", 895=>x"2a00", 896=>x"cd00",
---- 897=>x"c100", 898=>x"a800", 899=>x"8000", 900=>x"6500", 901=>x"5400", 902=>x"3300", 903=>x"2400",
---- 904=>x"d000", 905=>x"c300", 906=>x"b200", 907=>x"8e00", 908=>x"6b00", 909=>x"5600", 910=>x"3b00",
---- 911=>x"2e00", 912=>x"cf00", 913=>x"c700", 914=>x"b900", 915=>x"9700", 916=>x"7100", 917=>x"5500",
---- 918=>x"4100", 919=>x"2f00", 920=>x"d100", 921=>x"cc00", 922=>x"be00", 923=>x"9f00", 924=>x"7700",
---- 925=>x"5a00", 926=>x"4a00", 927=>x"2e00", 928=>x"d400", 929=>x"d000", 930=>x"c200", 931=>x"a600",
---- 932=>x"7e00", 933=>x"6300", 934=>x"4e00", 935=>x"3500", 936=>x"d600", 937=>x"d100", 938=>x"c800",
---- 939=>x"ac00", 940=>x"8a00", 941=>x"6700", 942=>x"5600", 943=>x"3d00", 944=>x"d500", 945=>x"d500",
---- 946=>x"cd00", 947=>x"b300", 948=>x"9300", 949=>x"6f00", 950=>x"a400", 951=>x"4b00", 952=>x"d500",
---- 953=>x"d100", 954=>x"cc00", 955=>x"be00", 956=>x"9c00", 957=>x"7500", 958=>x"5f00", 959=>x"5000",
---- 960=>x"d300", 961=>x"d200", 962=>x"cf00", 963=>x"c400", 964=>x"a200", 965=>x"7700", 966=>x"6000",
---- 967=>x"af00", 968=>x"d300", 969=>x"d000", 970=>x"3000", 971=>x"c600", 972=>x"a700", 973=>x"7f00",
---- 974=>x"5b00", 975=>x"4400", 976=>x"d100", 977=>x"cd00", 978=>x"c900", 979=>x"bd00", 980=>x"a300",
---- 981=>x"7800", 982=>x"b600", 983=>x"3600", 984=>x"ce00", 985=>x"c900", 986=>x"b900", 987=>x"a100",
---- 988=>x"8400", 989=>x"6200", 990=>x"4000", 991=>x"3500", 992=>x"bb00", 993=>x"a300", 994=>x"8900",
---- 995=>x"7600", 996=>x"6400", 997=>x"4e00", 998=>x"3b00", 999=>x"3600", 1000=>x"7300", 1001=>x"5e00",
---- 1002=>x"4f00", 1003=>x"4f00", 1004=>x"5d00", 1005=>x"5a00", 1006=>x"5500", 1007=>x"5300", 1008=>x"5c00",
---- 1009=>x"5e00", 1010=>x"6900", 1011=>x"6c00", 1012=>x"8600", 1013=>x"7700", 1014=>x"6c00", 1015=>x"6200",
---- 1016=>x"7b00", 1017=>x"9900", 1018=>x"6700", 1019=>x"6f00", 1020=>x"7500", 1021=>x"5f00", 1022=>x"5300",
---- 1023=>x"5000", 1024=>x"4d00", 1025=>x"3800", 1026=>x"3900", 1027=>x"4100", 1028=>x"4400", 1029=>x"4400",
---- 1030=>x"4700", 1031=>x"4400", 1032=>x"3000", 1033=>x"2f00", 1034=>x"3000", 1035=>x"3300", 1036=>x"3600",
---- 1037=>x"3800", 1038=>x"3d00", 1039=>x"4200", 1040=>x"3c00", 1041=>x"3100", 1042=>x"3100", 1043=>x"3400",
---- 1044=>x"3900", 1045=>x"3c00", 1046=>x"3600", 1047=>x"3d00", 1048=>x"7d00", 1049=>x"5800", 1050=>x"3400",
---- 1051=>x"2a00", 1052=>x"3200", 1053=>x"3700", 1054=>x"c700", 1055=>x"3800", 1056=>x"a500", 1057=>x"8500",
---- 1058=>x"4f00", 1059=>x"2c00", 1060=>x"2800", 1061=>x"3200", 1062=>x"3700", 1063=>x"3800", 1064=>x"aa00",
---- 1065=>x"9d00", 1066=>x"6600", 1067=>x"3c00", 1068=>x"2e00", 1069=>x"3500", 1070=>x"2f00", 1071=>x"3400",
---- 1072=>x"b000", 1073=>x"9d00", 1074=>x"7000", 1075=>x"4200", 1076=>x"2f00", 1077=>x"2c00", 1078=>x"d600",
---- 1079=>x"2e00", 1080=>x"b000", 1081=>x"9a00", 1082=>x"6d00", 1083=>x"4300", 1084=>x"3300", 1085=>x"2f00",
---- 1086=>x"2b00", 1087=>x"2f00", 1088=>x"ae00", 1089=>x"9500", 1090=>x"6700", 1091=>x"4200", 1092=>x"cc00",
---- 1093=>x"3200", 1094=>x"2f00", 1095=>x"3300", 1096=>x"9d00", 1097=>x"8000", 1098=>x"5a00", 1099=>x"3600",
---- 1100=>x"3600", 1101=>x"4100", 1102=>x"c900", 1103=>x"3700", 1104=>x"6700", 1105=>x"5700", 1106=>x"4000",
---- 1107=>x"3000", 1108=>x"4d00", 1109=>x"4f00", 1110=>x"3a00", 1111=>x"3800", 1112=>x"3d00", 1113=>x"4200",
---- 1114=>x"4c00", 1115=>x"5000", 1116=>x"5500", 1117=>x"5200", 1118=>x"3800", 1119=>x"3600", 1120=>x"5d00",
---- 1121=>x"5b00", 1122=>x"5400", 1123=>x"6100", 1124=>x"5a00", 1125=>x"5400", 1126=>x"3900", 1127=>x"3700",
---- 1128=>x"6800", 1129=>x"6700", 1130=>x"6300", 1131=>x"6800", 1132=>x"6200", 1133=>x"5a00", 1134=>x"3f00",
---- 1135=>x"3c00", 1136=>x"7a00", 1137=>x"7300", 1138=>x"7200", 1139=>x"7200", 1140=>x"6c00", 1141=>x"5c00",
---- 1142=>x"4300", 1143=>x"3f00", 1144=>x"7e00", 1145=>x"7700", 1146=>x"7400", 1147=>x"7200", 1148=>x"6e00",
---- 1149=>x"6100", 1150=>x"4500", 1151=>x"3e00", 1152=>x"8000", 1153=>x"7d00", 1154=>x"7a00", 1155=>x"7700",
---- 1156=>x"6e00", 1157=>x"6400", 1158=>x"4800", 1159=>x"3900", 1160=>x"8500", 1161=>x"7f00", 1162=>x"7c00",
---- 1163=>x"7900", 1164=>x"7400", 1165=>x"6800", 1166=>x"4c00", 1167=>x"3900", 1168=>x"8300", 1169=>x"8000",
---- 1170=>x"8100", 1171=>x"7c00", 1172=>x"7600", 1173=>x"6900", 1174=>x"4700", 1175=>x"3a00", 1176=>x"8200",
---- 1177=>x"8100", 1178=>x"8000", 1179=>x"7c00", 1180=>x"7900", 1181=>x"6900", 1182=>x"4500", 1183=>x"3a00",
---- 1184=>x"8500", 1185=>x"8100", 1186=>x"8000", 1187=>x"7e00", 1188=>x"7700", 1189=>x"6400", 1190=>x"3f00",
---- 1191=>x"3700", 1192=>x"8600", 1193=>x"8200", 1194=>x"8000", 1195=>x"7e00", 1196=>x"7400", 1197=>x"5e00",
---- 1198=>x"3e00", 1199=>x"3a00", 1200=>x"8500", 1201=>x"8200", 1202=>x"7f00", 1203=>x"7d00", 1204=>x"7400",
---- 1205=>x"5600", 1206=>x"3e00", 1207=>x"3700", 1208=>x"8700", 1209=>x"8200", 1210=>x"8000", 1211=>x"7a00",
---- 1212=>x"6f00", 1213=>x"5000", 1214=>x"3a00", 1215=>x"2a00", 1216=>x"8700", 1217=>x"8200", 1218=>x"8000",
---- 1219=>x"7b00", 1220=>x"6d00", 1221=>x"4a00", 1222=>x"3500", 1223=>x"2c00", 1224=>x"8500", 1225=>x"8200",
---- 1226=>x"7f00", 1227=>x"7b00", 1228=>x"6500", 1229=>x"4200", 1230=>x"2f00", 1231=>x"2a00", 1232=>x"8200",
---- 1233=>x"8400", 1234=>x"8000", 1235=>x"7300", 1236=>x"5b00", 1237=>x"4000", 1238=>x"2b00", 1239=>x"2e00",
---- 1240=>x"8300", 1241=>x"8200", 1242=>x"7d00", 1243=>x"6e00", 1244=>x"5700", 1245=>x"3300", 1246=>x"2600",
---- 1247=>x"3200", 1248=>x"8400", 1249=>x"8100", 1250=>x"7b00", 1251=>x"6700", 1252=>x"4c00", 1253=>x"2d00",
---- 1254=>x"2b00", 1255=>x"3000", 1256=>x"8100", 1257=>x"7e00", 1258=>x"7a00", 1259=>x"6500", 1260=>x"3a00",
---- 1261=>x"2800", 1262=>x"2b00", 1263=>x"3000", 1264=>x"8200", 1265=>x"7c00", 1266=>x"7400", 1267=>x"5900",
---- 1268=>x"2f00", 1269=>x"2b00", 1270=>x"2c00", 1271=>x"3500", 1272=>x"7f00", 1273=>x"7b00", 1274=>x"6f00",
---- 1275=>x"4100", 1276=>x"2700", 1277=>x"2b00", 1278=>x"2a00", 1279=>x"ce00", 1280=>x"7d00", 1281=>x"7a00",
---- 1282=>x"5800", 1283=>x"3100", 1284=>x"2700", 1285=>x"2b00", 1286=>x"2d00", 1287=>x"3400", 1288=>x"7d00",
---- 1289=>x"7000", 1290=>x"3d00", 1291=>x"2800", 1292=>x"2c00", 1293=>x"2d00", 1294=>x"2f00", 1295=>x"3700",
---- 1296=>x"7f00", 1297=>x"5b00", 1298=>x"2e00", 1299=>x"2d00", 1300=>x"2f00", 1301=>x"2b00", 1302=>x"3100",
---- 1303=>x"3600", 1304=>x"7600", 1305=>x"bc00", 1306=>x"d200", 1307=>x"3200", 1308=>x"3400", 1309=>x"2a00",
---- 1310=>x"3100", 1311=>x"3700", 1312=>x"6200", 1313=>x"3000", 1314=>x"2e00", 1315=>x"3400", 1316=>x"3200",
---- 1317=>x"2d00", 1318=>x"3200", 1319=>x"3900", 1320=>x"4600", 1321=>x"2d00", 1322=>x"2e00", 1323=>x"3000",
---- 1324=>x"2f00", 1325=>x"2e00", 1326=>x"3500", 1327=>x"3900", 1328=>x"3300", 1329=>x"3300", 1330=>x"2f00",
---- 1331=>x"2d00", 1332=>x"2e00", 1333=>x"3000", 1334=>x"3200", 1335=>x"3f00", 1336=>x"2e00", 1337=>x"3300",
---- 1338=>x"3100", 1339=>x"3100", 1340=>x"2f00", 1341=>x"2f00", 1342=>x"3b00", 1343=>x"4600", 1344=>x"3000",
---- 1345=>x"3200", 1346=>x"2f00", 1347=>x"2f00", 1348=>x"2e00", 1349=>x"2f00", 1350=>x"3e00", 1351=>x"4500",
---- 1352=>x"3000", 1353=>x"3200", 1354=>x"3000", 1355=>x"3200", 1356=>x"2d00", 1357=>x"3100", 1358=>x"3f00",
---- 1359=>x"4000", 1360=>x"2e00", 1361=>x"2e00", 1362=>x"3000", 1363=>x"3200", 1364=>x"2f00", 1365=>x"3200",
---- 1366=>x"4100", 1367=>x"3c00", 1368=>x"2d00", 1369=>x"3500", 1370=>x"ca00", 1371=>x"2f00", 1372=>x"2f00",
---- 1373=>x"3900", 1374=>x"3a00", 1375=>x"bf00", 1376=>x"2e00", 1377=>x"3b00", 1378=>x"3700", 1379=>x"2d00",
---- 1380=>x"3200", 1381=>x"3600", 1382=>x"3c00", 1383=>x"4500", 1384=>x"3200", 1385=>x"3500", 1386=>x"3100",
---- 1387=>x"3100", 1388=>x"3500", 1389=>x"3500", 1390=>x"4300", 1391=>x"4300", 1392=>x"3500", 1393=>x"2f00",
---- 1394=>x"3100", 1395=>x"3100", 1396=>x"3500", 1397=>x"3300", 1398=>x"4900", 1399=>x"3e00", 1400=>x"3800",
---- 1401=>x"3000", 1402=>x"2e00", 1403=>x"3100", 1404=>x"3600", 1405=>x"3c00", 1406=>x"4900", 1407=>x"3b00",
---- 1408=>x"3500", 1409=>x"2c00", 1410=>x"2b00", 1411=>x"3300", 1412=>x"3500", 1413=>x"4300", 1414=>x"4100",
---- 1415=>x"3600", 1416=>x"3300", 1417=>x"2e00", 1418=>x"2f00", 1419=>x"3400", 1420=>x"3b00", 1421=>x"4400",
---- 1422=>x"3800", 1423=>x"3c00", 1424=>x"3000", 1425=>x"2a00", 1426=>x"2c00", 1427=>x"3600", 1428=>x"3600",
---- 1429=>x"3500", 1430=>x"3300", 1431=>x"4100", 1432=>x"2e00", 1433=>x"2900", 1434=>x"2c00", 1435=>x"3300",
---- 1436=>x"4100", 1437=>x"3000", 1438=>x"2d00", 1439=>x"4100", 1440=>x"3100", 1441=>x"2e00", 1442=>x"3200",
---- 1443=>x"3100", 1444=>x"4000", 1445=>x"3100", 1446=>x"2f00", 1447=>x"4500", 1448=>x"3900", 1449=>x"3100",
---- 1450=>x"3700", 1451=>x"3400", 1452=>x"3f00", 1453=>x"3400", 1454=>x"3000", 1455=>x"4800", 1456=>x"3900",
---- 1457=>x"3700", 1458=>x"3500", 1459=>x"3500", 1460=>x"3900", 1461=>x"3400", 1462=>x"2f00", 1463=>x"5300",
---- 1464=>x"3a00", 1465=>x"4400", 1466=>x"3500", 1467=>x"3600", 1468=>x"3500", 1469=>x"3800", 1470=>x"2c00",
---- 1471=>x"5700", 1472=>x"3900", 1473=>x"3f00", 1474=>x"3400", 1475=>x"3400", 1476=>x"3200", 1477=>x"3500",
---- 1478=>x"2a00", 1479=>x"5300", 1480=>x"3700", 1481=>x"3d00", 1482=>x"3500", 1483=>x"3600", 1484=>x"3100",
---- 1485=>x"3400", 1486=>x"2c00", 1487=>x"5800", 1488=>x"3e00", 1489=>x"3f00", 1490=>x"3200", 1491=>x"3600",
---- 1492=>x"3100", 1493=>x"3300", 1494=>x"2f00", 1495=>x"6000", 1496=>x"3f00", 1497=>x"3400", 1498=>x"3700",
---- 1499=>x"4100", 1500=>x"2f00", 1501=>x"3200", 1502=>x"3600", 1503=>x"6000", 1504=>x"3e00", 1505=>x"2d00",
---- 1506=>x"3d00", 1507=>x"4000", 1508=>x"2e00", 1509=>x"3300", 1510=>x"3b00", 1511=>x"6400", 1512=>x"3600",
---- 1513=>x"2d00", 1514=>x"c700", 1515=>x"3700", 1516=>x"3000", 1517=>x"cc00", 1518=>x"3800", 1519=>x"6200",
---- 1520=>x"3200", 1521=>x"3200", 1522=>x"3500", 1523=>x"3400", 1524=>x"3300", 1525=>x"3400", 1526=>x"4000",
---- 1527=>x"6800", 1528=>x"3600", 1529=>x"3a00", 1530=>x"3500", 1531=>x"3400", 1532=>x"3700", 1533=>x"3400",
---- 1534=>x"4300", 1535=>x"6700", 1536=>x"3300", 1537=>x"3a00", 1538=>x"3800", 1539=>x"3300", 1540=>x"3400",
---- 1541=>x"3900", 1542=>x"4300", 1543=>x"6500", 1544=>x"3600", 1545=>x"3600", 1546=>x"3200", 1547=>x"3400",
---- 1548=>x"3100", 1549=>x"3e00", 1550=>x"4100", 1551=>x"6300", 1552=>x"3900", 1553=>x"3700", 1554=>x"3200",
---- 1555=>x"3600", 1556=>x"3000", 1557=>x"3e00", 1558=>x"3d00", 1559=>x"6100", 1560=>x"3500", 1561=>x"3100",
---- 1562=>x"d200", 1563=>x"3900", 1564=>x"3200", 1565=>x"3f00", 1566=>x"3e00", 1567=>x"5f00", 1568=>x"3200",
---- 1569=>x"2e00", 1570=>x"2c00", 1571=>x"3700", 1572=>x"3200", 1573=>x"3e00", 1574=>x"4900", 1575=>x"5900",
---- 1576=>x"3800", 1577=>x"3100", 1578=>x"3200", 1579=>x"3300", 1580=>x"3500", 1581=>x"4000", 1582=>x"5400",
---- 1583=>x"6100", 1584=>x"3400", 1585=>x"2a00", 1586=>x"2c00", 1587=>x"2800", 1588=>x"2e00", 1589=>x"3900",
---- 1590=>x"5000", 1591=>x"5600", 1592=>x"2a00", 1593=>x"2600", 1594=>x"2700", 1595=>x"2200", 1596=>x"2900",
---- 1597=>x"3700", 1598=>x"4d00", 1599=>x"5000", 1600=>x"5d00", 1601=>x"2b00", 1602=>x"2500", 1603=>x"2400",
---- 1604=>x"2800", 1605=>x"3900", 1606=>x"4b00", 1607=>x"5400", 1608=>x"c400", 1609=>x"8200", 1610=>x"3700",
---- 1611=>x"2300", 1612=>x"2600", 1613=>x"3c00", 1614=>x"4100", 1615=>x"4a00", 1616=>x"d500", 1617=>x"d300",
---- 1618=>x"9c00", 1619=>x"4800", 1620=>x"2700", 1621=>x"3400", 1622=>x"3500", 1623=>x"3f00", 1624=>x"d100",
---- 1625=>x"d400", 1626=>x"2800", 1627=>x"ae00", 1628=>x"4f00", 1629=>x"2e00", 1630=>x"d000", 1631=>x"3500",
---- 1632=>x"d300", 1633=>x"d200", 1634=>x"d400", 1635=>x"d800", 1636=>x"b400", 1637=>x"5500", 1638=>x"2900",
---- 1639=>x"3300", 1640=>x"d100", 1641=>x"d300", 1642=>x"d500", 1643=>x"d600", 1644=>x"db00", 1645=>x"b800",
---- 1646=>x"4f00", 1647=>x"3000", 1648=>x"d100", 1649=>x"d300", 1650=>x"d400", 1651=>x"d500", 1652=>x"d800",
---- 1653=>x"dc00", 1654=>x"ab00", 1655=>x"4200", 1656=>x"d100", 1657=>x"d100", 1658=>x"d400", 1659=>x"d600",
---- 1660=>x"d800", 1661=>x"d800", 1662=>x"dd00", 1663=>x"9c00", 1664=>x"d100", 1665=>x"d300", 1666=>x"d300",
---- 1667=>x"d500", 1668=>x"d800", 1669=>x"d900", 1670=>x"db00", 1671=>x"da00", 1672=>x"ce00", 1673=>x"d100",
---- 1674=>x"d200", 1675=>x"d400", 1676=>x"2900", 1677=>x"d900", 1678=>x"da00", 1679=>x"df00", 1680=>x"cc00",
---- 1681=>x"d000", 1682=>x"d000", 1683=>x"d100", 1684=>x"d700", 1685=>x"d800", 1686=>x"db00", 1687=>x"dd00",
---- 1688=>x"cd00", 1689=>x"d000", 1690=>x"cf00", 1691=>x"d200", 1692=>x"d500", 1693=>x"d500", 1694=>x"db00",
---- 1695=>x"de00", 1696=>x"ce00", 1697=>x"d000", 1698=>x"d000", 1699=>x"d100", 1700=>x"d500", 1701=>x"d700",
---- 1702=>x"da00", 1703=>x"2400", 1704=>x"ce00", 1705=>x"d100", 1706=>x"d200", 1707=>x"d300", 1708=>x"d500",
---- 1709=>x"d600", 1710=>x"d700", 1711=>x"dc00", 1712=>x"ce00", 1713=>x"d100", 1714=>x"d000", 1715=>x"d400",
---- 1716=>x"d500", 1717=>x"d300", 1718=>x"d800", 1719=>x"db00", 1720=>x"ce00", 1721=>x"d000", 1722=>x"cf00",
---- 1723=>x"d200", 1724=>x"d500", 1725=>x"d400", 1726=>x"d600", 1727=>x"d900", 1728=>x"cd00", 1729=>x"d000",
---- 1730=>x"d100", 1731=>x"d300", 1732=>x"d400", 1733=>x"d400", 1734=>x"d500", 1735=>x"d900", 1736=>x"ce00",
---- 1737=>x"ce00", 1738=>x"d300", 1739=>x"d200", 1740=>x"d100", 1741=>x"d600", 1742=>x"d600", 1743=>x"d900",
---- 1744=>x"cb00", 1745=>x"cf00", 1746=>x"cf00", 1747=>x"cf00", 1748=>x"d100", 1749=>x"d500", 1750=>x"d400",
---- 1751=>x"d600", 1752=>x"ca00", 1753=>x"cf00", 1754=>x"d100", 1755=>x"ce00", 1756=>x"d100", 1757=>x"d300",
---- 1758=>x"d400", 1759=>x"d500", 1760=>x"ca00", 1761=>x"d000", 1762=>x"ce00", 1763=>x"cf00", 1764=>x"d100",
---- 1765=>x"d300", 1766=>x"d400", 1767=>x"d400", 1768=>x"ca00", 1769=>x"cc00", 1770=>x"cd00", 1771=>x"cf00",
---- 1772=>x"d000", 1773=>x"d200", 1774=>x"2b00", 1775=>x"d400", 1776=>x"c900", 1777=>x"cc00", 1778=>x"cd00",
---- 1779=>x"ce00", 1780=>x"cf00", 1781=>x"d300", 1782=>x"d400", 1783=>x"d400", 1784=>x"c600", 1785=>x"ca00",
---- 1786=>x"cc00", 1787=>x"cd00", 1788=>x"cf00", 1789=>x"d100", 1790=>x"d200", 1791=>x"d300", 1792=>x"c500",
---- 1793=>x"c900", 1794=>x"cc00", 1795=>x"d000", 1796=>x"cf00", 1797=>x"d100", 1798=>x"d100", 1799=>x"d300",
---- 1800=>x"c700", 1801=>x"c800", 1802=>x"c900", 1803=>x"cd00", 1804=>x"cf00", 1805=>x"cd00", 1806=>x"d000",
---- 1807=>x"d200", 1808=>x"c600", 1809=>x"c800", 1810=>x"c900", 1811=>x"cb00", 1812=>x"cd00", 1813=>x"ce00",
---- 1814=>x"d000", 1815=>x"d200", 1816=>x"c300", 1817=>x"c800", 1818=>x"c800", 1819=>x"cb00", 1820=>x"cf00",
---- 1821=>x"cf00", 1822=>x"cf00", 1823=>x"d200", 1824=>x"c300", 1825=>x"c600", 1826=>x"c700", 1827=>x"c900",
---- 1828=>x"cd00", 1829=>x"2f00", 1830=>x"d000", 1831=>x"d300", 1832=>x"c200", 1833=>x"3a00", 1834=>x"c600",
---- 1835=>x"ca00", 1836=>x"cc00", 1837=>x"cf00", 1838=>x"2d00", 1839=>x"d100", 1840=>x"c200", 1841=>x"c400",
---- 1842=>x"c600", 1843=>x"ca00", 1844=>x"cb00", 1845=>x"cd00", 1846=>x"d000", 1847=>x"d300", 1848=>x"bf00",
---- 1849=>x"c200", 1850=>x"c300", 1851=>x"3700", 1852=>x"ca00", 1853=>x"cd00", 1854=>x"d100", 1855=>x"d200",
---- 1856=>x"bf00", 1857=>x"c000", 1858=>x"c100", 1859=>x"c800", 1860=>x"cc00", 1861=>x"ce00", 1862=>x"d000",
---- 1863=>x"d000", 1864=>x"be00", 1865=>x"bf00", 1866=>x"c400", 1867=>x"c800", 1868=>x"ca00", 1869=>x"cc00",
---- 1870=>x"cf00", 1871=>x"d000", 1872=>x"bc00", 1873=>x"bf00", 1874=>x"c500", 1875=>x"c700", 1876=>x"cb00",
---- 1877=>x"cb00", 1878=>x"ce00", 1879=>x"cf00", 1880=>x"bc00", 1881=>x"bd00", 1882=>x"c200", 1883=>x"c800",
---- 1884=>x"c800", 1885=>x"c900", 1886=>x"cf00", 1887=>x"ce00", 1888=>x"b800", 1889=>x"ba00", 1890=>x"bf00",
---- 1891=>x"c500", 1892=>x"c500", 1893=>x"c900", 1894=>x"cb00", 1895=>x"cd00", 1896=>x"b800", 1897=>x"bb00",
---- 1898=>x"c000", 1899=>x"3c00", 1900=>x"c400", 1901=>x"c700", 1902=>x"ca00", 1903=>x"ce00", 1904=>x"b700",
---- 1905=>x"ba00", 1906=>x"bf00", 1907=>x"c200", 1908=>x"c400", 1909=>x"c600", 1910=>x"c900", 1911=>x"cb00",
---- 1912=>x"b300", 1913=>x"ba00", 1914=>x"4100", 1915=>x"c100", 1916=>x"c500", 1917=>x"c700", 1918=>x"c700",
---- 1919=>x"cb00", 1920=>x"b300", 1921=>x"b900", 1922=>x"bb00", 1923=>x"c000", 1924=>x"c200", 1925=>x"c400",
---- 1926=>x"c800", 1927=>x"cb00", 1928=>x"b100", 1929=>x"b500", 1930=>x"b700", 1931=>x"bd00", 1932=>x"c000",
---- 1933=>x"c200", 1934=>x"c600", 1935=>x"c900", 1936=>x"ad00", 1937=>x"b000", 1938=>x"b600", 1939=>x"ba00",
---- 1940=>x"bf00", 1941=>x"c000", 1942=>x"c300", 1943=>x"c700", 1944=>x"ac00", 1945=>x"b100", 1946=>x"b300",
---- 1947=>x"b800", 1948=>x"bd00", 1949=>x"be00", 1950=>x"c200", 1951=>x"c500", 1952=>x"ad00", 1953=>x"af00",
---- 1954=>x"b200", 1955=>x"b700", 1956=>x"b900", 1957=>x"be00", 1958=>x"c100", 1959=>x"c400", 1960=>x"af00",
---- 1961=>x"af00", 1962=>x"b100", 1963=>x"b400", 1964=>x"b900", 1965=>x"bd00", 1966=>x"c000", 1967=>x"c200",
---- 1968=>x"b000", 1969=>x"b100", 1970=>x"b200", 1971=>x"b500", 1972=>x"b700", 1973=>x"ba00", 1974=>x"be00",
---- 1975=>x"bf00", 1976=>x"a900", 1977=>x"b000", 1978=>x"b300", 1979=>x"b700", 1980=>x"b900", 1981=>x"bb00",
---- 1982=>x"bd00", 1983=>x"bf00", 1984=>x"a900", 1985=>x"af00", 1986=>x"ae00", 1987=>x"b300", 1988=>x"b600",
---- 1989=>x"ba00", 1990=>x"bc00", 1991=>x"bd00", 1992=>x"a700", 1993=>x"aa00", 1994=>x"ab00", 1995=>x"b100",
---- 1996=>x"b300", 1997=>x"b300", 1998=>x"ba00", 1999=>x"bb00", 2000=>x"a800", 2001=>x"a900", 2002=>x"ad00",
---- 2003=>x"b200", 2004=>x"b400", 2005=>x"b300", 2006=>x"b800", 2007=>x"bb00", 2008=>x"aa00", 2009=>x"a900",
---- 2010=>x"ac00", 2011=>x"b000", 2012=>x"b400", 2013=>x"b500", 2014=>x"b600", 2015=>x"ba00", 2016=>x"a800",
---- 2017=>x"a500", 2018=>x"ad00", 2019=>x"b200", 2020=>x"b100", 2021=>x"b200", 2022=>x"b600", 2023=>x"b900",
---- 2024=>x"a200", 2025=>x"a600", 2026=>x"aa00", 2027=>x"af00", 2028=>x"ae00", 2029=>x"b200", 2030=>x"b800",
---- 2031=>x"4400", 2032=>x"a400", 2033=>x"a400", 2034=>x"a900", 2035=>x"ab00", 2036=>x"ad00", 2037=>x"b100",
---- 2038=>x"b500", 2039=>x"b900", 2040=>x"a500", 2041=>x"a400", 2042=>x"a900", 2043=>x"a800", 2044=>x"ae00",
---- 2045=>x"5100", 2046=>x"b100", 2047=>x"b600"),
---- 22 => (0=>x"9a00", 1=>x"9a00", 2=>x"9c00", 3=>x"9a00", 4=>x"9e00", 5=>x"9c00", 6=>x"9a00", 7=>x"9800",
---- 8=>x"9900", 9=>x"9c00", 10=>x"9b00", 11=>x"9a00", 12=>x"9e00", 13=>x"9e00", 14=>x"9a00",
---- 15=>x"9900", 16=>x"9900", 17=>x"9a00", 18=>x"9b00", 19=>x"9b00", 20=>x"9c00", 21=>x"9c00",
---- 22=>x"9b00", 23=>x"9900", 24=>x"9500", 25=>x"9900", 26=>x"9900", 27=>x"9800", 28=>x"9900",
---- 29=>x"9b00", 30=>x"9b00", 31=>x"9900", 32=>x"9900", 33=>x"9c00", 34=>x"9b00", 35=>x"9a00",
---- 36=>x"9b00", 37=>x"9b00", 38=>x"9a00", 39=>x"9c00", 40=>x"9a00", 41=>x"9d00", 42=>x"9e00",
---- 43=>x"9d00", 44=>x"9f00", 45=>x"9c00", 46=>x"9a00", 47=>x"6300", 48=>x"9b00", 49=>x"9d00",
---- 50=>x"a000", 51=>x"9e00", 52=>x"a000", 53=>x"9f00", 54=>x"9f00", 55=>x"9e00", 56=>x"9e00",
---- 57=>x"a100", 58=>x"a000", 59=>x"a200", 60=>x"a200", 61=>x"a200", 62=>x"a200", 63=>x"9e00",
---- 64=>x"9e00", 65=>x"a000", 66=>x"a100", 67=>x"a200", 68=>x"a100", 69=>x"a200", 70=>x"a200",
---- 71=>x"9f00", 72=>x"a200", 73=>x"9f00", 74=>x"a100", 75=>x"a300", 76=>x"a400", 77=>x"a000",
---- 78=>x"a200", 79=>x"a300", 80=>x"a300", 81=>x"9f00", 82=>x"a100", 83=>x"a300", 84=>x"a400",
---- 85=>x"a400", 86=>x"a200", 87=>x"a200", 88=>x"a100", 89=>x"a100", 90=>x"a000", 91=>x"a100",
---- 92=>x"a000", 93=>x"a200", 94=>x"a100", 95=>x"a100", 96=>x"a200", 97=>x"a500", 98=>x"a000",
---- 99=>x"9e00", 100=>x"a000", 101=>x"a100", 102=>x"a000", 103=>x"a000", 104=>x"a200", 105=>x"a300",
---- 106=>x"a000", 107=>x"9e00", 108=>x"9e00", 109=>x"9f00", 110=>x"9f00", 111=>x"9f00", 112=>x"a200",
---- 113=>x"a100", 114=>x"a100", 115=>x"a000", 116=>x"9d00", 117=>x"9e00", 118=>x"a000", 119=>x"9c00",
---- 120=>x"a000", 121=>x"a000", 122=>x"9f00", 123=>x"9c00", 124=>x"a000", 125=>x"9d00", 126=>x"a100",
---- 127=>x"9e00", 128=>x"a000", 129=>x"a200", 130=>x"9e00", 131=>x"9d00", 132=>x"9f00", 133=>x"9e00",
---- 134=>x"a000", 135=>x"a000", 136=>x"9f00", 137=>x"a100", 138=>x"9f00", 139=>x"9e00", 140=>x"9e00",
---- 141=>x"9d00", 142=>x"9f00", 143=>x"9e00", 144=>x"6300", 145=>x"9e00", 146=>x"9d00", 147=>x"9d00",
---- 148=>x"9c00", 149=>x"9d00", 150=>x"9d00", 151=>x"9d00", 152=>x"9c00", 153=>x"9e00", 154=>x"9d00",
---- 155=>x"a000", 156=>x"9c00", 157=>x"9d00", 158=>x"9d00", 159=>x"9d00", 160=>x"9900", 161=>x"9e00",
---- 162=>x"9a00", 163=>x"9e00", 164=>x"9d00", 165=>x"9c00", 166=>x"9d00", 167=>x"9c00", 168=>x"9a00",
---- 169=>x"9a00", 170=>x"9b00", 171=>x"9d00", 172=>x"9e00", 173=>x"9900", 174=>x"9c00", 175=>x"9c00",
---- 176=>x"9800", 177=>x"9700", 178=>x"9a00", 179=>x"9c00", 180=>x"9c00", 181=>x"9c00", 182=>x"9b00",
---- 183=>x"9800", 184=>x"9600", 185=>x"9500", 186=>x"9900", 187=>x"9c00", 188=>x"9a00", 189=>x"9b00",
---- 190=>x"9a00", 191=>x"9a00", 192=>x"9500", 193=>x"9600", 194=>x"9800", 195=>x"9a00", 196=>x"9a00",
---- 197=>x"9b00", 198=>x"9b00", 199=>x"9c00", 200=>x"9000", 201=>x"9600", 202=>x"9500", 203=>x"9700",
---- 204=>x"9a00", 205=>x"9a00", 206=>x"9a00", 207=>x"9b00", 208=>x"9200", 209=>x"9400", 210=>x"9400",
---- 211=>x"9700", 212=>x"9700", 213=>x"9a00", 214=>x"9a00", 215=>x"9a00", 216=>x"9300", 217=>x"9400",
---- 218=>x"9400", 219=>x"9600", 220=>x"9700", 221=>x"9800", 222=>x"9a00", 223=>x"9800", 224=>x"9100",
---- 225=>x"9500", 226=>x"9400", 227=>x"9400", 228=>x"9900", 229=>x"9800", 230=>x"9900", 231=>x"9700",
---- 232=>x"9100", 233=>x"9300", 234=>x"9300", 235=>x"9400", 236=>x"9300", 237=>x"9500", 238=>x"9700",
---- 239=>x"9800", 240=>x"8f00", 241=>x"9200", 242=>x"9400", 243=>x"9400", 244=>x"9000", 245=>x"9200",
---- 246=>x"9700", 247=>x"9a00", 248=>x"8f00", 249=>x"9200", 250=>x"9400", 251=>x"9300", 252=>x"9300",
---- 253=>x"9200", 254=>x"9400", 255=>x"9500", 256=>x"9100", 257=>x"9200", 258=>x"9100", 259=>x"9200",
---- 260=>x"9200", 261=>x"9100", 262=>x"9200", 263=>x"9300", 264=>x"9100", 265=>x"9000", 266=>x"9000",
---- 267=>x"9000", 268=>x"8f00", 269=>x"9000", 270=>x"9000", 271=>x"8e00", 272=>x"9200", 273=>x"9000",
---- 274=>x"8f00", 275=>x"8f00", 276=>x"8e00", 277=>x"9000", 278=>x"8e00", 279=>x"8c00", 280=>x"9600",
---- 281=>x"9300", 282=>x"9300", 283=>x"8d00", 284=>x"8a00", 285=>x"8c00", 286=>x"8c00", 287=>x"8b00",
---- 288=>x"9700", 289=>x"9400", 290=>x"9200", 291=>x"8e00", 292=>x"8800", 293=>x"8500", 294=>x"8600",
---- 295=>x"8600", 296=>x"9700", 297=>x"9400", 298=>x"9500", 299=>x"8f00", 300=>x"8800", 301=>x"8400",
---- 302=>x"8100", 303=>x"7f00", 304=>x"9700", 305=>x"9800", 306=>x"9700", 307=>x"8e00", 308=>x"8700",
---- 309=>x"8000", 310=>x"7a00", 311=>x"7600", 312=>x"9800", 313=>x"9800", 314=>x"9900", 315=>x"9200",
---- 316=>x"8900", 317=>x"7d00", 318=>x"7700", 319=>x"6c00", 320=>x"9900", 321=>x"9800", 322=>x"9900",
---- 323=>x"9200", 324=>x"8b00", 325=>x"7f00", 326=>x"7100", 327=>x"6400", 328=>x"6600", 329=>x"9a00",
---- 330=>x"9a00", 331=>x"9200", 332=>x"8f00", 333=>x"8300", 334=>x"7300", 335=>x"5e00", 336=>x"9700",
---- 337=>x"9900", 338=>x"9800", 339=>x"9100", 340=>x"8d00", 341=>x"8300", 342=>x"7500", 343=>x"5d00",
---- 344=>x"9900", 345=>x"9b00", 346=>x"9800", 347=>x"9200", 348=>x"8d00", 349=>x"8500", 350=>x"7700",
---- 351=>x"5c00", 352=>x"9800", 353=>x"9800", 354=>x"9800", 355=>x"9300", 356=>x"8f00", 357=>x"8500",
---- 358=>x"7a00", 359=>x"6400", 360=>x"9700", 361=>x"9800", 362=>x"9800", 363=>x"9700", 364=>x"9100",
---- 365=>x"8600", 366=>x"7a00", 367=>x"6600", 368=>x"9b00", 369=>x"9a00", 370=>x"9a00", 371=>x"9500",
---- 372=>x"9200", 373=>x"8d00", 374=>x"7e00", 375=>x"6a00", 376=>x"9a00", 377=>x"9b00", 378=>x"9a00",
---- 379=>x"9500", 380=>x"8f00", 381=>x"8700", 382=>x"7b00", 383=>x"6500", 384=>x"9800", 385=>x"9a00",
---- 386=>x"9800", 387=>x"9600", 388=>x"9200", 389=>x"8900", 390=>x"7b00", 391=>x"6400", 392=>x"9900",
---- 393=>x"9900", 394=>x"9900", 395=>x"9700", 396=>x"9300", 397=>x"8900", 398=>x"7c00", 399=>x"6400",
---- 400=>x"9800", 401=>x"9900", 402=>x"9b00", 403=>x"a100", 404=>x"9100", 405=>x"8700", 406=>x"7a00",
---- 407=>x"6500", 408=>x"9800", 409=>x"9a00", 410=>x"9c00", 411=>x"9800", 412=>x"8f00", 413=>x"8700",
---- 414=>x"7700", 415=>x"6600", 416=>x"9900", 417=>x"9900", 418=>x"9b00", 419=>x"9900", 420=>x"9000",
---- 421=>x"8800", 422=>x"7900", 423=>x"6700", 424=>x"9a00", 425=>x"9900", 426=>x"9900", 427=>x"9700",
---- 428=>x"9100", 429=>x"8700", 430=>x"7d00", 431=>x"6c00", 432=>x"9a00", 433=>x"9a00", 434=>x"9900",
---- 435=>x"9600", 436=>x"9000", 437=>x"8600", 438=>x"7b00", 439=>x"6900", 440=>x"9b00", 441=>x"9a00",
---- 442=>x"9900", 443=>x"9600", 444=>x"9000", 445=>x"8600", 446=>x"7a00", 447=>x"6700", 448=>x"6600",
---- 449=>x"9900", 450=>x"9b00", 451=>x"9b00", 452=>x"6d00", 453=>x"8600", 454=>x"7b00", 455=>x"6b00",
---- 456=>x"9a00", 457=>x"9900", 458=>x"9800", 459=>x"9a00", 460=>x"9400", 461=>x"8700", 462=>x"8100",
---- 463=>x"6700", 464=>x"9a00", 465=>x"9c00", 466=>x"9800", 467=>x"9a00", 468=>x"9400", 469=>x"8700",
---- 470=>x"7900", 471=>x"6c00", 472=>x"9800", 473=>x"9b00", 474=>x"9900", 475=>x"9800", 476=>x"9200",
---- 477=>x"8800", 478=>x"7800", 479=>x"6600", 480=>x"9900", 481=>x"9a00", 482=>x"9a00", 483=>x"9800",
---- 484=>x"9300", 485=>x"8800", 486=>x"7700", 487=>x"6500", 488=>x"9b00", 489=>x"9b00", 490=>x"9800",
---- 491=>x"9800", 492=>x"9200", 493=>x"8600", 494=>x"7a00", 495=>x"6500", 496=>x"9d00", 497=>x"9c00",
---- 498=>x"9b00", 499=>x"9700", 500=>x"9100", 501=>x"8600", 502=>x"7500", 503=>x"6000", 504=>x"9d00",
---- 505=>x"9b00", 506=>x"9b00", 507=>x"9500", 508=>x"8f00", 509=>x"8100", 510=>x"6e00", 511=>x"5f00",
---- 512=>x"9a00", 513=>x"9c00", 514=>x"9900", 515=>x"9200", 516=>x"8c00", 517=>x"7a00", 518=>x"6800",
---- 519=>x"5300", 520=>x"9b00", 521=>x"9a00", 522=>x"9400", 523=>x"9200", 524=>x"8800", 525=>x"7700",
---- 526=>x"6000", 527=>x"4700", 528=>x"9a00", 529=>x"9700", 530=>x"9400", 531=>x"8f00", 532=>x"8400",
---- 533=>x"6e00", 534=>x"5500", 535=>x"6000", 536=>x"9600", 537=>x"9600", 538=>x"9000", 539=>x"8700",
---- 540=>x"7c00", 541=>x"7300", 542=>x"9100", 543=>x"c600", 544=>x"9600", 545=>x"9400", 546=>x"8b00",
---- 547=>x"8700", 548=>x"6200", 549=>x"bb00", 550=>x"da00", 551=>x"d600", 552=>x"8e00", 553=>x"8d00",
---- 554=>x"9a00", 555=>x"bb00", 556=>x"d700", 557=>x"d700", 558=>x"c700", 559=>x"bc00", 560=>x"9300",
---- 561=>x"ab00", 562=>x"c900", 563=>x"d600", 564=>x"c900", 565=>x"be00", 566=>x"ba00", 567=>x"ba00",
---- 568=>x"c100", 569=>x"d200", 570=>x"cd00", 571=>x"c400", 572=>x"c100", 573=>x"bf00", 574=>x"bd00",
---- 575=>x"bf00", 576=>x"d100", 577=>x"be00", 578=>x"b800", 579=>x"bf00", 580=>x"bf00", 581=>x"c400",
---- 582=>x"c900", 583=>x"d000", 584=>x"c000", 585=>x"bb00", 586=>x"be00", 587=>x"be00", 588=>x"c500",
---- 589=>x"cf00", 590=>x"d000", 591=>x"cd00", 592=>x"c300", 593=>x"c300", 594=>x"c600", 595=>x"ce00",
---- 596=>x"d200", 597=>x"d100", 598=>x"cc00", 599=>x"c800", 600=>x"c400", 601=>x"c600", 602=>x"cf00",
---- 603=>x"d300", 604=>x"d100", 605=>x"ce00", 606=>x"3b00", 607=>x"c100", 608=>x"cb00", 609=>x"cf00",
---- 610=>x"cf00", 611=>x"ce00", 612=>x"cd00", 613=>x"c600", 614=>x"c100", 615=>x"c700", 616=>x"cf00",
---- 617=>x"cb00", 618=>x"cb00", 619=>x"ca00", 620=>x"c600", 621=>x"c400", 622=>x"3a00", 623=>x"c900",
---- 624=>x"c600", 625=>x"c400", 626=>x"c400", 627=>x"c300", 628=>x"c400", 629=>x"c500", 630=>x"c400",
---- 631=>x"c900", 632=>x"c000", 633=>x"bc00", 634=>x"c000", 635=>x"c000", 636=>x"c400", 637=>x"c300",
---- 638=>x"c600", 639=>x"c800", 640=>x"c300", 641=>x"c100", 642=>x"be00", 643=>x"c200", 644=>x"c500",
---- 645=>x"c500", 646=>x"c900", 647=>x"c900", 648=>x"c200", 649=>x"c000", 650=>x"bf00", 651=>x"c500",
---- 652=>x"c600", 653=>x"c800", 654=>x"c900", 655=>x"c900", 656=>x"c200", 657=>x"c300", 658=>x"c300",
---- 659=>x"c700", 660=>x"c800", 661=>x"ca00", 662=>x"c900", 663=>x"cc00", 664=>x"c300", 665=>x"3b00",
---- 666=>x"c700", 667=>x"c900", 668=>x"ca00", 669=>x"cb00", 670=>x"cc00", 671=>x"cc00", 672=>x"c400",
---- 673=>x"c600", 674=>x"ca00", 675=>x"cb00", 676=>x"cc00", 677=>x"cc00", 678=>x"cb00", 679=>x"cb00",
---- 680=>x"c700", 681=>x"c900", 682=>x"cd00", 683=>x"ca00", 684=>x"cc00", 685=>x"ca00", 686=>x"cb00",
---- 687=>x"cc00", 688=>x"c700", 689=>x"ca00", 690=>x"c900", 691=>x"cd00", 692=>x"cd00", 693=>x"ca00",
---- 694=>x"cc00", 695=>x"cc00", 696=>x"c900", 697=>x"cb00", 698=>x"cb00", 699=>x"cd00", 700=>x"cb00",
---- 701=>x"3500", 702=>x"cc00", 703=>x"cc00", 704=>x"c900", 705=>x"ca00", 706=>x"cc00", 707=>x"ce00",
---- 708=>x"ca00", 709=>x"ca00", 710=>x"cb00", 711=>x"cb00", 712=>x"c700", 713=>x"cb00", 714=>x"ce00",
---- 715=>x"cd00", 716=>x"cb00", 717=>x"ce00", 718=>x"cc00", 719=>x"cb00", 720=>x"c600", 721=>x"cd00",
---- 722=>x"d000", 723=>x"cc00", 724=>x"cc00", 725=>x"cf00", 726=>x"d200", 727=>x"d200", 728=>x"c300",
---- 729=>x"d000", 730=>x"cc00", 731=>x"cc00", 732=>x"d300", 733=>x"d300", 734=>x"c000", 735=>x"9800",
---- 736=>x"cb00", 737=>x"cf00", 738=>x"d000", 739=>x"d500", 740=>x"bf00", 741=>x"8900", 742=>x"6900",
---- 743=>x"5400", 744=>x"ce00", 745=>x"d500", 746=>x"cf00", 747=>x"a600", 748=>x"6800", 749=>x"5300",
---- 750=>x"5b00", 751=>x"5c00", 752=>x"c900", 753=>x"ad00", 754=>x"9600", 755=>x"7700", 756=>x"5e00",
---- 757=>x"5e00", 758=>x"6100", 759=>x"5c00", 760=>x"7f00", 761=>x"5d00", 762=>x"8100", 763=>x"8600",
---- 764=>x"7300", 765=>x"6000", 766=>x"6000", 767=>x"5900", 768=>x"6600", 769=>x"6900", 770=>x"8400",
---- 771=>x"8c00", 772=>x"8100", 773=>x"8c00", 774=>x"7200", 775=>x"7b00", 776=>x"6a00", 777=>x"6700",
---- 778=>x"7a00", 779=>x"8d00", 780=>x"9200", 781=>x"9c00", 782=>x"9e00", 783=>x"a200", 784=>x"6500",
---- 785=>x"6a00", 786=>x"6c00", 787=>x"8d00", 788=>x"9900", 789=>x"a700", 790=>x"a300", 791=>x"a500",
---- 792=>x"6800", 793=>x"7700", 794=>x"6a00", 795=>x"8600", 796=>x"9800", 797=>x"a400", 798=>x"a000",
---- 799=>x"a800", 800=>x"7200", 801=>x"7800", 802=>x"7800", 803=>x"7600", 804=>x"9500", 805=>x"9700",
---- 806=>x"9d00", 807=>x"ab00", 808=>x"8c00", 809=>x"7200", 810=>x"7f00", 811=>x"6b00", 812=>x"8800",
---- 813=>x"9800", 814=>x"9a00", 815=>x"a700", 816=>x"7f00", 817=>x"8100", 818=>x"7500", 819=>x"6a00",
---- 820=>x"7900", 821=>x"9700", 822=>x"9800", 823=>x"a600", 824=>x"7400", 825=>x"8b00", 826=>x"7b00",
---- 827=>x"7800", 828=>x"7a00", 829=>x"9400", 830=>x"9c00", 831=>x"b000", 832=>x"5900", 833=>x"8000",
---- 834=>x"8900", 835=>x"8300", 836=>x"7f00", 837=>x"9000", 838=>x"a400", 839=>x"bb00", 840=>x"4900",
---- 841=>x"5300", 842=>x"8b00", 843=>x"8700", 844=>x"8200", 845=>x"8a00", 846=>x"a200", 847=>x"9f00",
---- 848=>x"5b00", 849=>x"4500", 850=>x"6e00", 851=>x"8a00", 852=>x"8700", 853=>x"8f00", 854=>x"9a00",
---- 855=>x"8700", 856=>x"6300", 857=>x"4a00", 858=>x"5100", 859=>x"8300", 860=>x"8500", 861=>x"9300",
---- 862=>x"9a00", 863=>x"8e00", 864=>x"5e00", 865=>x"5600", 866=>x"b300", 867=>x"7700", 868=>x"8600",
---- 869=>x"8900", 870=>x"9700", 871=>x"9200", 872=>x"c600", 873=>x"5600", 874=>x"b800", 875=>x"6300",
---- 876=>x"8e00", 877=>x"8900", 878=>x"9900", 879=>x"9800", 880=>x"2900", 881=>x"5100", 882=>x"4900",
---- 883=>x"5100", 884=>x"9200", 885=>x"9200", 886=>x"a200", 887=>x"9c00", 888=>x"2e00", 889=>x"3f00",
---- 890=>x"4c00", 891=>x"4700", 892=>x"8b00", 893=>x"9b00", 894=>x"a700", 895=>x"9900", 896=>x"2a00",
---- 897=>x"3200", 898=>x"4a00", 899=>x"4300", 900=>x"6f00", 901=>x"9f00", 902=>x"ac00", 903=>x"9c00",
---- 904=>x"2800", 905=>x"2900", 906=>x"3a00", 907=>x"4500", 908=>x"4f00", 909=>x"9800", 910=>x"a400",
---- 911=>x"a500", 912=>x"2400", 913=>x"2500", 914=>x"2e00", 915=>x"4800", 916=>x"4400", 917=>x"8d00",
---- 918=>x"a600", 919=>x"a200", 920=>x"2200", 921=>x"2400", 922=>x"2800", 923=>x"4700", 924=>x"4400",
---- 925=>x"8200", 926=>x"ae00", 927=>x"6100", 928=>x"2700", 929=>x"2600", 930=>x"2900", 931=>x"3800",
---- 932=>x"4700", 933=>x"9500", 934=>x"b200", 935=>x"a000", 936=>x"2d00", 937=>x"2b00", 938=>x"2900",
---- 939=>x"3000", 940=>x"4700", 941=>x"5700", 942=>x"a800", 943=>x"aa00", 944=>x"3100", 945=>x"2c00",
---- 946=>x"2800", 947=>x"2700", 948=>x"4b00", 949=>x"5500", 950=>x"9700", 951=>x"b100", 952=>x"3300",
---- 953=>x"2700", 954=>x"2900", 955=>x"2700", 956=>x"4200", 957=>x"5100", 958=>x"8d00", 959=>x"b500",
---- 960=>x"3100", 961=>x"2600", 962=>x"2b00", 963=>x"2900", 964=>x"3d00", 965=>x"4a00", 966=>x"7b00",
---- 967=>x"b600", 968=>x"3000", 969=>x"2700", 970=>x"2800", 971=>x"d600", 972=>x"3800", 973=>x"4100",
---- 974=>x"7100", 975=>x"b800", 976=>x"2f00", 977=>x"2a00", 978=>x"2700", 979=>x"2700", 980=>x"3200",
---- 981=>x"4300", 982=>x"6000", 983=>x"b800", 984=>x"2d00", 985=>x"2700", 986=>x"2600", 987=>x"2600",
---- 988=>x"3500", 989=>x"4b00", 990=>x"4e00", 991=>x"b700", 992=>x"2c00", 993=>x"2700", 994=>x"2900",
---- 995=>x"2900", 996=>x"3400", 997=>x"4200", 998=>x"3f00", 999=>x"ab00", 1000=>x"3700", 1001=>x"2c00",
---- 1002=>x"2d00", 1003=>x"2a00", 1004=>x"3100", 1005=>x"3b00", 1006=>x"4000", 1007=>x"a800", 1008=>x"4000",
---- 1009=>x"3400", 1010=>x"2d00", 1011=>x"2700", 1012=>x"2a00", 1013=>x"3d00", 1014=>x"4000", 1015=>x"a200",
---- 1016=>x"3d00", 1017=>x"4200", 1018=>x"3000", 1019=>x"2c00", 1020=>x"2d00", 1021=>x"4100", 1022=>x"3a00",
---- 1023=>x"9700", 1024=>x"4500", 1025=>x"4000", 1026=>x"2b00", 1027=>x"2700", 1028=>x"2c00", 1029=>x"4500",
---- 1030=>x"3d00", 1031=>x"9500", 1032=>x"4600", 1033=>x"2f00", 1034=>x"2c00", 1035=>x"2700", 1036=>x"2500",
---- 1037=>x"4700", 1038=>x"3900", 1039=>x"8d00", 1040=>x"3900", 1041=>x"2c00", 1042=>x"2d00", 1043=>x"2800",
---- 1044=>x"2900", 1045=>x"4200", 1046=>x"3600", 1047=>x"8600", 1048=>x"2e00", 1049=>x"3100", 1050=>x"3100",
---- 1051=>x"2800", 1052=>x"2c00", 1053=>x"4400", 1054=>x"3400", 1055=>x"8100", 1056=>x"3000", 1057=>x"3000",
---- 1058=>x"3100", 1059=>x"2500", 1060=>x"2b00", 1061=>x"4700", 1062=>x"3000", 1063=>x"7b00", 1064=>x"3100",
---- 1065=>x"2f00", 1066=>x"3200", 1067=>x"2f00", 1068=>x"2e00", 1069=>x"4f00", 1070=>x"2d00", 1071=>x"7a00",
---- 1072=>x"2f00", 1073=>x"2c00", 1074=>x"3100", 1075=>x"2f00", 1076=>x"3100", 1077=>x"5200", 1078=>x"2a00",
---- 1079=>x"7400", 1080=>x"2a00", 1081=>x"2d00", 1082=>x"2800", 1083=>x"2600", 1084=>x"3900", 1085=>x"5600",
---- 1086=>x"2900", 1087=>x"6e00", 1088=>x"cc00", 1089=>x"2c00", 1090=>x"3000", 1091=>x"2d00", 1092=>x"3c00",
---- 1093=>x"5100", 1094=>x"2d00", 1095=>x"6300", 1096=>x"3600", 1097=>x"3000", 1098=>x"3800", 1099=>x"3100",
---- 1100=>x"4000", 1101=>x"5200", 1102=>x"2d00", 1103=>x"6000", 1104=>x"3600", 1105=>x"2d00", 1106=>x"3c00",
---- 1107=>x"3300", 1108=>x"4200", 1109=>x"4a00", 1110=>x"2800", 1111=>x"5b00", 1112=>x"3400", 1113=>x"2900",
---- 1114=>x"3300", 1115=>x"3400", 1116=>x"4b00", 1117=>x"4c00", 1118=>x"2c00", 1119=>x"5800", 1120=>x"2f00",
---- 1121=>x"2900", 1122=>x"3400", 1123=>x"3100", 1124=>x"4800", 1125=>x"b600", 1126=>x"2a00", 1127=>x"5700",
---- 1128=>x"2e00", 1129=>x"2b00", 1130=>x"3400", 1131=>x"3400", 1132=>x"4000", 1133=>x"4600", 1134=>x"2a00",
---- 1135=>x"5400", 1136=>x"3000", 1137=>x"2d00", 1138=>x"3500", 1139=>x"3600", 1140=>x"4200", 1141=>x"4900",
---- 1142=>x"2c00", 1143=>x"5100", 1144=>x"3300", 1145=>x"2e00", 1146=>x"3500", 1147=>x"3c00", 1148=>x"4100",
---- 1149=>x"4100", 1150=>x"2900", 1151=>x"4b00", 1152=>x"3200", 1153=>x"d200", 1154=>x"3700", 1155=>x"3900",
---- 1156=>x"4100", 1157=>x"4400", 1158=>x"2200", 1159=>x"4400", 1160=>x"3300", 1161=>x"3100", 1162=>x"3b00",
---- 1163=>x"3700", 1164=>x"4700", 1165=>x"4200", 1166=>x"2000", 1167=>x"4100", 1168=>x"3200", 1169=>x"3400",
---- 1170=>x"4000", 1171=>x"3900", 1172=>x"4800", 1173=>x"3d00", 1174=>x"2700", 1175=>x"3800", 1176=>x"3200",
---- 1177=>x"3500", 1178=>x"3e00", 1179=>x"3900", 1180=>x"4d00", 1181=>x"3d00", 1182=>x"2600", 1183=>x"3400",
---- 1184=>x"3100", 1185=>x"3700", 1186=>x"3600", 1187=>x"c600", 1188=>x"5500", 1189=>x"3b00", 1190=>x"2700",
---- 1191=>x"3100", 1192=>x"2e00", 1193=>x"3800", 1194=>x"3300", 1195=>x"3b00", 1196=>x"5600", 1197=>x"3600",
---- 1198=>x"2400", 1199=>x"2d00", 1200=>x"2c00", 1201=>x"3600", 1202=>x"3000", 1203=>x"3a00", 1204=>x"5600",
---- 1205=>x"3500", 1206=>x"2400", 1207=>x"2900", 1208=>x"3000", 1209=>x"3300", 1210=>x"3100", 1211=>x"3c00",
---- 1212=>x"5600", 1213=>x"3400", 1214=>x"2600", 1215=>x"2400", 1216=>x"3500", 1217=>x"3600", 1218=>x"3800",
---- 1219=>x"4000", 1220=>x"5700", 1221=>x"3100", 1222=>x"2300", 1223=>x"2200", 1224=>x"3600", 1225=>x"3c00",
---- 1226=>x"3a00", 1227=>x"3d00", 1228=>x"5900", 1229=>x"3600", 1230=>x"2300", 1231=>x"2600", 1232=>x"3200",
---- 1233=>x"3b00", 1234=>x"4300", 1235=>x"4600", 1236=>x"5500", 1237=>x"3800", 1238=>x"2300", 1239=>x"2600",
---- 1240=>x"2f00", 1241=>x"3800", 1242=>x"4200", 1243=>x"4700", 1244=>x"4f00", 1245=>x"3800", 1246=>x"1e00",
---- 1247=>x"2300", 1248=>x"3400", 1249=>x"4000", 1250=>x"4100", 1251=>x"4300", 1252=>x"4e00", 1253=>x"3800",
---- 1254=>x"2200", 1255=>x"2200", 1256=>x"3000", 1257=>x"3b00", 1258=>x"4500", 1259=>x"4a00", 1260=>x"4400",
---- 1261=>x"3d00", 1262=>x"2500", 1263=>x"2400", 1264=>x"2e00", 1265=>x"3c00", 1266=>x"4700", 1267=>x"4a00",
---- 1268=>x"4700", 1269=>x"3800", 1270=>x"2500", 1271=>x"2500", 1272=>x"3200", 1273=>x"3e00", 1274=>x"4500",
---- 1275=>x"4800", 1276=>x"4700", 1277=>x"3500", 1278=>x"2a00", 1279=>x"2700", 1280=>x"3200", 1281=>x"3b00",
---- 1282=>x"4600", 1283=>x"4300", 1284=>x"4700", 1285=>x"3100", 1286=>x"2e00", 1287=>x"2b00", 1288=>x"3600",
---- 1289=>x"3e00", 1290=>x"4a00", 1291=>x"3e00", 1292=>x"ba00", 1293=>x"3200", 1294=>x"3000", 1295=>x"2b00",
---- 1296=>x"3300", 1297=>x"4400", 1298=>x"b600", 1299=>x"3f00", 1300=>x"4a00", 1301=>x"3200", 1302=>x"3100",
---- 1303=>x"3300", 1304=>x"c800", 1305=>x"4500", 1306=>x"4b00", 1307=>x"3c00", 1308=>x"4b00", 1309=>x"3200",
---- 1310=>x"2f00", 1311=>x"3900", 1312=>x"3700", 1313=>x"4b00", 1314=>x"5300", 1315=>x"4000", 1316=>x"4c00",
---- 1317=>x"3100", 1318=>x"2e00", 1319=>x"3300", 1320=>x"3b00", 1321=>x"5100", 1322=>x"5200", 1323=>x"4800",
---- 1324=>x"4800", 1325=>x"3800", 1326=>x"3700", 1327=>x"3500", 1328=>x"3900", 1329=>x"5c00", 1330=>x"4900",
---- 1331=>x"4b00", 1332=>x"4c00", 1333=>x"3400", 1334=>x"4000", 1335=>x"3600", 1336=>x"3900", 1337=>x"5b00",
---- 1338=>x"4900", 1339=>x"4700", 1340=>x"4800", 1341=>x"3900", 1342=>x"3f00", 1343=>x"3900", 1344=>x"3e00",
---- 1345=>x"5b00", 1346=>x"4400", 1347=>x"4600", 1348=>x"4600", 1349=>x"3900", 1350=>x"3e00", 1351=>x"3100",
---- 1352=>x"4200", 1353=>x"5700", 1354=>x"4600", 1355=>x"4600", 1356=>x"4700", 1357=>x"3f00", 1358=>x"3d00",
---- 1359=>x"2f00", 1360=>x"4a00", 1361=>x"5500", 1362=>x"4800", 1363=>x"4800", 1364=>x"3e00", 1365=>x"3d00",
---- 1366=>x"3a00", 1367=>x"3400", 1368=>x"4a00", 1369=>x"5000", 1370=>x"4800", 1371=>x"4800", 1372=>x"3b00",
---- 1373=>x"3c00", 1374=>x"3c00", 1375=>x"3200", 1376=>x"b300", 1377=>x"5300", 1378=>x"4700", 1379=>x"4700",
---- 1380=>x"4b00", 1381=>x"4100", 1382=>x"4300", 1383=>x"3400", 1384=>x"4600", 1385=>x"5500", 1386=>x"4c00",
---- 1387=>x"4b00", 1388=>x"4e00", 1389=>x"3d00", 1390=>x"4400", 1391=>x"3800", 1392=>x"4500", 1393=>x"4d00",
---- 1394=>x"4900", 1395=>x"5200", 1396=>x"4800", 1397=>x"3800", 1398=>x"3e00", 1399=>x"3d00", 1400=>x"4d00",
---- 1401=>x"4800", 1402=>x"4600", 1403=>x"5200", 1404=>x"4700", 1405=>x"2f00", 1406=>x"3e00", 1407=>x"4900",
---- 1408=>x"4f00", 1409=>x"4c00", 1410=>x"4800", 1411=>x"5200", 1412=>x"4500", 1413=>x"2c00", 1414=>x"4000",
---- 1415=>x"5300", 1416=>x"5400", 1417=>x"4800", 1418=>x"4c00", 1419=>x"5200", 1420=>x"4c00", 1421=>x"3400",
---- 1422=>x"3f00", 1423=>x"5800", 1424=>x"5900", 1425=>x"4600", 1426=>x"4b00", 1427=>x"4f00", 1428=>x"3e00",
---- 1429=>x"3300", 1430=>x"4100", 1431=>x"5500", 1432=>x"6000", 1433=>x"4700", 1434=>x"5300", 1435=>x"5400",
---- 1436=>x"4100", 1437=>x"3b00", 1438=>x"4200", 1439=>x"5500", 1440=>x"5d00", 1441=>x"4100", 1442=>x"4f00",
---- 1443=>x"5900", 1444=>x"4200", 1445=>x"4400", 1446=>x"3c00", 1447=>x"5300", 1448=>x"5900", 1449=>x"3f00",
---- 1450=>x"5000", 1451=>x"5400", 1452=>x"4900", 1453=>x"4300", 1454=>x"3600", 1455=>x"5a00", 1456=>x"5700",
---- 1457=>x"4600", 1458=>x"5000", 1459=>x"5300", 1460=>x"4800", 1461=>x"3f00", 1462=>x"3800", 1463=>x"5400",
---- 1464=>x"5e00", 1465=>x"4400", 1466=>x"5000", 1467=>x"5d00", 1468=>x"4700", 1469=>x"3f00", 1470=>x"3f00",
---- 1471=>x"5100", 1472=>x"5e00", 1473=>x"4900", 1474=>x"5000", 1475=>x"5900", 1476=>x"4500", 1477=>x"4000",
---- 1478=>x"3c00", 1479=>x"5000", 1480=>x"6100", 1481=>x"4400", 1482=>x"4e00", 1483=>x"5700", 1484=>x"4b00",
---- 1485=>x"4600", 1486=>x"4500", 1487=>x"5000", 1488=>x"6200", 1489=>x"4600", 1490=>x"5400", 1491=>x"5400",
---- 1492=>x"4b00", 1493=>x"4600", 1494=>x"4a00", 1495=>x"5300", 1496=>x"6200", 1497=>x"4900", 1498=>x"5700",
---- 1499=>x"5c00", 1500=>x"4a00", 1501=>x"4100", 1502=>x"4b00", 1503=>x"5200", 1504=>x"6800", 1505=>x"4a00",
---- 1506=>x"5500", 1507=>x"5b00", 1508=>x"4800", 1509=>x"4600", 1510=>x"4a00", 1511=>x"4b00", 1512=>x"6900",
---- 1513=>x"4900", 1514=>x"5900", 1515=>x"5800", 1516=>x"4800", 1517=>x"4d00", 1518=>x"af00", 1519=>x"4c00",
---- 1520=>x"6300", 1521=>x"4700", 1522=>x"5900", 1523=>x"5400", 1524=>x"4400", 1525=>x"4e00", 1526=>x"4f00",
---- 1527=>x"4b00", 1528=>x"6400", 1529=>x"5000", 1530=>x"5700", 1531=>x"5500", 1532=>x"4b00", 1533=>x"ae00",
---- 1534=>x"5400", 1535=>x"5200", 1536=>x"6500", 1537=>x"5300", 1538=>x"5600", 1539=>x"5700", 1540=>x"4c00",
---- 1541=>x"5400", 1542=>x"5900", 1543=>x"aa00", 1544=>x"6800", 1545=>x"5400", 1546=>x"5a00", 1547=>x"5700",
---- 1548=>x"4d00", 1549=>x"5000", 1550=>x"5500", 1551=>x"5800", 1552=>x"6800", 1553=>x"5100", 1554=>x"5c00",
---- 1555=>x"5900", 1556=>x"4e00", 1557=>x"af00", 1558=>x"5700", 1559=>x"5200", 1560=>x"6a00", 1561=>x"4f00",
---- 1562=>x"5a00", 1563=>x"5a00", 1564=>x"4e00", 1565=>x"4f00", 1566=>x"5600", 1567=>x"5a00", 1568=>x"6a00",
---- 1569=>x"4e00", 1570=>x"5600", 1571=>x"5800", 1572=>x"5400", 1573=>x"4c00", 1574=>x"5000", 1575=>x"5900",
---- 1576=>x"6b00", 1577=>x"4f00", 1578=>x"5300", 1579=>x"5900", 1580=>x"4f00", 1581=>x"4e00", 1582=>x"5400",
---- 1583=>x"5900", 1584=>x"6900", 1585=>x"4e00", 1586=>x"5100", 1587=>x"5400", 1588=>x"4c00", 1589=>x"4900",
---- 1590=>x"5300", 1591=>x"5700", 1592=>x"6600", 1593=>x"4b00", 1594=>x"4f00", 1595=>x"5500", 1596=>x"4f00",
---- 1597=>x"4c00", 1598=>x"5000", 1599=>x"5000", 1600=>x"9b00", 1601=>x"4d00", 1602=>x"4d00", 1603=>x"5200",
---- 1604=>x"4e00", 1605=>x"4600", 1606=>x"4d00", 1607=>x"b400", 1608=>x"6500", 1609=>x"4b00", 1610=>x"4800",
---- 1611=>x"4e00", 1612=>x"4900", 1613=>x"4300", 1614=>x"4b00", 1615=>x"4a00", 1616=>x"6600", 1617=>x"4a00",
---- 1618=>x"4600", 1619=>x"4e00", 1620=>x"4800", 1621=>x"4900", 1622=>x"5200", 1623=>x"4a00", 1624=>x"5d00",
---- 1625=>x"4600", 1626=>x"4100", 1627=>x"4800", 1628=>x"4200", 1629=>x"4200", 1630=>x"4e00", 1631=>x"4900",
---- 1632=>x"5300", 1633=>x"4000", 1634=>x"3700", 1635=>x"4400", 1636=>x"3b00", 1637=>x"4400", 1638=>x"4e00",
---- 1639=>x"4500", 1640=>x"af00", 1641=>x"4500", 1642=>x"3b00", 1643=>x"3d00", 1644=>x"3e00", 1645=>x"4d00",
---- 1646=>x"4f00", 1647=>x"4700", 1648=>x"3800", 1649=>x"4000", 1650=>x"3000", 1651=>x"3800", 1652=>x"3700",
---- 1653=>x"4900", 1654=>x"4700", 1655=>x"4600", 1656=>x"3400", 1657=>x"3400", 1658=>x"2c00", 1659=>x"2f00",
---- 1660=>x"3600", 1661=>x"4900", 1662=>x"3f00", 1663=>x"4400", 1664=>x"7d00", 1665=>x"3300", 1666=>x"2d00",
---- 1667=>x"2b00", 1668=>x"3400", 1669=>x"4400", 1670=>x"3a00", 1671=>x"3e00", 1672=>x"ca00", 1673=>x"5d00",
---- 1674=>x"2b00", 1675=>x"2d00", 1676=>x"3200", 1677=>x"3c00", 1678=>x"3200", 1679=>x"3b00", 1680=>x"df00",
---- 1681=>x"aa00", 1682=>x"3400", 1683=>x"2500", 1684=>x"3000", 1685=>x"4200", 1686=>x"2e00", 1687=>x"3700",
---- 1688=>x"dd00", 1689=>x"d900", 1690=>x"6c00", 1691=>x"2300", 1692=>x"2c00", 1693=>x"3d00", 1694=>x"2c00",
---- 1695=>x"3600", 1696=>x"db00", 1697=>x"e200", 1698=>x"b300", 1699=>x"3500", 1700=>x"2700", 1701=>x"2f00",
---- 1702=>x"2c00", 1703=>x"2e00", 1704=>x"dc00", 1705=>x"dc00", 1706=>x"db00", 1707=>x"6700", 1708=>x"2100",
---- 1709=>x"3100", 1710=>x"2800", 1711=>x"2a00", 1712=>x"dc00", 1713=>x"dd00", 1714=>x"e300", 1715=>x"a700",
---- 1716=>x"2a00", 1717=>x"2500", 1718=>x"2300", 1719=>x"2800", 1720=>x"db00", 1721=>x"dd00", 1722=>x"df00",
---- 1723=>x"d500", 1724=>x"5400", 1725=>x"1f00", 1726=>x"2700", 1727=>x"2500", 1728=>x"d800", 1729=>x"dd00",
---- 1730=>x"dc00", 1731=>x"e200", 1732=>x"9000", 1733=>x"2700", 1734=>x"2400", 1735=>x"2400", 1736=>x"d700",
---- 1737=>x"db00", 1738=>x"dd00", 1739=>x"e200", 1740=>x"be00", 1741=>x"3100", 1742=>x"1800", 1743=>x"2100",
---- 1744=>x"d800", 1745=>x"da00", 1746=>x"dc00", 1747=>x"de00", 1748=>x"d800", 1749=>x"5a00", 1750=>x"1800",
---- 1751=>x"df00", 1752=>x"d700", 1753=>x"d800", 1754=>x"da00", 1755=>x"dc00", 1756=>x"e000", 1757=>x"8b00",
---- 1758=>x"1900", 1759=>x"1f00", 1760=>x"d500", 1761=>x"d700", 1762=>x"da00", 1763=>x"da00", 1764=>x"e100",
---- 1765=>x"b600", 1766=>x"2800", 1767=>x"1a00", 1768=>x"d700", 1769=>x"d800", 1770=>x"d800", 1771=>x"da00",
---- 1772=>x"de00", 1773=>x"d000", 1774=>x"4b00", 1775=>x"1500", 1776=>x"d500", 1777=>x"d700", 1778=>x"d800",
---- 1779=>x"d900", 1780=>x"d900", 1781=>x"dd00", 1782=>x"7500", 1783=>x"1600", 1784=>x"d300", 1785=>x"d600",
---- 1786=>x"d600", 1787=>x"da00", 1788=>x"d600", 1789=>x"df00", 1790=>x"a000", 1791=>x"1a00", 1792=>x"d500",
---- 1793=>x"d500", 1794=>x"d600", 1795=>x"d600", 1796=>x"d600", 1797=>x"dc00", 1798=>x"c000", 1799=>x"2d00",
---- 1800=>x"d500", 1801=>x"d400", 1802=>x"d700", 1803=>x"d500", 1804=>x"d700", 1805=>x"d900", 1806=>x"d500",
---- 1807=>x"4f00", 1808=>x"d200", 1809=>x"d600", 1810=>x"d500", 1811=>x"d600", 1812=>x"d600", 1813=>x"d500",
---- 1814=>x"dd00", 1815=>x"8200", 1816=>x"d200", 1817=>x"d400", 1818=>x"d400", 1819=>x"d400", 1820=>x"d500",
---- 1821=>x"d500", 1822=>x"dc00", 1823=>x"ae00", 1824=>x"d600", 1825=>x"d300", 1826=>x"d500", 1827=>x"d300",
---- 1828=>x"d500", 1829=>x"d500", 1830=>x"d800", 1831=>x"c900", 1832=>x"d200", 1833=>x"d400", 1834=>x"d500",
---- 1835=>x"d600", 1836=>x"d500", 1837=>x"d500", 1838=>x"d600", 1839=>x"d900", 1840=>x"d300", 1841=>x"d300",
---- 1842=>x"d400", 1843=>x"d600", 1844=>x"d600", 1845=>x"d400", 1846=>x"d600", 1847=>x"dc00", 1848=>x"d200",
---- 1849=>x"d500", 1850=>x"d600", 1851=>x"d600", 1852=>x"d600", 1853=>x"d600", 1854=>x"d700", 1855=>x"dc00",
---- 1856=>x"d200", 1857=>x"d500", 1858=>x"2b00", 1859=>x"d500", 1860=>x"d600", 1861=>x"d800", 1862=>x"da00",
---- 1863=>x"db00", 1864=>x"d100", 1865=>x"d400", 1866=>x"d500", 1867=>x"d400", 1868=>x"d500", 1869=>x"d700",
---- 1870=>x"d900", 1871=>x"d900", 1872=>x"d100", 1873=>x"d300", 1874=>x"d300", 1875=>x"d300", 1876=>x"d500",
---- 1877=>x"d700", 1878=>x"d900", 1879=>x"d800", 1880=>x"d000", 1881=>x"d100", 1882=>x"d200", 1883=>x"d400",
---- 1884=>x"d400", 1885=>x"d500", 1886=>x"d800", 1887=>x"d900", 1888=>x"ce00", 1889=>x"d000", 1890=>x"d100",
---- 1891=>x"d400", 1892=>x"d500", 1893=>x"d600", 1894=>x"d900", 1895=>x"d800", 1896=>x"d000", 1897=>x"d100",
---- 1898=>x"d000", 1899=>x"d300", 1900=>x"d500", 1901=>x"d500", 1902=>x"d700", 1903=>x"d800", 1904=>x"3100",
---- 1905=>x"d000", 1906=>x"d200", 1907=>x"d300", 1908=>x"d100", 1909=>x"d400", 1910=>x"d600", 1911=>x"d700",
---- 1912=>x"cd00", 1913=>x"ce00", 1914=>x"d000", 1915=>x"d100", 1916=>x"d100", 1917=>x"d400", 1918=>x"d500",
---- 1919=>x"2800", 1920=>x"ce00", 1921=>x"d100", 1922=>x"cf00", 1923=>x"d000", 1924=>x"d100", 1925=>x"d400",
---- 1926=>x"d600", 1927=>x"d300", 1928=>x"cc00", 1929=>x"ce00", 1930=>x"ce00", 1931=>x"d100", 1932=>x"d300",
---- 1933=>x"d400", 1934=>x"d400", 1935=>x"d300", 1936=>x"c900", 1937=>x"cc00", 1938=>x"cf00", 1939=>x"d000",
---- 1940=>x"d200", 1941=>x"d100", 1942=>x"d500", 1943=>x"d400", 1944=>x"c800", 1945=>x"cb00", 1946=>x"cd00",
---- 1947=>x"ce00", 1948=>x"d200", 1949=>x"d300", 1950=>x"d500", 1951=>x"d400", 1952=>x"c800", 1953=>x"c800",
---- 1954=>x"cd00", 1955=>x"ce00", 1956=>x"d100", 1957=>x"d300", 1958=>x"d500", 1959=>x"d400", 1960=>x"c700",
---- 1961=>x"c900", 1962=>x"cc00", 1963=>x"cc00", 1964=>x"d100", 1965=>x"d000", 1966=>x"d200", 1967=>x"d200",
---- 1968=>x"c400", 1969=>x"c800", 1970=>x"cb00", 1971=>x"ce00", 1972=>x"cf00", 1973=>x"d000", 1974=>x"d300",
---- 1975=>x"d400", 1976=>x"c300", 1977=>x"c500", 1978=>x"c900", 1979=>x"cb00", 1980=>x"cd00", 1981=>x"cf00",
---- 1982=>x"d300", 1983=>x"d500", 1984=>x"c000", 1985=>x"c400", 1986=>x"c600", 1987=>x"c800", 1988=>x"cc00",
---- 1989=>x"cd00", 1990=>x"d200", 1991=>x"d400", 1992=>x"bd00", 1993=>x"c300", 1994=>x"c300", 1995=>x"c500",
---- 1996=>x"ca00", 1997=>x"cb00", 1998=>x"d100", 1999=>x"d300", 2000=>x"bb00", 2001=>x"c100", 2002=>x"c500",
---- 2003=>x"c700", 2004=>x"ca00", 2005=>x"cb00", 2006=>x"ce00", 2007=>x"d100", 2008=>x"ba00", 2009=>x"bd00",
---- 2010=>x"c600", 2011=>x"c700", 2012=>x"c900", 2013=>x"cb00", 2014=>x"cd00", 2015=>x"cd00", 2016=>x"bc00",
---- 2017=>x"bd00", 2018=>x"c400", 2019=>x"c500", 2020=>x"c900", 2021=>x"ca00", 2022=>x"cd00", 2023=>x"ce00",
---- 2024=>x"b800", 2025=>x"bc00", 2026=>x"c100", 2027=>x"c300", 2028=>x"c700", 2029=>x"c900", 2030=>x"cb00",
---- 2031=>x"ce00", 2032=>x"bb00", 2033=>x"bf00", 2034=>x"c100", 2035=>x"c400", 2036=>x"c500", 2037=>x"c800",
---- 2038=>x"ca00", 2039=>x"cc00", 2040=>x"b900", 2041=>x"bf00", 2042=>x"c000", 2043=>x"c200", 2044=>x"c200",
---- 2045=>x"c500", 2046=>x"c800", 2047=>x"ca00"),
---- 23 => (0=>x"9a00", 1=>x"9800", 2=>x"9a00", 3=>x"9900", 4=>x"9800", 5=>x"9900", 6=>x"9c00", 7=>x"9900",
---- 8=>x"9a00", 9=>x"9800", 10=>x"9a00", 11=>x"9900", 12=>x"9800", 13=>x"9900", 14=>x"9c00",
---- 15=>x"9800", 16=>x"9900", 17=>x"9900", 18=>x"9900", 19=>x"9900", 20=>x"9800", 21=>x"9900",
---- 22=>x"9d00", 23=>x"9a00", 24=>x"9900", 25=>x"9800", 26=>x"9700", 27=>x"9a00", 28=>x"9c00",
---- 29=>x"9a00", 30=>x"9b00", 31=>x"9800", 32=>x"9c00", 33=>x"9c00", 34=>x"6400", 35=>x"9800",
---- 36=>x"9a00", 37=>x"9900", 38=>x"9900", 39=>x"9900", 40=>x"9d00", 41=>x"9d00", 42=>x"9a00",
---- 43=>x"9b00", 44=>x"9a00", 45=>x"9d00", 46=>x"9b00", 47=>x"6600", 48=>x"9d00", 49=>x"9c00",
---- 50=>x"9c00", 51=>x"9b00", 52=>x"9c00", 53=>x"9c00", 54=>x"9b00", 55=>x"9900", 56=>x"9d00",
---- 57=>x"9c00", 58=>x"9c00", 59=>x"9b00", 60=>x"9d00", 61=>x"9b00", 62=>x"9800", 63=>x"9a00",
---- 64=>x"9e00", 65=>x"9e00", 66=>x"9e00", 67=>x"9e00", 68=>x"9d00", 69=>x"9a00", 70=>x"9900",
---- 71=>x"9a00", 72=>x"9f00", 73=>x"9e00", 74=>x"9e00", 75=>x"a000", 76=>x"9f00", 77=>x"9d00",
---- 78=>x"9b00", 79=>x"9a00", 80=>x"a000", 81=>x"9d00", 82=>x"9c00", 83=>x"9f00", 84=>x"9e00",
---- 85=>x"9f00", 86=>x"9a00", 87=>x"9c00", 88=>x"a100", 89=>x"a100", 90=>x"9c00", 91=>x"9a00",
---- 92=>x"9d00", 93=>x"9b00", 94=>x"9b00", 95=>x"9b00", 96=>x"a100", 97=>x"a100", 98=>x"9e00",
---- 99=>x"9a00", 100=>x"9b00", 101=>x"9d00", 102=>x"9c00", 103=>x"9b00", 104=>x"9e00", 105=>x"9f00",
---- 106=>x"a000", 107=>x"9b00", 108=>x"9c00", 109=>x"9e00", 110=>x"9b00", 111=>x"9b00", 112=>x"9f00",
---- 113=>x"9f00", 114=>x"9e00", 115=>x"9c00", 116=>x"9d00", 117=>x"9b00", 118=>x"9c00", 119=>x"9e00",
---- 120=>x"9e00", 121=>x"9e00", 122=>x"9d00", 123=>x"9e00", 124=>x"9e00", 125=>x"9b00", 126=>x"9a00",
---- 127=>x"9c00", 128=>x"9d00", 129=>x"9e00", 130=>x"9e00", 131=>x"9a00", 132=>x"9d00", 133=>x"9b00",
---- 134=>x"9d00", 135=>x"9c00", 136=>x"9f00", 137=>x"9d00", 138=>x"9e00", 139=>x"9c00", 140=>x"9d00",
---- 141=>x"9d00", 142=>x"9c00", 143=>x"9c00", 144=>x"9f00", 145=>x"9b00", 146=>x"9b00", 147=>x"9a00",
---- 148=>x"a000", 149=>x"9e00", 150=>x"9a00", 151=>x"9f00", 152=>x"9d00", 153=>x"9e00", 154=>x"9b00",
---- 155=>x"9b00", 156=>x"9d00", 157=>x"9d00", 158=>x"9900", 159=>x"9900", 160=>x"9c00", 161=>x"9b00",
---- 162=>x"9b00", 163=>x"9b00", 164=>x"9b00", 165=>x"9a00", 166=>x"9800", 167=>x"9800", 168=>x"9900",
---- 169=>x"9b00", 170=>x"9b00", 171=>x"9a00", 172=>x"9b00", 173=>x"9900", 174=>x"9900", 175=>x"9a00",
---- 176=>x"9a00", 177=>x"9b00", 178=>x"9a00", 179=>x"9a00", 180=>x"9b00", 181=>x"9900", 182=>x"9b00",
---- 183=>x"9c00", 184=>x"9900", 185=>x"9900", 186=>x"9900", 187=>x"9900", 188=>x"9a00", 189=>x"9a00",
---- 190=>x"9b00", 191=>x"9a00", 192=>x"9800", 193=>x"9700", 194=>x"9900", 195=>x"9a00", 196=>x"6600",
---- 197=>x"6600", 198=>x"9c00", 199=>x"9a00", 200=>x"9800", 201=>x"9900", 202=>x"9a00", 203=>x"9900",
---- 204=>x"9900", 205=>x"9900", 206=>x"9a00", 207=>x"9900", 208=>x"9900", 209=>x"9900", 210=>x"9800",
---- 211=>x"9700", 212=>x"9a00", 213=>x"9800", 214=>x"9700", 215=>x"9800", 216=>x"9a00", 217=>x"9800",
---- 218=>x"9500", 219=>x"9600", 220=>x"9800", 221=>x"9700", 222=>x"9400", 223=>x"9200", 224=>x"9800",
---- 225=>x"9800", 226=>x"9600", 227=>x"9400", 228=>x"9600", 229=>x"9600", 230=>x"9300", 231=>x"9300",
---- 232=>x"9600", 233=>x"9a00", 234=>x"9600", 235=>x"9200", 236=>x"6c00", 237=>x"9200", 238=>x"9400",
---- 239=>x"9300", 240=>x"9700", 241=>x"9800", 242=>x"9800", 243=>x"9500", 244=>x"9300", 245=>x"8e00",
---- 246=>x"9200", 247=>x"9100", 248=>x"9500", 249=>x"9600", 250=>x"9900", 251=>x"9800", 252=>x"9500",
---- 253=>x"9200", 254=>x"9000", 255=>x"8d00", 256=>x"9300", 257=>x"9400", 258=>x"9800", 259=>x"9800",
---- 260=>x"9500", 261=>x"9200", 262=>x"8e00", 263=>x"8e00", 264=>x"9000", 265=>x"9200", 266=>x"9600",
---- 267=>x"9600", 268=>x"9700", 269=>x"9000", 270=>x"8e00", 271=>x"8b00", 272=>x"8d00", 273=>x"8e00",
---- 274=>x"9000", 275=>x"9500", 276=>x"9900", 277=>x"9200", 278=>x"8f00", 279=>x"8f00", 280=>x"7600",
---- 281=>x"8b00", 282=>x"8d00", 283=>x"9300", 284=>x"9600", 285=>x"9400", 286=>x"9100", 287=>x"9100",
---- 288=>x"8200", 289=>x"8500", 290=>x"8800", 291=>x"8d00", 292=>x"9500", 293=>x"9600", 294=>x"9300",
---- 295=>x"6e00", 296=>x"7c00", 297=>x"7f00", 298=>x"8300", 299=>x"8a00", 300=>x"9200", 301=>x"9700",
---- 302=>x"9500", 303=>x"9100", 304=>x"7400", 305=>x"7800", 306=>x"8000", 307=>x"8700", 308=>x"8e00",
---- 309=>x"9300", 310=>x"9600", 311=>x"6c00", 312=>x"6b00", 313=>x"6e00", 314=>x"7500", 315=>x"7f00",
---- 316=>x"8b00", 317=>x"8f00", 318=>x"9400", 319=>x"9500", 320=>x"5f00", 321=>x"5f00", 322=>x"6900",
---- 323=>x"7800", 324=>x"8300", 325=>x"8a00", 326=>x"9200", 327=>x"9700", 328=>x"5500", 329=>x"5400",
---- 330=>x"5900", 331=>x"6900", 332=>x"7b00", 333=>x"8800", 334=>x"8e00", 335=>x"9300", 336=>x"4d00",
---- 337=>x"4400", 338=>x"4900", 339=>x"5e00", 340=>x"7300", 341=>x"8200", 342=>x"8800", 343=>x"9000",
---- 344=>x"4100", 345=>x"3700", 346=>x"3900", 347=>x"5300", 348=>x"6b00", 349=>x"7b00", 350=>x"8500",
---- 351=>x"8a00", 352=>x"4700", 353=>x"3400", 354=>x"3200", 355=>x"4300", 356=>x"a500", 357=>x"7100",
---- 358=>x"7d00", 359=>x"8800", 360=>x"4c00", 361=>x"3000", 362=>x"2a00", 363=>x"3500", 364=>x"4e00",
---- 365=>x"6600", 366=>x"7300", 367=>x"7f00", 368=>x"4c00", 369=>x"2f00", 370=>x"2900", 371=>x"2e00",
---- 372=>x"4500", 373=>x"6000", 374=>x"6b00", 375=>x"7800", 376=>x"4c00", 377=>x"2f00", 378=>x"2400",
---- 379=>x"2c00", 380=>x"3b00", 381=>x"5600", 382=>x"6800", 383=>x"7400", 384=>x"4a00", 385=>x"2e00",
---- 386=>x"2b00", 387=>x"3100", 388=>x"3400", 389=>x"4d00", 390=>x"6100", 391=>x"6b00", 392=>x"4c00",
---- 393=>x"3100", 394=>x"2900", 395=>x"2e00", 396=>x"3700", 397=>x"3400", 398=>x"4e00", 399=>x"6100",
---- 400=>x"4f00", 401=>x"3300", 402=>x"2d00", 403=>x"2a00", 404=>x"2700", 405=>x"2d00", 406=>x"3b00",
---- 407=>x"5200", 408=>x"4e00", 409=>x"3600", 410=>x"3100", 411=>x"2c00", 412=>x"2500", 413=>x"2d00",
---- 414=>x"3100", 415=>x"4600", 416=>x"5200", 417=>x"3500", 418=>x"2d00", 419=>x"2a00", 420=>x"2800",
---- 421=>x"2900", 422=>x"2b00", 423=>x"3600", 424=>x"5300", 425=>x"3800", 426=>x"2c00", 427=>x"2c00",
---- 428=>x"2f00", 429=>x"2900", 430=>x"2900", 431=>x"2c00", 432=>x"5000", 433=>x"3a00", 434=>x"2e00",
---- 435=>x"2d00", 436=>x"2d00", 437=>x"2b00", 438=>x"2800", 439=>x"2700", 440=>x"5300", 441=>x"3c00",
---- 442=>x"3000", 443=>x"2d00", 444=>x"2e00", 445=>x"2d00", 446=>x"2900", 447=>x"2800", 448=>x"5200",
---- 449=>x"c200", 450=>x"3000", 451=>x"2c00", 452=>x"2c00", 453=>x"2e00", 454=>x"2b00", 455=>x"2a00",
---- 456=>x"5100", 457=>x"3900", 458=>x"2f00", 459=>x"2b00", 460=>x"2f00", 461=>x"2c00", 462=>x"2c00",
---- 463=>x"2700", 464=>x"5500", 465=>x"3900", 466=>x"2e00", 467=>x"2d00", 468=>x"2e00", 469=>x"2b00",
---- 470=>x"2700", 471=>x"2600", 472=>x"5100", 473=>x"3900", 474=>x"2c00", 475=>x"2900", 476=>x"2a00",
---- 477=>x"2600", 478=>x"2600", 479=>x"2400", 480=>x"5100", 481=>x"3500", 482=>x"2c00", 483=>x"2800",
---- 484=>x"2800", 485=>x"2700", 486=>x"2100", 487=>x"3300", 488=>x"4a00", 489=>x"2e00", 490=>x"2800",
---- 491=>x"2500", 492=>x"2400", 493=>x"2200", 494=>x"4600", 495=>x"a200", 496=>x"4200", 497=>x"2900",
---- 498=>x"db00", 499=>x"2200", 500=>x"2300", 501=>x"5c00", 502=>x"b700", 503=>x"d900", 504=>x"3f00",
---- 505=>x"2700", 506=>x"1e00", 507=>x"d300", 508=>x"7300", 509=>x"c800", 510=>x"de00", 511=>x"d100",
---- 512=>x"3200", 513=>x"2500", 514=>x"4500", 515=>x"9300", 516=>x"d500", 517=>x"db00", 518=>x"ce00",
---- 519=>x"a900", 520=>x"3d00", 521=>x"7300", 522=>x"ba00", 523=>x"dc00", 524=>x"d200", 525=>x"c000",
---- 526=>x"ac00", 527=>x"b600", 528=>x"9e00", 529=>x"d700", 530=>x"d700", 531=>x"c800", 532=>x"b900",
---- 533=>x"ad00", 534=>x"bc00", 535=>x"d400", 536=>x"de00", 537=>x"cf00", 538=>x"be00", 539=>x"b900",
---- 540=>x"b900", 541=>x"c400", 542=>x"d300", 543=>x"d500", 544=>x"c500", 545=>x"bc00", 546=>x"b800",
---- 547=>x"bc00", 548=>x"c900", 549=>x"d300", 550=>x"d500", 551=>x"d200", 552=>x"bd00", 553=>x"b600",
---- 554=>x"be00", 555=>x"cc00", 556=>x"d400", 557=>x"d300", 558=>x"d000", 559=>x"cf00", 560=>x"b900",
---- 561=>x"c800", 562=>x"d400", 563=>x"d300", 564=>x"d100", 565=>x"ce00", 566=>x"cb00", 567=>x"ca00",
---- 568=>x"cd00", 569=>x"d500", 570=>x"d100", 571=>x"ce00", 572=>x"cc00", 573=>x"c800", 574=>x"c700",
---- 575=>x"c900", 576=>x"d300", 577=>x"d000", 578=>x"cc00", 579=>x"cc00", 580=>x"c800", 581=>x"c800",
---- 582=>x"c900", 583=>x"c900", 584=>x"cd00", 585=>x"cc00", 586=>x"ca00", 587=>x"c900", 588=>x"c900",
---- 589=>x"c700", 590=>x"c500", 591=>x"c800", 592=>x"c900", 593=>x"ca00", 594=>x"c900", 595=>x"c800",
---- 596=>x"ca00", 597=>x"c600", 598=>x"c600", 599=>x"c900", 600=>x"c800", 601=>x"c800", 602=>x"c800",
---- 603=>x"c900", 604=>x"c600", 605=>x"c600", 606=>x"3800", 607=>x"ca00", 608=>x"c800", 609=>x"c900",
---- 610=>x"c700", 611=>x"c700", 612=>x"c500", 613=>x"c600", 614=>x"c900", 615=>x"cc00", 616=>x"c800",
---- 617=>x"c800", 618=>x"c600", 619=>x"c700", 620=>x"c900", 621=>x"c900", 622=>x"cb00", 623=>x"cc00",
---- 624=>x"c800", 625=>x"c700", 626=>x"c600", 627=>x"c900", 628=>x"ca00", 629=>x"c900", 630=>x"cb00",
---- 631=>x"3200", 632=>x"c700", 633=>x"c900", 634=>x"c500", 635=>x"c900", 636=>x"ca00", 637=>x"ca00",
---- 638=>x"cc00", 639=>x"cc00", 640=>x"c900", 641=>x"ca00", 642=>x"c800", 643=>x"cb00", 644=>x"c700",
---- 645=>x"cd00", 646=>x"cf00", 647=>x"ce00", 648=>x"c800", 649=>x"c700", 650=>x"ca00", 651=>x"ca00",
---- 652=>x"ca00", 653=>x"3100", 654=>x"d000", 655=>x"cf00", 656=>x"c800", 657=>x"cb00", 658=>x"cb00",
---- 659=>x"cb00", 660=>x"cd00", 661=>x"ce00", 662=>x"d100", 663=>x"d200", 664=>x"ca00", 665=>x"ca00",
---- 666=>x"cb00", 667=>x"cc00", 668=>x"d000", 669=>x"d200", 670=>x"d100", 671=>x"d300", 672=>x"c900",
---- 673=>x"cb00", 674=>x"3400", 675=>x"ce00", 676=>x"d100", 677=>x"d100", 678=>x"d500", 679=>x"ca00",
---- 680=>x"ca00", 681=>x"cd00", 682=>x"cc00", 683=>x"d000", 684=>x"d300", 685=>x"d100", 686=>x"d600",
---- 687=>x"ac00", 688=>x"c900", 689=>x"ce00", 690=>x"cd00", 691=>x"d100", 692=>x"d300", 693=>x"d600",
---- 694=>x"c200", 695=>x"9b00", 696=>x"cc00", 697=>x"cf00", 698=>x"d000", 699=>x"d200", 700=>x"d900",
---- 701=>x"cb00", 702=>x"a900", 703=>x"a600", 704=>x"cc00", 705=>x"ce00", 706=>x"d300", 707=>x"d500",
---- 708=>x"c900", 709=>x"af00", 710=>x"9700", 711=>x"8400", 712=>x"ce00", 713=>x"d300", 714=>x"ce00",
---- 715=>x"b800", 716=>x"9a00", 717=>x"7e00", 718=>x"6500", 719=>x"5000", 720=>x"ca00", 721=>x"ad00",
---- 722=>x"8800", 723=>x"6e00", 724=>x"6200", 725=>x"5b00", 726=>x"5600", 727=>x"5500", 728=>x"7700",
---- 729=>x"5d00", 730=>x"5500", 731=>x"5500", 732=>x"5b00", 733=>x"5d00", 734=>x"5b00", 735=>x"5800",
---- 736=>x"5300", 737=>x"5600", 738=>x"5600", 739=>x"5900", 740=>x"9f00", 741=>x"5a00", 742=>x"5c00",
---- 743=>x"6000", 744=>x"5c00", 745=>x"5a00", 746=>x"5600", 747=>x"5900", 748=>x"6000", 749=>x"6600",
---- 750=>x"6e00", 751=>x"7900", 752=>x"5900", 753=>x"5700", 754=>x"5800", 755=>x"5f00", 756=>x"7200",
---- 757=>x"8300", 758=>x"9500", 759=>x"9d00", 760=>x"5b00", 761=>x"6900", 762=>x"7500", 763=>x"8700",
---- 764=>x"9b00", 765=>x"9f00", 766=>x"a800", 767=>x"aa00", 768=>x"8800", 769=>x"9b00", 770=>x"a300",
---- 771=>x"a800", 772=>x"a900", 773=>x"a500", 774=>x"a500", 775=>x"ad00", 776=>x"a700", 777=>x"a700",
---- 778=>x"a700", 779=>x"a600", 780=>x"aa00", 781=>x"a800", 782=>x"a800", 783=>x"b200", 784=>x"a600",
---- 785=>x"a700", 786=>x"a600", 787=>x"a600", 788=>x"a900", 789=>x"b000", 790=>x"b700", 791=>x"c900",
---- 792=>x"aa00", 793=>x"aa00", 794=>x"aa00", 795=>x"ac00", 796=>x"b200", 797=>x"b900", 798=>x"c900",
---- 799=>x"d500", 800=>x"ab00", 801=>x"ac00", 802=>x"b000", 803=>x"b100", 804=>x"b900", 805=>x"ce00",
---- 806=>x"b600", 807=>x"6900", 808=>x"a700", 809=>x"ac00", 810=>x"ae00", 811=>x"be00", 812=>x"d000",
---- 813=>x"a300", 814=>x"3f00", 815=>x"2100", 816=>x"ae00", 817=>x"b500", 818=>x"c300", 819=>x"ce00",
---- 820=>x"8a00", 821=>x"3300", 822=>x"2500", 823=>x"2f00", 824=>x"c000", 825=>x"ce00", 826=>x"4900",
---- 827=>x"7100", 828=>x"2e00", 829=>x"2a00", 830=>x"2a00", 831=>x"2c00", 832=>x"bd00", 833=>x"9100",
---- 834=>x"4b00", 835=>x"2a00", 836=>x"2b00", 837=>x"2f00", 838=>x"2d00", 839=>x"2d00", 840=>x"8300",
---- 841=>x"5000", 842=>x"2800", 843=>x"2c00", 844=>x"2900", 845=>x"2e00", 846=>x"2c00", 847=>x"3100",
---- 848=>x"7400", 849=>x"5800", 850=>x"2b00", 851=>x"2500", 852=>x"2c00", 853=>x"2e00", 854=>x"2a00",
---- 855=>x"2c00", 856=>x"7600", 857=>x"4a00", 858=>x"2f00", 859=>x"2900", 860=>x"2900", 861=>x"2600",
---- 862=>x"2c00", 863=>x"2e00", 864=>x"7600", 865=>x"3e00", 866=>x"2c00", 867=>x"2b00", 868=>x"2a00",
---- 869=>x"2a00", 870=>x"2f00", 871=>x"2e00", 872=>x"6400", 873=>x"3500", 874=>x"3400", 875=>x"3000",
---- 876=>x"3000", 877=>x"3000", 878=>x"2e00", 879=>x"2f00", 880=>x"5500", 881=>x"2e00", 882=>x"3200",
---- 883=>x"2f00", 884=>x"2c00", 885=>x"2d00", 886=>x"2f00", 887=>x"3100", 888=>x"4d00", 889=>x"2a00",
---- 890=>x"3000", 891=>x"2b00", 892=>x"2d00", 893=>x"3000", 894=>x"2e00", 895=>x"3300", 896=>x"4e00",
---- 897=>x"2d00", 898=>x"3400", 899=>x"2f00", 900=>x"3400", 901=>x"3800", 902=>x"3600", 903=>x"3700",
---- 904=>x"5f00", 905=>x"3400", 906=>x"3c00", 907=>x"3000", 908=>x"3100", 909=>x"3200", 910=>x"3400",
---- 911=>x"3800", 912=>x"6a00", 913=>x"3500", 914=>x"3200", 915=>x"3900", 916=>x"3000", 917=>x"3300",
---- 918=>x"3300", 919=>x"3700", 920=>x"6600", 921=>x"3e00", 922=>x"3300", 923=>x"3800", 924=>x"3500",
---- 925=>x"3900", 926=>x"3500", 927=>x"3700", 928=>x"6d00", 929=>x"b300", 930=>x"2e00", 931=>x"2f00",
---- 932=>x"3000", 933=>x"3900", 934=>x"3a00", 935=>x"3600", 936=>x"7400", 937=>x"4600", 938=>x"2900",
---- 939=>x"3200", 940=>x"3400", 941=>x"3800", 942=>x"3700", 943=>x"3b00", 944=>x"7500", 945=>x"bf00",
---- 946=>x"3b00", 947=>x"3000", 948=>x"3000", 949=>x"3a00", 950=>x"3800", 951=>x"3b00", 952=>x"8400",
---- 953=>x"4600", 954=>x"3500", 955=>x"3100", 956=>x"2f00", 957=>x"3900", 958=>x"3700", 959=>x"3800",
---- 960=>x"8f00", 961=>x"4f00", 962=>x"3500", 963=>x"3800", 964=>x"3a00", 965=>x"4100", 966=>x"3a00",
---- 967=>x"3c00", 968=>x"9600", 969=>x"5100", 970=>x"4400", 971=>x"3b00", 972=>x"3d00", 973=>x"4900",
---- 974=>x"3b00", 975=>x"3800", 976=>x"9e00", 977=>x"5a00", 978=>x"3f00", 979=>x"3a00", 980=>x"3d00",
---- 981=>x"3c00", 982=>x"3f00", 983=>x"3c00", 984=>x"a300", 985=>x"6e00", 986=>x"3800", 987=>x"3600",
---- 988=>x"4500", 989=>x"3f00", 990=>x"3700", 991=>x"3b00", 992=>x"ac00", 993=>x"7c00", 994=>x"3d00",
---- 995=>x"3000", 996=>x"3d00", 997=>x"4500", 998=>x"3e00", 999=>x"3d00", 1000=>x"a900", 1001=>x"8400",
---- 1002=>x"4800", 1003=>x"3500", 1004=>x"3600", 1005=>x"4400", 1006=>x"4600", 1007=>x"4300", 1008=>x"a800",
---- 1009=>x"8400", 1010=>x"5400", 1011=>x"3400", 1012=>x"3400", 1013=>x"b900", 1014=>x"3f00", 1015=>x"3c00",
---- 1016=>x"ad00", 1017=>x"8000", 1018=>x"5f00", 1019=>x"3600", 1020=>x"2e00", 1021=>x"3e00", 1022=>x"3e00",
---- 1023=>x"3e00", 1024=>x"b100", 1025=>x"7900", 1026=>x"6a00", 1027=>x"3b00", 1028=>x"2c00", 1029=>x"4300",
---- 1030=>x"4500", 1031=>x"4000", 1032=>x"b300", 1033=>x"8200", 1034=>x"6700", 1035=>x"4c00", 1036=>x"3100",
---- 1037=>x"c200", 1038=>x"4700", 1039=>x"3c00", 1040=>x"b400", 1041=>x"8200", 1042=>x"6100", 1043=>x"4e00",
---- 1044=>x"3c00", 1045=>x"3a00", 1046=>x"4400", 1047=>x"3a00", 1048=>x"b800", 1049=>x"8900", 1050=>x"5a00",
---- 1051=>x"4b00", 1052=>x"3900", 1053=>x"4300", 1054=>x"4b00", 1055=>x"3c00", 1056=>x"b700", 1057=>x"8900",
---- 1058=>x"5c00", 1059=>x"5800", 1060=>x"3d00", 1061=>x"4700", 1062=>x"4a00", 1063=>x"3c00", 1064=>x"b600",
---- 1065=>x"8f00", 1066=>x"5b00", 1067=>x"5d00", 1068=>x"4400", 1069=>x"4c00", 1070=>x"4400", 1071=>x"3b00",
---- 1072=>x"b800", 1073=>x"9c00", 1074=>x"5600", 1075=>x"5d00", 1076=>x"4c00", 1077=>x"5300", 1078=>x"4100",
---- 1079=>x"3c00", 1080=>x"b700", 1081=>x"a000", 1082=>x"5900", 1083=>x"5200", 1084=>x"ad00", 1085=>x"5300",
---- 1086=>x"3f00", 1087=>x"3700", 1088=>x"b300", 1089=>x"a500", 1090=>x"5e00", 1091=>x"4c00", 1092=>x"5900",
---- 1093=>x"5700", 1094=>x"4200", 1095=>x"3100", 1096=>x"b100", 1097=>x"ad00", 1098=>x"6a00", 1099=>x"4f00",
---- 1100=>x"5f00", 1101=>x"4d00", 1102=>x"3d00", 1103=>x"3700", 1104=>x"a700", 1105=>x"b100", 1106=>x"7700",
---- 1107=>x"4d00", 1108=>x"5c00", 1109=>x"4c00", 1110=>x"3d00", 1111=>x"3700", 1112=>x"a700", 1113=>x"b400",
---- 1114=>x"8500", 1115=>x"4f00", 1116=>x"5600", 1117=>x"5300", 1118=>x"3500", 1119=>x"3000", 1120=>x"a100",
---- 1121=>x"b700", 1122=>x"6d00", 1123=>x"5600", 1124=>x"4f00", 1125=>x"4f00", 1126=>x"3200", 1127=>x"3500",
---- 1128=>x"a000", 1129=>x"b400", 1130=>x"9300", 1131=>x"5b00", 1132=>x"4200", 1133=>x"4c00", 1134=>x"3300",
---- 1135=>x"3200", 1136=>x"a000", 1137=>x"b500", 1138=>x"9500", 1139=>x"6000", 1140=>x"4500", 1141=>x"4e00",
---- 1142=>x"3000", 1143=>x"3400", 1144=>x"9e00", 1145=>x"b300", 1146=>x"a100", 1147=>x"6100", 1148=>x"4000",
---- 1149=>x"4b00", 1150=>x"2b00", 1151=>x"3700", 1152=>x"9c00", 1153=>x"b400", 1154=>x"aa00", 1155=>x"6700",
---- 1156=>x"3b00", 1157=>x"4400", 1158=>x"2600", 1159=>x"3700", 1160=>x"9a00", 1161=>x"ad00", 1162=>x"a800",
---- 1163=>x"9100", 1164=>x"3900", 1165=>x"3a00", 1166=>x"2400", 1167=>x"3c00", 1168=>x"9300", 1169=>x"af00",
---- 1170=>x"a500", 1171=>x"8100", 1172=>x"3c00", 1173=>x"3900", 1174=>x"2600", 1175=>x"3700", 1176=>x"8e00",
---- 1177=>x"ac00", 1178=>x"9d00", 1179=>x"9400", 1180=>x"4200", 1181=>x"3100", 1182=>x"2900", 1183=>x"2d00",
---- 1184=>x"8800", 1185=>x"ac00", 1186=>x"8d00", 1187=>x"9b00", 1188=>x"4d00", 1189=>x"2800", 1190=>x"2400",
---- 1191=>x"2b00", 1192=>x"8000", 1193=>x"ad00", 1194=>x"8a00", 1195=>x"a200", 1196=>x"5d00", 1197=>x"2400",
---- 1198=>x"2a00", 1199=>x"2d00", 1200=>x"7f00", 1201=>x"b300", 1202=>x"9100", 1203=>x"a100", 1204=>x"6d00",
---- 1205=>x"2500", 1206=>x"2800", 1207=>x"2b00", 1208=>x"7300", 1209=>x"4800", 1210=>x"9400", 1211=>x"9800",
---- 1212=>x"8200", 1213=>x"3000", 1214=>x"2700", 1215=>x"2500", 1216=>x"6a00", 1217=>x"ad00", 1218=>x"9600",
---- 1219=>x"9100", 1220=>x"8400", 1221=>x"4300", 1222=>x"2b00", 1223=>x"2a00", 1224=>x"6000", 1225=>x"a700",
---- 1226=>x"9400", 1227=>x"8e00", 1228=>x"8900", 1229=>x"4c00", 1230=>x"2300", 1231=>x"2d00", 1232=>x"5700",
---- 1233=>x"a300", 1234=>x"9a00", 1235=>x"9100", 1236=>x"9300", 1237=>x"5200", 1238=>x"1b00", 1239=>x"2b00",
---- 1240=>x"4e00", 1241=>x"9900", 1242=>x"a300", 1243=>x"9100", 1244=>x"9700", 1245=>x"5600", 1246=>x"1c00",
---- 1247=>x"3000", 1248=>x"4900", 1249=>x"9200", 1250=>x"a400", 1251=>x"8e00", 1252=>x"9900", 1253=>x"6000",
---- 1254=>x"2400", 1255=>x"2f00", 1256=>x"4000", 1257=>x"8300", 1258=>x"a400", 1259=>x"9000", 1260=>x"9a00",
---- 1261=>x"7300", 1262=>x"3300", 1263=>x"2b00", 1264=>x"3200", 1265=>x"7a00", 1266=>x"a700", 1267=>x"9800",
---- 1268=>x"9c00", 1269=>x"8200", 1270=>x"3c00", 1271=>x"2d00", 1272=>x"2d00", 1273=>x"6e00", 1274=>x"a800",
---- 1275=>x"9d00", 1276=>x"9600", 1277=>x"8500", 1278=>x"4600", 1279=>x"2c00", 1280=>x"2900", 1281=>x"6000",
---- 1282=>x"a500", 1283=>x"a400", 1284=>x"9400", 1285=>x"8200", 1286=>x"5000", 1287=>x"2a00", 1288=>x"2300",
---- 1289=>x"5500", 1290=>x"a200", 1291=>x"a800", 1292=>x"8f00", 1293=>x"8900", 1294=>x"5700", 1295=>x"2800",
---- 1296=>x"2100", 1297=>x"4600", 1298=>x"9a00", 1299=>x"ab00", 1300=>x"8500", 1301=>x"8d00", 1302=>x"5f00",
---- 1303=>x"2700", 1304=>x"2100", 1305=>x"3700", 1306=>x"9100", 1307=>x"ac00", 1308=>x"8a00", 1309=>x"8f00",
---- 1310=>x"6a00", 1311=>x"2b00", 1312=>x"dc00", 1313=>x"2d00", 1314=>x"8800", 1315=>x"af00", 1316=>x"8b00",
---- 1317=>x"8d00", 1318=>x"7100", 1319=>x"3600", 1320=>x"2900", 1321=>x"2800", 1322=>x"7a00", 1323=>x"ae00",
---- 1324=>x"8b00", 1325=>x"8600", 1326=>x"6c00", 1327=>x"3f00", 1328=>x"2900", 1329=>x"2300", 1330=>x"6900",
---- 1331=>x"ac00", 1332=>x"9000", 1333=>x"8200", 1334=>x"6800", 1335=>x"4600", 1336=>x"3000", 1337=>x"2400",
---- 1338=>x"5900", 1339=>x"a800", 1340=>x"9700", 1341=>x"8700", 1342=>x"6700", 1343=>x"4f00", 1344=>x"2b00",
---- 1345=>x"2300", 1346=>x"4a00", 1347=>x"9d00", 1348=>x"9f00", 1349=>x"8900", 1350=>x"6600", 1351=>x"5e00",
---- 1352=>x"2800", 1353=>x"2300", 1354=>x"4300", 1355=>x"9500", 1356=>x"9b00", 1357=>x"8500", 1358=>x"6600",
---- 1359=>x"6200", 1360=>x"2c00", 1361=>x"2600", 1362=>x"4500", 1363=>x"8e00", 1364=>x"9f00", 1365=>x"8000",
---- 1366=>x"6700", 1367=>x"6b00", 1368=>x"2b00", 1369=>x"2300", 1370=>x"c100", 1371=>x"8800", 1372=>x"a300",
---- 1373=>x"8400", 1374=>x"6d00", 1375=>x"6600", 1376=>x"2800", 1377=>x"2300", 1378=>x"3300", 1379=>x"8000",
---- 1380=>x"a600", 1381=>x"8500", 1382=>x"7100", 1383=>x"6f00", 1384=>x"2700", 1385=>x"2700", 1386=>x"2d00",
---- 1387=>x"7800", 1388=>x"a700", 1389=>x"8100", 1390=>x"7400", 1391=>x"7900", 1392=>x"2600", 1393=>x"2700",
---- 1394=>x"2a00", 1395=>x"6c00", 1396=>x"a500", 1397=>x"7e00", 1398=>x"7700", 1399=>x"8200", 1400=>x"2e00",
---- 1401=>x"2800", 1402=>x"2a00", 1403=>x"5e00", 1404=>x"a000", 1405=>x"8700", 1406=>x"8600", 1407=>x"8800",
---- 1408=>x"2f00", 1409=>x"2a00", 1410=>x"2c00", 1411=>x"5300", 1412=>x"9c00", 1413=>x"8d00", 1414=>x"8a00",
---- 1415=>x"9000", 1416=>x"3100", 1417=>x"2d00", 1418=>x"2b00", 1419=>x"4b00", 1420=>x"9500", 1421=>x"9400",
---- 1422=>x"8a00", 1423=>x"9500", 1424=>x"3600", 1425=>x"2800", 1426=>x"2d00", 1427=>x"4a00", 1428=>x"9700",
---- 1429=>x"9d00", 1430=>x"8e00", 1431=>x"9500", 1432=>x"3e00", 1433=>x"d300", 1434=>x"2e00", 1435=>x"4900",
---- 1436=>x"9100", 1437=>x"a000", 1438=>x"9000", 1439=>x"9700", 1440=>x"3e00", 1441=>x"2f00", 1442=>x"3000",
---- 1443=>x"4800", 1444=>x"8e00", 1445=>x"a300", 1446=>x"9600", 1447=>x"9a00", 1448=>x"4300", 1449=>x"3000",
---- 1450=>x"2f00", 1451=>x"4300", 1452=>x"9000", 1453=>x"a400", 1454=>x"9700", 1455=>x"9900", 1456=>x"4400",
---- 1457=>x"2e00", 1458=>x"2f00", 1459=>x"4000", 1460=>x"8800", 1461=>x"a600", 1462=>x"9300", 1463=>x"9900",
---- 1464=>x"4300", 1465=>x"3700", 1466=>x"3700", 1467=>x"3f00", 1468=>x"8900", 1469=>x"ae00", 1470=>x"9600",
---- 1471=>x"9c00", 1472=>x"4d00", 1473=>x"3100", 1474=>x"3200", 1475=>x"3700", 1476=>x"8600", 1477=>x"ac00",
---- 1478=>x"6700", 1479=>x"9c00", 1480=>x"4a00", 1481=>x"3100", 1482=>x"3800", 1483=>x"3500", 1484=>x"8300",
---- 1485=>x"ad00", 1486=>x"9e00", 1487=>x"9e00", 1488=>x"4800", 1489=>x"3800", 1490=>x"3900", 1491=>x"3600",
---- 1492=>x"8000", 1493=>x"b000", 1494=>x"9f00", 1495=>x"a300", 1496=>x"4000", 1497=>x"4500", 1498=>x"3800",
---- 1499=>x"3500", 1500=>x"8400", 1501=>x"ae00", 1502=>x"9c00", 1503=>x"a200", 1504=>x"3d00", 1505=>x"4e00",
---- 1506=>x"3300", 1507=>x"3000", 1508=>x"8200", 1509=>x"af00", 1510=>x"9e00", 1511=>x"a000", 1512=>x"3e00",
---- 1513=>x"4f00", 1514=>x"3d00", 1515=>x"3000", 1516=>x"7d00", 1517=>x"b500", 1518=>x"9f00", 1519=>x"a100",
---- 1520=>x"3f00", 1521=>x"5100", 1522=>x"3c00", 1523=>x"3000", 1524=>x"8000", 1525=>x"b100", 1526=>x"9d00",
---- 1527=>x"a300", 1528=>x"4400", 1529=>x"5600", 1530=>x"3c00", 1531=>x"3000", 1532=>x"8200", 1533=>x"ae00",
---- 1534=>x"9a00", 1535=>x"9f00", 1536=>x"4400", 1537=>x"5400", 1538=>x"3f00", 1539=>x"3600", 1540=>x"8d00",
---- 1541=>x"ad00", 1542=>x"9900", 1543=>x"9d00", 1544=>x"4200", 1545=>x"4e00", 1546=>x"4600", 1547=>x"3a00",
---- 1548=>x"8c00", 1549=>x"ae00", 1550=>x"9900", 1551=>x"9900", 1552=>x"4100", 1553=>x"4b00", 1554=>x"4600",
---- 1555=>x"4100", 1556=>x"9300", 1557=>x"ac00", 1558=>x"9700", 1559=>x"9200", 1560=>x"4600", 1561=>x"4c00",
---- 1562=>x"4400", 1563=>x"4500", 1564=>x"9900", 1565=>x"a300", 1566=>x"9a00", 1567=>x"8900", 1568=>x"4b00",
---- 1569=>x"4e00", 1570=>x"4200", 1571=>x"4600", 1572=>x"9c00", 1573=>x"a100", 1574=>x"9900", 1575=>x"8300",
---- 1576=>x"4900", 1577=>x"5200", 1578=>x"4a00", 1579=>x"b200", 1580=>x"a400", 1581=>x"9d00", 1582=>x"6b00",
---- 1583=>x"8000", 1584=>x"4400", 1585=>x"4e00", 1586=>x"4500", 1587=>x"5000", 1588=>x"aa00", 1589=>x"9b00",
---- 1590=>x"9000", 1591=>x"7e00", 1592=>x"4500", 1593=>x"4600", 1594=>x"3c00", 1595=>x"5700", 1596=>x"a700",
---- 1597=>x"9700", 1598=>x"8f00", 1599=>x"8000", 1600=>x"4700", 1601=>x"4b00", 1602=>x"3e00", 1603=>x"a200",
---- 1604=>x"a600", 1605=>x"9600", 1606=>x"8f00", 1607=>x"8800", 1608=>x"4b00", 1609=>x"4700", 1610=>x"3900",
---- 1611=>x"6500", 1612=>x"a500", 1613=>x"9500", 1614=>x"7500", 1615=>x"8b00", 1616=>x"4600", 1617=>x"4000",
---- 1618=>x"3700", 1619=>x"7500", 1620=>x"a700", 1621=>x"9200", 1622=>x"8600", 1623=>x"8e00", 1624=>x"4600",
---- 1625=>x"3900", 1626=>x"3600", 1627=>x"7c00", 1628=>x"a300", 1629=>x"8f00", 1630=>x"8900", 1631=>x"9500",
---- 1632=>x"ba00", 1633=>x"3200", 1634=>x"3100", 1635=>x"8100", 1636=>x"a100", 1637=>x"9000", 1638=>x"8600",
---- 1639=>x"9500", 1640=>x"4300", 1641=>x"3300", 1642=>x"3800", 1643=>x"8d00", 1644=>x"a000", 1645=>x"9000",
---- 1646=>x"8800", 1647=>x"9400", 1648=>x"4d00", 1649=>x"2f00", 1650=>x"3c00", 1651=>x"6600", 1652=>x"9900",
---- 1653=>x"8e00", 1654=>x"8a00", 1655=>x"9300", 1656=>x"4600", 1657=>x"2c00", 1658=>x"4500", 1659=>x"9d00",
---- 1660=>x"9400", 1661=>x"8a00", 1662=>x"8d00", 1663=>x"9300", 1664=>x"c500", 1665=>x"2400", 1666=>x"4d00",
---- 1667=>x"a500", 1668=>x"9000", 1669=>x"8b00", 1670=>x"9100", 1671=>x"9400", 1672=>x"3b00", 1673=>x"2400",
---- 1674=>x"5b00", 1675=>x"a400", 1676=>x"8b00", 1677=>x"8800", 1678=>x"9000", 1679=>x"9100", 1680=>x"3800",
---- 1681=>x"2300", 1682=>x"6900", 1683=>x"a200", 1684=>x"8600", 1685=>x"8900", 1686=>x"8f00", 1687=>x"9300",
---- 1688=>x"2d00", 1689=>x"2200", 1690=>x"7000", 1691=>x"9e00", 1692=>x"8600", 1693=>x"8800", 1694=>x"9400",
---- 1695=>x"9600", 1696=>x"2500", 1697=>x"2a00", 1698=>x"7d00", 1699=>x"a100", 1700=>x"8900", 1701=>x"8900",
---- 1702=>x"9500", 1703=>x"9600", 1704=>x"2200", 1705=>x"2d00", 1706=>x"8600", 1707=>x"9d00", 1708=>x"8c00",
---- 1709=>x"8900", 1710=>x"9800", 1711=>x"6a00", 1712=>x"1e00", 1713=>x"3400", 1714=>x"8b00", 1715=>x"9c00",
---- 1716=>x"8d00", 1717=>x"8d00", 1718=>x"9600", 1719=>x"9600", 1720=>x"1f00", 1721=>x"3f00", 1722=>x"8e00",
---- 1723=>x"9600", 1724=>x"8d00", 1725=>x"8f00", 1726=>x"9600", 1727=>x"9300", 1728=>x"1b00", 1729=>x"4900",
---- 1730=>x"9600", 1731=>x"8d00", 1732=>x"8e00", 1733=>x"9400", 1734=>x"9500", 1735=>x"9400", 1736=>x"1b00",
---- 1737=>x"5900", 1738=>x"9300", 1739=>x"8e00", 1740=>x"8e00", 1741=>x"9700", 1742=>x"9400", 1743=>x"9500",
---- 1744=>x"1d00", 1745=>x"6300", 1746=>x"8f00", 1747=>x"8e00", 1748=>x"8f00", 1749=>x"9b00", 1750=>x"9300",
---- 1751=>x"9400", 1752=>x"2300", 1753=>x"6e00", 1754=>x"8c00", 1755=>x"8d00", 1756=>x"8f00", 1757=>x"9900",
---- 1758=>x"9600", 1759=>x"9000", 1760=>x"2500", 1761=>x"7400", 1762=>x"8b00", 1763=>x"8b00", 1764=>x"9100",
---- 1765=>x"9400", 1766=>x"9700", 1767=>x"8f00", 1768=>x"2b00", 1769=>x"7700", 1770=>x"8c00", 1771=>x"8c00",
---- 1772=>x"9200", 1773=>x"9700", 1774=>x"9b00", 1775=>x"8f00", 1776=>x"3300", 1777=>x"7d00", 1778=>x"8a00",
---- 1779=>x"8e00", 1780=>x"9100", 1781=>x"9000", 1782=>x"6700", 1783=>x"9500", 1784=>x"3b00", 1785=>x"8500",
---- 1786=>x"8b00", 1787=>x"8f00", 1788=>x"8f00", 1789=>x"9100", 1790=>x"9500", 1791=>x"9800", 1792=>x"3e00",
---- 1793=>x"8400", 1794=>x"8b00", 1795=>x"8e00", 1796=>x"9200", 1797=>x"9500", 1798=>x"9400", 1799=>x"9700",
---- 1800=>x"3f00", 1801=>x"8500", 1802=>x"8d00", 1803=>x"9200", 1804=>x"9400", 1805=>x"9700", 1806=>x"9300",
---- 1807=>x"9200", 1808=>x"4700", 1809=>x"8500", 1810=>x"8f00", 1811=>x"8f00", 1812=>x"8e00", 1813=>x"9600",
---- 1814=>x"9500", 1815=>x"9100", 1816=>x"5f00", 1817=>x"8700", 1818=>x"9000", 1819=>x"8c00", 1820=>x"7f00",
---- 1821=>x"8900", 1822=>x"8c00", 1823=>x"8d00", 1824=>x"7b00", 1825=>x"8600", 1826=>x"9300", 1827=>x"8300",
---- 1828=>x"7100", 1829=>x"7900", 1830=>x"7f00", 1831=>x"8000", 1832=>x"9a00", 1833=>x"8800", 1834=>x"8f00",
---- 1835=>x"7100", 1836=>x"6000", 1837=>x"6b00", 1838=>x"6d00", 1839=>x"7200", 1840=>x"b600", 1841=>x"8700",
---- 1842=>x"7900", 1843=>x"6100", 1844=>x"4f00", 1845=>x"5f00", 1846=>x"5f00", 1847=>x"5d00", 1848=>x"cd00",
---- 1849=>x"7800", 1850=>x"5b00", 1851=>x"4f00", 1852=>x"4500", 1853=>x"5200", 1854=>x"5000", 1855=>x"5000",
---- 1856=>x"da00", 1857=>x"8900", 1858=>x"4800", 1859=>x"4f00", 1860=>x"4800", 1861=>x"5000", 1862=>x"4500",
---- 1863=>x"4700", 1864=>x"df00", 1865=>x"9f00", 1866=>x"4800", 1867=>x"5500", 1868=>x"5300", 1869=>x"5c00",
---- 1870=>x"4d00", 1871=>x"4d00", 1872=>x"df00", 1873=>x"b900", 1874=>x"5000", 1875=>x"5000", 1876=>x"5800",
---- 1877=>x"5d00", 1878=>x"5900", 1879=>x"5900", 1880=>x"db00", 1881=>x"d200", 1882=>x"6200", 1883=>x"4900",
---- 1884=>x"5d00", 1885=>x"5f00", 1886=>x"6200", 1887=>x"5d00", 1888=>x"d800", 1889=>x"dc00", 1890=>x"8a00",
---- 1891=>x"4a00", 1892=>x"5d00", 1893=>x"6200", 1894=>x"6700", 1895=>x"6500", 1896=>x"d700", 1897=>x"dd00",
---- 1898=>x"ae00", 1899=>x"5100", 1900=>x"5b00", 1901=>x"6200", 1902=>x"6a00", 1903=>x"6900", 1904=>x"d700",
---- 1905=>x"dc00", 1906=>x"c700", 1907=>x"6400", 1908=>x"5500", 1909=>x"6200", 1910=>x"6500", 1911=>x"6a00",
---- 1912=>x"d700", 1913=>x"d900", 1914=>x"d900", 1915=>x"7c00", 1916=>x"4b00", 1917=>x"5d00", 1918=>x"6500",
---- 1919=>x"6a00", 1920=>x"d500", 1921=>x"d700", 1922=>x"dc00", 1923=>x"9c00", 1924=>x"4b00", 1925=>x"5900",
---- 1926=>x"6300", 1927=>x"6b00", 1928=>x"d400", 1929=>x"d800", 1930=>x"db00", 1931=>x"bc00", 1932=>x"5a00",
---- 1933=>x"5300", 1934=>x"5d00", 1935=>x"6300", 1936=>x"d400", 1937=>x"d800", 1938=>x"d800", 1939=>x"d200",
---- 1940=>x"7300", 1941=>x"4d00", 1942=>x"5c00", 1943=>x"6100", 1944=>x"d500", 1945=>x"d800", 1946=>x"d700",
---- 1947=>x"d900", 1948=>x"8b00", 1949=>x"4a00", 1950=>x"5b00", 1951=>x"6100", 1952=>x"2a00", 1953=>x"d700",
---- 1954=>x"d600", 1955=>x"da00", 1956=>x"ab00", 1957=>x"4e00", 1958=>x"5300", 1959=>x"5f00", 1960=>x"d300",
---- 1961=>x"d700", 1962=>x"d500", 1963=>x"d700", 1964=>x"c700", 1965=>x"6100", 1966=>x"4e00", 1967=>x"5a00",
---- 1968=>x"d400", 1969=>x"d700", 1970=>x"d700", 1971=>x"d600", 1972=>x"d400", 1973=>x"7700", 1974=>x"4900",
---- 1975=>x"5700", 1976=>x"d400", 1977=>x"d400", 1978=>x"d600", 1979=>x"d600", 1980=>x"db00", 1981=>x"9700",
---- 1982=>x"4900", 1983=>x"5300", 1984=>x"d300", 1985=>x"d400", 1986=>x"d500", 1987=>x"d500", 1988=>x"d800",
---- 1989=>x"b500", 1990=>x"5400", 1991=>x"4c00", 1992=>x"d200", 1993=>x"d200", 1994=>x"d400", 1995=>x"d500",
---- 1996=>x"d700", 1997=>x"c600", 1998=>x"6100", 1999=>x"4400", 2000=>x"d200", 2001=>x"d000", 2002=>x"d100",
---- 2003=>x"d300", 2004=>x"d500", 2005=>x"d300", 2006=>x"7900", 2007=>x"4000", 2008=>x"d000", 2009=>x"d100",
---- 2010=>x"d100", 2011=>x"d200", 2012=>x"d600", 2013=>x"d800", 2014=>x"9800", 2015=>x"4500", 2016=>x"cf00",
---- 2017=>x"d200", 2018=>x"d300", 2019=>x"d300", 2020=>x"d300", 2021=>x"d900", 2022=>x"b500", 2023=>x"4d00",
---- 2024=>x"cd00", 2025=>x"d000", 2026=>x"d300", 2027=>x"d300", 2028=>x"d300", 2029=>x"d500", 2030=>x"c900",
---- 2031=>x"6400", 2032=>x"cd00", 2033=>x"d000", 2034=>x"d200", 2035=>x"d000", 2036=>x"d400", 2037=>x"d500",
---- 2038=>x"2800", 2039=>x"8200", 2040=>x"cc00", 2041=>x"cf00", 2042=>x"d100", 2043=>x"d100", 2044=>x"d300",
---- 2045=>x"d300", 2046=>x"d700", 2047=>x"9b00"),
---- 24 => (0=>x"9b00", 1=>x"9c00", 2=>x"9e00", 3=>x"9b00", 4=>x"9c00", 5=>x"a000", 6=>x"9d00", 7=>x"9b00",
---- 8=>x"9a00", 9=>x"9c00", 10=>x"9e00", 11=>x"9b00", 12=>x"9c00", 13=>x"a000", 14=>x"9c00",
---- 15=>x"9b00", 16=>x"9a00", 17=>x"9c00", 18=>x"9e00", 19=>x"9b00", 20=>x"9c00", 21=>x"9e00",
---- 22=>x"9d00", 23=>x"9b00", 24=>x"9700", 25=>x"9a00", 26=>x"9b00", 27=>x"9a00", 28=>x"9c00",
---- 29=>x"9b00", 30=>x"9c00", 31=>x"9a00", 32=>x"9b00", 33=>x"9b00", 34=>x"9a00", 35=>x"9a00",
---- 36=>x"9b00", 37=>x"9c00", 38=>x"9900", 39=>x"9a00", 40=>x"6500", 41=>x"9c00", 42=>x"9800",
---- 43=>x"9a00", 44=>x"9900", 45=>x"9900", 46=>x"9900", 47=>x"9800", 48=>x"9900", 49=>x"9900",
---- 50=>x"9800", 51=>x"9900", 52=>x"9900", 53=>x"9a00", 54=>x"9a00", 55=>x"9800", 56=>x"9b00",
---- 57=>x"9b00", 58=>x"9800", 59=>x"9800", 60=>x"9500", 61=>x"9800", 62=>x"9900", 63=>x"9900",
---- 64=>x"9900", 65=>x"9b00", 66=>x"9b00", 67=>x"9700", 68=>x"9800", 69=>x"9500", 70=>x"9900",
---- 71=>x"9800", 72=>x"6700", 73=>x"9b00", 74=>x"9b00", 75=>x"9900", 76=>x"9800", 77=>x"9700",
---- 78=>x"9800", 79=>x"9800", 80=>x"9d00", 81=>x"9c00", 82=>x"9900", 83=>x"9800", 84=>x"9700",
---- 85=>x"9700", 86=>x"9700", 87=>x"9b00", 88=>x"9a00", 89=>x"9a00", 90=>x"9700", 91=>x"9a00",
---- 92=>x"9700", 93=>x"9800", 94=>x"9700", 95=>x"9700", 96=>x"9b00", 97=>x"9a00", 98=>x"9900",
---- 99=>x"9700", 100=>x"9700", 101=>x"9800", 102=>x"9700", 103=>x"9700", 104=>x"9b00", 105=>x"9a00",
---- 106=>x"9900", 107=>x"9900", 108=>x"9900", 109=>x"9900", 110=>x"9800", 111=>x"9800", 112=>x"9d00",
---- 113=>x"9a00", 114=>x"9c00", 115=>x"9a00", 116=>x"9a00", 117=>x"9c00", 118=>x"6300", 119=>x"9600",
---- 120=>x"9d00", 121=>x"6400", 122=>x"9b00", 123=>x"9c00", 124=>x"9c00", 125=>x"6200", 126=>x"9b00",
---- 127=>x"9b00", 128=>x"9e00", 129=>x"9d00", 130=>x"9b00", 131=>x"9c00", 132=>x"9d00", 133=>x"9d00",
---- 134=>x"9a00", 135=>x"9b00", 136=>x"9d00", 137=>x"9d00", 138=>x"9c00", 139=>x"9a00", 140=>x"9c00",
---- 141=>x"9a00", 142=>x"9b00", 143=>x"9e00", 144=>x"9d00", 145=>x"9c00", 146=>x"9c00", 147=>x"9b00",
---- 148=>x"9d00", 149=>x"9b00", 150=>x"9a00", 151=>x"9b00", 152=>x"9c00", 153=>x"9e00", 154=>x"9e00",
---- 155=>x"9d00", 156=>x"9c00", 157=>x"9d00", 158=>x"9b00", 159=>x"9a00", 160=>x"9a00", 161=>x"9c00",
---- 162=>x"9f00", 163=>x"9d00", 164=>x"9b00", 165=>x"9b00", 166=>x"9c00", 167=>x"9900", 168=>x"9900",
---- 169=>x"9800", 170=>x"9900", 171=>x"9c00", 172=>x"9d00", 173=>x"9b00", 174=>x"9a00", 175=>x"9800",
---- 176=>x"9b00", 177=>x"9a00", 178=>x"9700", 179=>x"9c00", 180=>x"9b00", 181=>x"9800", 182=>x"6700",
---- 183=>x"9600", 184=>x"9b00", 185=>x"9b00", 186=>x"9900", 187=>x"9900", 188=>x"9800", 189=>x"9800",
---- 190=>x"9600", 191=>x"9500", 192=>x"9900", 193=>x"9b00", 194=>x"9700", 195=>x"9600", 196=>x"9700",
---- 197=>x"9800", 198=>x"9600", 199=>x"9400", 200=>x"9a00", 201=>x"9b00", 202=>x"9600", 203=>x"9800",
---- 204=>x"9800", 205=>x"9400", 206=>x"9300", 207=>x"9400", 208=>x"9700", 209=>x"9800", 210=>x"9700",
---- 211=>x"9700", 212=>x"9300", 213=>x"9100", 214=>x"9200", 215=>x"9100", 216=>x"9300", 217=>x"9500",
---- 218=>x"9400", 219=>x"9400", 220=>x"9200", 221=>x"9100", 222=>x"8f00", 223=>x"8e00", 224=>x"9100",
---- 225=>x"9400", 226=>x"9200", 227=>x"9200", 228=>x"9100", 229=>x"9100", 230=>x"9000", 231=>x"9100",
---- 232=>x"9100", 233=>x"9100", 234=>x"9200", 235=>x"9100", 236=>x"9300", 237=>x"9000", 238=>x"8f00",
---- 239=>x"8f00", 240=>x"9100", 241=>x"8f00", 242=>x"9100", 243=>x"9200", 244=>x"9200", 245=>x"9300",
---- 246=>x"9000", 247=>x"8f00", 248=>x"8e00", 249=>x"8f00", 250=>x"9000", 251=>x"9100", 252=>x"9200",
---- 253=>x"9200", 254=>x"8e00", 255=>x"9000", 256=>x"8c00", 257=>x"8e00", 258=>x"8e00", 259=>x"8f00",
---- 260=>x"8f00", 261=>x"8f00", 262=>x"8f00", 263=>x"9000", 264=>x"8b00", 265=>x"8f00", 266=>x"8d00",
---- 267=>x"8e00", 268=>x"8e00", 269=>x"9300", 270=>x"9300", 271=>x"8e00", 272=>x"8d00", 273=>x"8d00",
---- 274=>x"8e00", 275=>x"9000", 276=>x"9100", 277=>x"9200", 278=>x"9300", 279=>x"8f00", 280=>x"8e00",
---- 281=>x"8f00", 282=>x"9100", 283=>x"9000", 284=>x"9100", 285=>x"9100", 286=>x"9300", 287=>x"8f00",
---- 288=>x"8f00", 289=>x"8e00", 290=>x"9000", 291=>x"8f00", 292=>x"9100", 293=>x"9200", 294=>x"9000",
---- 295=>x"8f00", 296=>x"9000", 297=>x"8e00", 298=>x"9000", 299=>x"9300", 300=>x"9300", 301=>x"9500",
---- 302=>x"9400", 303=>x"8e00", 304=>x"9100", 305=>x"8f00", 306=>x"9100", 307=>x"9300", 308=>x"9400",
---- 309=>x"9500", 310=>x"9400", 311=>x"8f00", 312=>x"9200", 313=>x"9100", 314=>x"9100", 315=>x"9100",
---- 316=>x"9200", 317=>x"9300", 318=>x"9200", 319=>x"8f00", 320=>x"9400", 321=>x"9300", 322=>x"8e00",
---- 323=>x"9100", 324=>x"8f00", 325=>x"9100", 326=>x"9200", 327=>x"9000", 328=>x"9600", 329=>x"9300",
---- 330=>x"9000", 331=>x"8d00", 332=>x"9000", 333=>x"9200", 334=>x"9200", 335=>x"9000", 336=>x"9400",
---- 337=>x"9300", 338=>x"9400", 339=>x"9000", 340=>x"9100", 341=>x"9400", 342=>x"9300", 343=>x"9200",
---- 344=>x"9200", 345=>x"9400", 346=>x"9400", 347=>x"9000", 348=>x"8e00", 349=>x"8f00", 350=>x"9200",
---- 351=>x"9300", 352=>x"8f00", 353=>x"9500", 354=>x"9600", 355=>x"9400", 356=>x"8f00", 357=>x"9000",
---- 358=>x"9000", 359=>x"9200", 360=>x"8c00", 361=>x"9300", 362=>x"9400", 363=>x"9600", 364=>x"9100",
---- 365=>x"8f00", 366=>x"9200", 367=>x"9100", 368=>x"8600", 369=>x"9000", 370=>x"9300", 371=>x"9600",
---- 372=>x"9500", 373=>x"8f00", 374=>x"9200", 375=>x"9000", 376=>x"8200", 377=>x"8c00", 378=>x"6f00",
---- 379=>x"9500", 380=>x"9600", 381=>x"9300", 382=>x"9000", 383=>x"9200", 384=>x"7b00", 385=>x"8600",
---- 386=>x"8b00", 387=>x"9300", 388=>x"9500", 389=>x"9400", 390=>x"9100", 391=>x"8f00", 392=>x"7300",
---- 393=>x"7e00", 394=>x"8600", 395=>x"8f00", 396=>x"9300", 397=>x"9500", 398=>x"9300", 399=>x"9100",
---- 400=>x"6500", 401=>x"7800", 402=>x"8100", 403=>x"8700", 404=>x"9200", 405=>x"9500", 406=>x"9300",
---- 407=>x"9200", 408=>x"5d00", 409=>x"6b00", 410=>x"7d00", 411=>x"8600", 412=>x"8d00", 413=>x"9400",
---- 414=>x"9400", 415=>x"9200", 416=>x"4b00", 417=>x"5e00", 418=>x"8800", 419=>x"7f00", 420=>x"8700",
---- 421=>x"8f00", 422=>x"6d00", 423=>x"9400", 424=>x"c500", 425=>x"5300", 426=>x"6500", 427=>x"7800",
---- 428=>x"8200", 429=>x"8900", 430=>x"8f00", 431=>x"9300", 432=>x"2f00", 433=>x"4100", 434=>x"5800",
---- 435=>x"6d00", 436=>x"7900", 437=>x"8200", 438=>x"8900", 439=>x"8d00", 440=>x"2900", 441=>x"2f00",
---- 442=>x"4400", 443=>x"5a00", 444=>x"6a00", 445=>x"7200", 446=>x"8300", 447=>x"9500", 448=>x"2700",
---- 449=>x"2600", 450=>x"2f00", 451=>x"4000", 452=>x"5800", 453=>x"8a00", 454=>x"b700", 455=>x"ca00",
---- 456=>x"2500", 457=>x"2400", 458=>x"2200", 459=>x"4d00", 460=>x"a200", 461=>x"d100", 462=>x"dc00",
---- 463=>x"dd00", 464=>x"2700", 465=>x"2000", 466=>x"5100", 467=>x"b400", 468=>x"dc00", 469=>x"dd00",
---- 470=>x"d500", 471=>x"c300", 472=>x"2800", 473=>x"6a00", 474=>x"3f00", 475=>x"df00", 476=>x"db00",
---- 477=>x"c400", 478=>x"b900", 479=>x"c400", 480=>x"8400", 481=>x"ce00", 482=>x"de00", 483=>x"d600",
---- 484=>x"b300", 485=>x"af00", 486=>x"cd00", 487=>x"d900", 488=>x"d500", 489=>x"d900", 490=>x"c900",
---- 491=>x"a600", 492=>x"b200", 493=>x"d300", 494=>x"da00", 495=>x"2400", 496=>x"d900", 497=>x"bc00",
---- 498=>x"9f00", 499=>x"b200", 500=>x"d600", 501=>x"db00", 502=>x"da00", 503=>x"d600", 504=>x"af00",
---- 505=>x"9b00", 506=>x"c100", 507=>x"d600", 508=>x"db00", 509=>x"da00", 510=>x"d600", 511=>x"d300",
---- 512=>x"a200", 513=>x"c300", 514=>x"d700", 515=>x"d700", 516=>x"2900", 517=>x"d400", 518=>x"d500",
---- 519=>x"d100", 520=>x"d000", 521=>x"d900", 522=>x"d800", 523=>x"d500", 524=>x"d400", 525=>x"d100",
---- 526=>x"d000", 527=>x"ca00", 528=>x"2900", 529=>x"d800", 530=>x"2e00", 531=>x"cf00", 532=>x"d100",
---- 533=>x"ce00", 534=>x"cb00", 535=>x"c800", 536=>x"d400", 537=>x"d200", 538=>x"ce00", 539=>x"cb00",
---- 540=>x"ce00", 541=>x"ca00", 542=>x"c800", 543=>x"c800", 544=>x"d100", 545=>x"ce00", 546=>x"cb00",
---- 547=>x"cc00", 548=>x"cc00", 549=>x"c800", 550=>x"c800", 551=>x"cb00", 552=>x"cd00", 553=>x"c800",
---- 554=>x"ca00", 555=>x"c900", 556=>x"c800", 557=>x"ca00", 558=>x"cb00", 559=>x"cc00", 560=>x"c800",
---- 561=>x"c900", 562=>x"c800", 563=>x"cb00", 564=>x"cc00", 565=>x"cd00", 566=>x"cb00", 567=>x"cb00",
---- 568=>x"c900", 569=>x"c800", 570=>x"c900", 571=>x"cb00", 572=>x"cd00", 573=>x"cc00", 574=>x"cc00",
---- 575=>x"cc00", 576=>x"c800", 577=>x"ca00", 578=>x"cd00", 579=>x"ce00", 580=>x"cd00", 581=>x"cb00",
---- 582=>x"cb00", 583=>x"c900", 584=>x"c800", 585=>x"cb00", 586=>x"cd00", 587=>x"cd00", 588=>x"cb00",
---- 589=>x"cc00", 590=>x"c900", 591=>x"c300", 592=>x"ca00", 593=>x"cb00", 594=>x"ca00", 595=>x"cd00",
---- 596=>x"cd00", 597=>x"cb00", 598=>x"bf00", 599=>x"c100", 600=>x"ca00", 601=>x"cd00", 602=>x"cc00",
---- 603=>x"cc00", 604=>x"d000", 605=>x"bd00", 606=>x"b200", 607=>x"bc00", 608=>x"cc00", 609=>x"cb00",
---- 610=>x"cd00", 611=>x"d100", 612=>x"c000", 613=>x"a900", 614=>x"a800", 615=>x"b200", 616=>x"ca00",
---- 617=>x"ce00", 618=>x"cd00", 619=>x"c700", 620=>x"ac00", 621=>x"9f00", 622=>x"a200", 623=>x"a700",
---- 624=>x"cf00", 625=>x"cc00", 626=>x"cd00", 627=>x"b500", 628=>x"a200", 629=>x"9c00", 630=>x"9a00",
---- 631=>x"5600", 632=>x"ce00", 633=>x"cd00", 634=>x"c400", 635=>x"a200", 636=>x"9900", 637=>x"9d00",
---- 638=>x"a900", 639=>x"bc00", 640=>x"ce00", 641=>x"d000", 642=>x"aa00", 643=>x"9900", 644=>x"9c00",
---- 645=>x"aa00", 646=>x"bd00", 647=>x"9900", 648=>x"d200", 649=>x"bd00", 650=>x"9800", 651=>x"9e00",
---- 652=>x"ab00", 653=>x"b700", 654=>x"9a00", 655=>x"8000", 656=>x"cf00", 657=>x"a300", 658=>x"9600",
---- 659=>x"a700", 660=>x"b700", 661=>x"9c00", 662=>x"8600", 663=>x"9d00", 664=>x"b300", 665=>x"9200",
---- 666=>x"9f00", 667=>x"af00", 668=>x"9700", 669=>x"8f00", 670=>x"a900", 671=>x"ab00", 672=>x"9600",
---- 673=>x"9e00", 674=>x"ac00", 675=>x"9700", 676=>x"9700", 677=>x"a600", 678=>x"9700", 679=>x"7c00",
---- 680=>x"9800", 681=>x"a700", 682=>x"9800", 683=>x"9700", 684=>x"8b00", 685=>x"7500", 686=>x"5d00",
---- 687=>x"6700", 688=>x"a500", 689=>x"9c00", 690=>x"8d00", 691=>x"6a00", 692=>x"4f00", 693=>x"5900",
---- 694=>x"5f00", 695=>x"7a00", 696=>x"9200", 697=>x"7300", 698=>x"5100", 699=>x"5000", 700=>x"5700",
---- 701=>x"6200", 702=>x"6f00", 703=>x"6800", 704=>x"5b00", 705=>x"4d00", 706=>x"5700", 707=>x"5f00",
---- 708=>x"6000", 709=>x"6b00", 710=>x"8900", 711=>x"b500", 712=>x"5200", 713=>x"5700", 714=>x"5c00",
---- 715=>x"5e00", 716=>x"6600", 717=>x"8200", 718=>x"b000", 719=>x"c700", 720=>x"5700", 721=>x"5c00",
---- 722=>x"5900", 723=>x"9b00", 724=>x"8600", 725=>x"a900", 726=>x"bf00", 727=>x"cc00", 728=>x"5a00",
---- 729=>x"6600", 730=>x"7200", 731=>x"8900", 732=>x"ae00", 733=>x"ba00", 734=>x"c900", 735=>x"db00",
---- 736=>x"6700", 737=>x"8100", 738=>x"9800", 739=>x"ad00", 740=>x"be00", 741=>x"cd00", 742=>x"b900",
---- 743=>x"6d00", 744=>x"8d00", 745=>x"a600", 746=>x"b800", 747=>x"c200", 748=>x"cd00", 749=>x"ba00",
---- 750=>x"4400", 751=>x"2100", 752=>x"a700", 753=>x"b500", 754=>x"bf00", 755=>x"3500", 756=>x"d100",
---- 757=>x"5f00", 758=>x"1f00", 759=>x"3000", 760=>x"b000", 761=>x"b400", 762=>x"c500", 763=>x"c800",
---- 764=>x"6b00", 765=>x"2400", 766=>x"2e00", 767=>x"3100", 768=>x"b000", 769=>x"c300", 770=>x"3400",
---- 771=>x"6100", 772=>x"2300", 773=>x"2a00", 774=>x"2b00", 775=>x"2d00", 776=>x"c400", 777=>x"d300",
---- 778=>x"6a00", 779=>x"1f00", 780=>x"2a00", 781=>x"2b00", 782=>x"2e00", 783=>x"3200", 784=>x"d200",
---- 785=>x"7700", 786=>x"2500", 787=>x"2900", 788=>x"2700", 789=>x"2b00", 790=>x"3000", 791=>x"3300",
---- 792=>x"7900", 793=>x"2000", 794=>x"2b00", 795=>x"2900", 796=>x"2c00", 797=>x"2f00", 798=>x"3100",
---- 799=>x"3300", 800=>x"2b00", 801=>x"2600", 802=>x"2b00", 803=>x"2b00", 804=>x"2f00", 805=>x"3000",
---- 806=>x"3500", 807=>x"3300", 808=>x"2d00", 809=>x"2600", 810=>x"2800", 811=>x"2e00", 812=>x"2e00",
---- 813=>x"3100", 814=>x"3300", 815=>x"3700", 816=>x"2e00", 817=>x"2900", 818=>x"2c00", 819=>x"2f00",
---- 820=>x"3500", 821=>x"3300", 822=>x"3000", 823=>x"3600", 824=>x"2d00", 825=>x"2b00", 826=>x"3100",
---- 827=>x"3500", 828=>x"3700", 829=>x"3700", 830=>x"3200", 831=>x"3400", 832=>x"2a00", 833=>x"2e00",
---- 834=>x"3600", 835=>x"3700", 836=>x"3900", 837=>x"3400", 838=>x"3300", 839=>x"3600", 840=>x"2f00",
---- 841=>x"2f00", 842=>x"3300", 843=>x"3800", 844=>x"3900", 845=>x"3700", 846=>x"3700", 847=>x"3b00",
---- 848=>x"3100", 849=>x"3500", 850=>x"3500", 851=>x"3700", 852=>x"3a00", 853=>x"3a00", 854=>x"ca00",
---- 855=>x"3800", 856=>x"3600", 857=>x"3b00", 858=>x"3700", 859=>x"3600", 860=>x"3800", 861=>x"3d00",
---- 862=>x"3c00", 863=>x"3d00", 864=>x"2f00", 865=>x"3700", 866=>x"3700", 867=>x"3900", 868=>x"3700",
---- 869=>x"3600", 870=>x"3c00", 871=>x"3c00", 872=>x"3400", 873=>x"ca00", 874=>x"3900", 875=>x"3b00",
---- 876=>x"3800", 877=>x"4100", 878=>x"3e00", 879=>x"3d00", 880=>x"3300", 881=>x"3700", 882=>x"3900",
---- 883=>x"3800", 884=>x"3c00", 885=>x"3f00", 886=>x"3e00", 887=>x"3c00", 888=>x"3400", 889=>x"3700",
---- 890=>x"3700", 891=>x"3800", 892=>x"3b00", 893=>x"3c00", 894=>x"4200", 895=>x"3800", 896=>x"3700",
---- 897=>x"3700", 898=>x"3700", 899=>x"3900", 900=>x"3d00", 901=>x"3f00", 902=>x"3e00", 903=>x"3300",
---- 904=>x"3700", 905=>x"3800", 906=>x"3900", 907=>x"3c00", 908=>x"4100", 909=>x"4100", 910=>x"3b00",
---- 911=>x"cb00", 912=>x"3900", 913=>x"3b00", 914=>x"c400", 915=>x"3a00", 916=>x"4100", 917=>x"4000",
---- 918=>x"3700", 919=>x"3200", 920=>x"3b00", 921=>x"3a00", 922=>x"3c00", 923=>x"3d00", 924=>x"4100",
---- 925=>x"3f00", 926=>x"3800", 927=>x"2f00", 928=>x"3a00", 929=>x"3b00", 930=>x"3b00", 931=>x"3b00",
---- 932=>x"4200", 933=>x"3e00", 934=>x"3800", 935=>x"2f00", 936=>x"3b00", 937=>x"3900", 938=>x"3900",
---- 939=>x"3a00", 940=>x"3d00", 941=>x"3900", 942=>x"3700", 943=>x"3300", 944=>x"3e00", 945=>x"3d00",
---- 946=>x"3c00", 947=>x"3f00", 948=>x"3d00", 949=>x"3400", 950=>x"3000", 951=>x"3400", 952=>x"3a00",
---- 953=>x"3f00", 954=>x"4100", 955=>x"4000", 956=>x"3e00", 957=>x"3300", 958=>x"2c00", 959=>x"3000",
---- 960=>x"3c00", 961=>x"3c00", 962=>x"4300", 963=>x"3e00", 964=>x"3a00", 965=>x"3300", 966=>x"3100",
---- 967=>x"3500", 968=>x"3c00", 969=>x"3f00", 970=>x"3e00", 971=>x"3f00", 972=>x"3500", 973=>x"2e00",
---- 974=>x"3400", 975=>x"3500", 976=>x"3e00", 977=>x"4700", 978=>x"4a00", 979=>x"3b00", 980=>x"3400",
---- 981=>x"3000", 982=>x"3200", 983=>x"3000", 984=>x"3e00", 985=>x"4600", 986=>x"4300", 987=>x"3800",
---- 988=>x"3000", 989=>x"3000", 990=>x"3200", 991=>x"3300", 992=>x"3e00", 993=>x"4000", 994=>x"3900",
---- 995=>x"3600", 996=>x"3400", 997=>x"3000", 998=>x"3300", 999=>x"3300", 1000=>x"4200", 1001=>x"3e00",
---- 1002=>x"3800", 1003=>x"2f00", 1004=>x"3300", 1005=>x"3000", 1006=>x"2e00", 1007=>x"2f00", 1008=>x"4000",
---- 1009=>x"4200", 1010=>x"3700", 1011=>x"3100", 1012=>x"3000", 1013=>x"3300", 1014=>x"cb00", 1015=>x"3400",
---- 1016=>x"4100", 1017=>x"4100", 1018=>x"3500", 1019=>x"3100", 1020=>x"3200", 1021=>x"3500", 1022=>x"3400",
---- 1023=>x"3500", 1024=>x"4000", 1025=>x"3800", 1026=>x"3300", 1027=>x"3000", 1028=>x"3000", 1029=>x"3200",
---- 1030=>x"3200", 1031=>x"3600", 1032=>x"3f00", 1033=>x"3700", 1034=>x"3000", 1035=>x"3100", 1036=>x"3300",
---- 1037=>x"2f00", 1038=>x"3200", 1039=>x"ca00", 1040=>x"3d00", 1041=>x"3300", 1042=>x"2d00", 1043=>x"3000",
---- 1044=>x"3200", 1045=>x"3200", 1046=>x"3800", 1047=>x"3800", 1048=>x"3800", 1049=>x"3000", 1050=>x"2e00",
---- 1051=>x"3200", 1052=>x"3100", 1053=>x"3200", 1054=>x"3400", 1055=>x"3500", 1056=>x"3d00", 1057=>x"2e00",
---- 1058=>x"2e00", 1059=>x"3200", 1060=>x"3400", 1061=>x"3600", 1062=>x"3200", 1063=>x"2f00", 1064=>x"ca00",
---- 1065=>x"3000", 1066=>x"3000", 1067=>x"3400", 1068=>x"3000", 1069=>x"3500", 1070=>x"2f00", 1071=>x"2c00",
---- 1072=>x"3300", 1073=>x"2e00", 1074=>x"3200", 1075=>x"3200", 1076=>x"3400", 1077=>x"3300", 1078=>x"3100",
---- 1079=>x"3000", 1080=>x"3400", 1081=>x"3300", 1082=>x"3500", 1083=>x"3200", 1084=>x"3c00", 1085=>x"3600",
---- 1086=>x"2e00", 1087=>x"2d00", 1088=>x"3200", 1089=>x"3200", 1090=>x"3100", 1091=>x"2f00", 1092=>x"3600",
---- 1093=>x"3700", 1094=>x"3000", 1095=>x"2c00", 1096=>x"2b00", 1097=>x"2f00", 1098=>x"2d00", 1099=>x"2e00",
---- 1100=>x"3500", 1101=>x"3700", 1102=>x"2d00", 1103=>x"2d00", 1104=>x"2e00", 1105=>x"3100", 1106=>x"3000",
---- 1107=>x"2d00", 1108=>x"3b00", 1109=>x"3900", 1110=>x"2e00", 1111=>x"4300", 1112=>x"3000", 1113=>x"3400",
---- 1114=>x"2c00", 1115=>x"3200", 1116=>x"3b00", 1117=>x"3400", 1118=>x"3100", 1119=>x"4400", 1120=>x"2f00",
---- 1121=>x"2f00", 1122=>x"2900", 1123=>x"3c00", 1124=>x"3b00", 1125=>x"2e00", 1126=>x"2c00", 1127=>x"4800",
---- 1128=>x"3400", 1129=>x"3000", 1130=>x"2e00", 1131=>x"4100", 1132=>x"3800", 1133=>x"2900", 1134=>x"2b00",
---- 1135=>x"5000", 1136=>x"3300", 1137=>x"2d00", 1138=>x"3000", 1139=>x"c700", 1140=>x"3200", 1141=>x"2900",
---- 1142=>x"3000", 1143=>x"5f00", 1144=>x"3100", 1145=>x"2500", 1146=>x"3200", 1147=>x"3600", 1148=>x"2a00",
---- 1149=>x"2900", 1150=>x"3800", 1151=>x"6b00", 1152=>x"3200", 1153=>x"2c00", 1154=>x"3300", 1155=>x"3400",
---- 1156=>x"2d00", 1157=>x"2c00", 1158=>x"4600", 1159=>x"7700", 1160=>x"2f00", 1161=>x"2a00", 1162=>x"3700",
---- 1163=>x"3200", 1164=>x"2d00", 1165=>x"d100", 1166=>x"5900", 1167=>x"8300", 1168=>x"2e00", 1169=>x"2f00",
---- 1170=>x"3700", 1171=>x"2f00", 1172=>x"2c00", 1173=>x"3500", 1174=>x"6900", 1175=>x"8900", 1176=>x"2d00",
---- 1177=>x"3100", 1178=>x"3500", 1179=>x"2b00", 1180=>x"2800", 1181=>x"4000", 1182=>x"7400", 1183=>x"8b00",
---- 1184=>x"3700", 1185=>x"3200", 1186=>x"3300", 1187=>x"2d00", 1188=>x"2b00", 1189=>x"4b00", 1190=>x"7e00",
---- 1191=>x"8f00", 1192=>x"4000", 1193=>x"3600", 1194=>x"3200", 1195=>x"2b00", 1196=>x"2e00", 1197=>x"5a00",
---- 1198=>x"8300", 1199=>x"8d00", 1200=>x"3e00", 1201=>x"3b00", 1202=>x"3200", 1203=>x"2c00", 1204=>x"3800",
---- 1205=>x"6c00", 1206=>x"8a00", 1207=>x"8c00", 1208=>x"3c00", 1209=>x"3b00", 1210=>x"3300", 1211=>x"3100",
---- 1212=>x"ba00", 1213=>x"7800", 1214=>x"8c00", 1215=>x"8a00", 1216=>x"3800", 1217=>x"3700", 1218=>x"2f00",
---- 1219=>x"2b00", 1220=>x"5600", 1221=>x"8300", 1222=>x"8c00", 1223=>x"8900", 1224=>x"3a00", 1225=>x"3500",
---- 1226=>x"2b00", 1227=>x"3300", 1228=>x"6600", 1229=>x"8800", 1230=>x"8c00", 1231=>x"7600", 1232=>x"3600",
---- 1233=>x"2e00", 1234=>x"2700", 1235=>x"3f00", 1236=>x"7400", 1237=>x"8d00", 1238=>x"8c00", 1239=>x"8700",
---- 1240=>x"3000", 1241=>x"2c00", 1242=>x"2c00", 1243=>x"4d00", 1244=>x"7e00", 1245=>x"8e00", 1246=>x"8900",
---- 1247=>x"8900", 1248=>x"2b00", 1249=>x"2b00", 1250=>x"3700", 1251=>x"5a00", 1252=>x"8700", 1253=>x"8d00",
---- 1254=>x"8a00", 1255=>x"8a00", 1256=>x"2500", 1257=>x"2500", 1258=>x"4000", 1259=>x"6800", 1260=>x"8d00",
---- 1261=>x"8f00", 1262=>x"8a00", 1263=>x"8c00", 1264=>x"2400", 1265=>x"2700", 1266=>x"4c00", 1267=>x"7900",
---- 1268=>x"9100", 1269=>x"9200", 1270=>x"8e00", 1271=>x"9000", 1272=>x"2200", 1273=>x"2400", 1274=>x"5700",
---- 1275=>x"8600", 1276=>x"9100", 1277=>x"9200", 1278=>x"8b00", 1279=>x"9400", 1280=>x"2400", 1281=>x"2500",
---- 1282=>x"5c00", 1283=>x"8f00", 1284=>x"9200", 1285=>x"9000", 1286=>x"8d00", 1287=>x"9b00", 1288=>x"2a00",
---- 1289=>x"3200", 1290=>x"7000", 1291=>x"9100", 1292=>x"9400", 1293=>x"9000", 1294=>x"9000", 1295=>x"9d00",
---- 1296=>x"3300", 1297=>x"4500", 1298=>x"7d00", 1299=>x"9500", 1300=>x"9500", 1301=>x"8f00", 1302=>x"9400",
---- 1303=>x"9f00", 1304=>x"3000", 1305=>x"5d00", 1306=>x"8700", 1307=>x"9400", 1308=>x"9300", 1309=>x"9100",
---- 1310=>x"9500", 1311=>x"9f00", 1312=>x"2d00", 1313=>x"6d00", 1314=>x"8e00", 1315=>x"9500", 1316=>x"9200",
---- 1317=>x"8e00", 1318=>x"9a00", 1319=>x"9f00", 1320=>x"3400", 1321=>x"7a00", 1322=>x"9200", 1323=>x"9200",
---- 1324=>x"9200", 1325=>x"9200", 1326=>x"9c00", 1327=>x"9e00", 1328=>x"4900", 1329=>x"8200", 1330=>x"9400",
---- 1331=>x"9100", 1332=>x"9200", 1333=>x"9500", 1334=>x"9e00", 1335=>x"9c00", 1336=>x"5e00", 1337=>x"8800",
---- 1338=>x"9400", 1339=>x"9000", 1340=>x"9200", 1341=>x"9500", 1342=>x"9f00", 1343=>x"9d00", 1344=>x"6c00",
---- 1345=>x"8d00", 1346=>x"9500", 1347=>x"8d00", 1348=>x"9200", 1349=>x"9900", 1350=>x"9f00", 1351=>x"9b00",
---- 1352=>x"7900", 1353=>x"8e00", 1354=>x"9400", 1355=>x"9000", 1356=>x"9100", 1357=>x"9b00", 1358=>x"9e00",
---- 1359=>x"9900", 1360=>x"8500", 1361=>x"8d00", 1362=>x"9000", 1363=>x"9100", 1364=>x"9400", 1365=>x"9d00",
---- 1366=>x"9900", 1367=>x"9a00", 1368=>x"8a00", 1369=>x"8c00", 1370=>x"8f00", 1371=>x"9300", 1372=>x"9700",
---- 1373=>x"9c00", 1374=>x"9b00", 1375=>x"9b00", 1376=>x"8c00", 1377=>x"8c00", 1378=>x"9000", 1379=>x"9100",
---- 1380=>x"9500", 1381=>x"9c00", 1382=>x"9b00", 1383=>x"9900", 1384=>x"8f00", 1385=>x"9100", 1386=>x"9000",
---- 1387=>x"9000", 1388=>x"9700", 1389=>x"9d00", 1390=>x"9b00", 1391=>x"9b00", 1392=>x"9500", 1393=>x"9100",
---- 1394=>x"9300", 1395=>x"8e00", 1396=>x"9800", 1397=>x"9c00", 1398=>x"9a00", 1399=>x"9c00", 1400=>x"9200",
---- 1401=>x"9000", 1402=>x"9500", 1403=>x"9300", 1404=>x"9a00", 1405=>x"9b00", 1406=>x"9f00", 1407=>x"9b00",
---- 1408=>x"9500", 1409=>x"9300", 1410=>x"9600", 1411=>x"9300", 1412=>x"9a00", 1413=>x"9d00", 1414=>x"9d00",
---- 1415=>x"9a00", 1416=>x"9500", 1417=>x"9300", 1418=>x"9500", 1419=>x"9500", 1420=>x"9a00", 1421=>x"9a00",
---- 1422=>x"9a00", 1423=>x"9900", 1424=>x"9600", 1425=>x"9300", 1426=>x"9500", 1427=>x"9700", 1428=>x"9b00",
---- 1429=>x"9d00", 1430=>x"9c00", 1431=>x"9a00", 1432=>x"9a00", 1433=>x"9400", 1434=>x"9600", 1435=>x"9500",
---- 1436=>x"9c00", 1437=>x"9e00", 1438=>x"9c00", 1439=>x"9d00", 1440=>x"9900", 1441=>x"9600", 1442=>x"9500",
---- 1443=>x"9700", 1444=>x"9b00", 1445=>x"9c00", 1446=>x"9c00", 1447=>x"9c00", 1448=>x"9900", 1449=>x"9800",
---- 1450=>x"9700", 1451=>x"9a00", 1452=>x"9a00", 1453=>x"9c00", 1454=>x"9a00", 1455=>x"9b00", 1456=>x"9a00",
---- 1457=>x"9500", 1458=>x"9500", 1459=>x"9a00", 1460=>x"9b00", 1461=>x"9900", 1462=>x"6600", 1463=>x"9b00",
---- 1464=>x"9800", 1465=>x"9300", 1466=>x"9600", 1467=>x"9b00", 1468=>x"9a00", 1469=>x"9c00", 1470=>x"9800",
---- 1471=>x"9d00", 1472=>x"9900", 1473=>x"9100", 1474=>x"9900", 1475=>x"9900", 1476=>x"9b00", 1477=>x"9d00",
---- 1478=>x"9a00", 1479=>x"9b00", 1480=>x"9700", 1481=>x"8e00", 1482=>x"9c00", 1483=>x"9a00", 1484=>x"9c00",
---- 1485=>x"9c00", 1486=>x"9d00", 1487=>x"9d00", 1488=>x"9400", 1489=>x"9100", 1490=>x"9b00", 1491=>x"9d00",
---- 1492=>x"9e00", 1493=>x"9c00", 1494=>x"9c00", 1495=>x"9d00", 1496=>x"9200", 1497=>x"9300", 1498=>x"9800",
---- 1499=>x"9f00", 1500=>x"9e00", 1501=>x"9d00", 1502=>x"9900", 1503=>x"9c00", 1504=>x"9200", 1505=>x"9400",
---- 1506=>x"9700", 1507=>x"9f00", 1508=>x"9d00", 1509=>x"9c00", 1510=>x"9b00", 1511=>x"9a00", 1512=>x"9500",
---- 1513=>x"9100", 1514=>x"9a00", 1515=>x"9e00", 1516=>x"9d00", 1517=>x"9d00", 1518=>x"9c00", 1519=>x"9800",
---- 1520=>x"9700", 1521=>x"9200", 1522=>x"9700", 1523=>x"9700", 1524=>x"9a00", 1525=>x"9d00", 1526=>x"9a00",
---- 1527=>x"9800", 1528=>x"9400", 1529=>x"8d00", 1530=>x"8c00", 1531=>x"9000", 1532=>x"9300", 1533=>x"9300",
---- 1534=>x"9400", 1535=>x"9400", 1536=>x"8e00", 1537=>x"8100", 1538=>x"7e00", 1539=>x"8400", 1540=>x"8900",
---- 1541=>x"8b00", 1542=>x"8c00", 1543=>x"8d00", 1544=>x"8300", 1545=>x"7900", 1546=>x"7100", 1547=>x"7600",
---- 1548=>x"7c00", 1549=>x"8200", 1550=>x"8300", 1551=>x"8600", 1552=>x"7500", 1553=>x"7600", 1554=>x"6e00",
---- 1555=>x"6e00", 1556=>x"7300", 1557=>x"7a00", 1558=>x"7c00", 1559=>x"7c00", 1560=>x"7000", 1561=>x"7200",
---- 1562=>x"7200", 1563=>x"6900", 1564=>x"6f00", 1565=>x"6e00", 1566=>x"7500", 1567=>x"7600", 1568=>x"7200",
---- 1569=>x"7200", 1570=>x"7a00", 1571=>x"7200", 1572=>x"6d00", 1573=>x"7000", 1574=>x"6f00", 1575=>x"7200",
---- 1576=>x"7800", 1577=>x"7f00", 1578=>x"7f00", 1579=>x"8200", 1580=>x"7500", 1581=>x"7700", 1582=>x"7300",
---- 1583=>x"7300", 1584=>x"7c00", 1585=>x"8800", 1586=>x"8100", 1587=>x"8600", 1588=>x"8400", 1589=>x"7d00",
---- 1590=>x"7c00", 1591=>x"7a00", 1592=>x"8600", 1593=>x"8a00", 1594=>x"8400", 1595=>x"8700", 1596=>x"8e00",
---- 1597=>x"8100", 1598=>x"8000", 1599=>x"8000", 1600=>x"8e00", 1601=>x"8b00", 1602=>x"8a00", 1603=>x"8a00",
---- 1604=>x"8e00", 1605=>x"8a00", 1606=>x"8500", 1607=>x"8400", 1608=>x"9300", 1609=>x"8f00", 1610=>x"8d00",
---- 1611=>x"8c00", 1612=>x"8d00", 1613=>x"8e00", 1614=>x"8700", 1615=>x"8600", 1616=>x"9500", 1617=>x"9200",
---- 1618=>x"9100", 1619=>x"9100", 1620=>x"8e00", 1621=>x"8d00", 1622=>x"8900", 1623=>x"8b00", 1624=>x"9700",
---- 1625=>x"9400", 1626=>x"9100", 1627=>x"9200", 1628=>x"9100", 1629=>x"8e00", 1630=>x"8e00", 1631=>x"8d00",
---- 1632=>x"9500", 1633=>x"9400", 1634=>x"9200", 1635=>x"9100", 1636=>x"9200", 1637=>x"8f00", 1638=>x"8f00",
---- 1639=>x"8f00", 1640=>x"9500", 1641=>x"9700", 1642=>x"9100", 1643=>x"9100", 1644=>x"9100", 1645=>x"6f00",
---- 1646=>x"9200", 1647=>x"8f00", 1648=>x"6c00", 1649=>x"9600", 1650=>x"9300", 1651=>x"9100", 1652=>x"9100",
---- 1653=>x"8c00", 1654=>x"9000", 1655=>x"9100", 1656=>x"9600", 1657=>x"9600", 1658=>x"9400", 1659=>x"9200",
---- 1660=>x"9000", 1661=>x"8d00", 1662=>x"7100", 1663=>x"8e00", 1664=>x"9400", 1665=>x"9400", 1666=>x"9100",
---- 1667=>x"9000", 1668=>x"9200", 1669=>x"8f00", 1670=>x"9000", 1671=>x"8c00", 1672=>x"9200", 1673=>x"9300",
---- 1674=>x"9400", 1675=>x"9200", 1676=>x"9100", 1677=>x"8f00", 1678=>x"9100", 1679=>x"9200", 1680=>x"9300",
---- 1681=>x"9000", 1682=>x"9300", 1683=>x"9100", 1684=>x"9000", 1685=>x"9000", 1686=>x"9100", 1687=>x"9000",
---- 1688=>x"9200", 1689=>x"9300", 1690=>x"9100", 1691=>x"9100", 1692=>x"9000", 1693=>x"8d00", 1694=>x"9300",
---- 1695=>x"8e00", 1696=>x"9200", 1697=>x"9200", 1698=>x"9000", 1699=>x"9100", 1700=>x"9000", 1701=>x"8e00",
---- 1702=>x"9100", 1703=>x"8f00", 1704=>x"9300", 1705=>x"9400", 1706=>x"9100", 1707=>x"9200", 1708=>x"9000",
---- 1709=>x"9100", 1710=>x"9100", 1711=>x"8f00", 1712=>x"9500", 1713=>x"9900", 1714=>x"9100", 1715=>x"9100",
---- 1716=>x"9200", 1717=>x"9100", 1718=>x"9000", 1719=>x"9000", 1720=>x"9500", 1721=>x"9500", 1722=>x"9200",
---- 1723=>x"9200", 1724=>x"9200", 1725=>x"9200", 1726=>x"8f00", 1727=>x"8e00", 1728=>x"9200", 1729=>x"6c00",
---- 1730=>x"9100", 1731=>x"9300", 1732=>x"9300", 1733=>x"9100", 1734=>x"8f00", 1735=>x"8f00", 1736=>x"9200",
---- 1737=>x"9100", 1738=>x"9100", 1739=>x"8e00", 1740=>x"9200", 1741=>x"9100", 1742=>x"8f00", 1743=>x"8e00",
---- 1744=>x"9300", 1745=>x"9100", 1746=>x"8f00", 1747=>x"9000", 1748=>x"9100", 1749=>x"9000", 1750=>x"8e00",
---- 1751=>x"8d00", 1752=>x"9100", 1753=>x"9200", 1754=>x"9200", 1755=>x"9000", 1756=>x"6f00", 1757=>x"8e00",
---- 1758=>x"8b00", 1759=>x"8c00", 1760=>x"6e00", 1761=>x"9000", 1762=>x"9000", 1763=>x"8f00", 1764=>x"8e00",
---- 1765=>x"8c00", 1766=>x"8d00", 1767=>x"8c00", 1768=>x"8d00", 1769=>x"8f00", 1770=>x"8f00", 1771=>x"8d00",
---- 1772=>x"8d00", 1773=>x"8b00", 1774=>x"8c00", 1775=>x"8a00", 1776=>x"9000", 1777=>x"8e00", 1778=>x"8e00",
---- 1779=>x"8c00", 1780=>x"8d00", 1781=>x"8c00", 1782=>x"8c00", 1783=>x"8900", 1784=>x"8f00", 1785=>x"8f00",
---- 1786=>x"8f00", 1787=>x"8f00", 1788=>x"8e00", 1789=>x"8900", 1790=>x"8a00", 1791=>x"8b00", 1792=>x"8d00",
---- 1793=>x"9000", 1794=>x"8f00", 1795=>x"9000", 1796=>x"8e00", 1797=>x"8b00", 1798=>x"8a00", 1799=>x"8c00",
---- 1800=>x"9000", 1801=>x"8f00", 1802=>x"8e00", 1803=>x"8e00", 1804=>x"9300", 1805=>x"8c00", 1806=>x"8c00",
---- 1807=>x"8d00", 1808=>x"9000", 1809=>x"8e00", 1810=>x"8f00", 1811=>x"8f00", 1812=>x"8d00", 1813=>x"9000",
---- 1814=>x"9000", 1815=>x"8e00", 1816=>x"8e00", 1817=>x"9100", 1818=>x"9000", 1819=>x"9300", 1820=>x"9200",
---- 1821=>x"9300", 1822=>x"9100", 1823=>x"8f00", 1824=>x"8500", 1825=>x"8900", 1826=>x"8900", 1827=>x"8e00",
---- 1828=>x"9300", 1829=>x"9200", 1830=>x"9100", 1831=>x"9200", 1832=>x"7400", 1833=>x"7c00", 1834=>x"7e00",
---- 1835=>x"8400", 1836=>x"8900", 1837=>x"8c00", 1838=>x"9000", 1839=>x"9000", 1840=>x"6600", 1841=>x"6a00",
---- 1842=>x"7000", 1843=>x"7900", 1844=>x"7c00", 1845=>x"8000", 1846=>x"8400", 1847=>x"8a00", 1848=>x"5700",
---- 1849=>x"5d00", 1850=>x"6200", 1851=>x"6500", 1852=>x"6b00", 1853=>x"6f00", 1854=>x"7400", 1855=>x"7b00",
---- 1856=>x"4800", 1857=>x"4e00", 1858=>x"5500", 1859=>x"5300", 1860=>x"5c00", 1861=>x"6000", 1862=>x"6100",
---- 1863=>x"6a00", 1864=>x"b300", 1865=>x"4a00", 1866=>x"4d00", 1867=>x"4c00", 1868=>x"4f00", 1869=>x"5300",
---- 1870=>x"5200", 1871=>x"5200", 1872=>x"5400", 1873=>x"5200", 1874=>x"5200", 1875=>x"4c00", 1876=>x"4600",
---- 1877=>x"4600", 1878=>x"4300", 1879=>x"4200", 1880=>x"5a00", 1881=>x"5b00", 1882=>x"5700", 1883=>x"5300",
---- 1884=>x"5100", 1885=>x"4a00", 1886=>x"4400", 1887=>x"4100", 1888=>x"6400", 1889=>x"6100", 1890=>x"5e00",
---- 1891=>x"5900", 1892=>x"5900", 1893=>x"5100", 1894=>x"4b00", 1895=>x"4400", 1896=>x"6800", 1897=>x"6700",
---- 1898=>x"6500", 1899=>x"5f00", 1900=>x"5c00", 1901=>x"5700", 1902=>x"5200", 1903=>x"4d00", 1904=>x"9400",
---- 1905=>x"6b00", 1906=>x"6900", 1907=>x"6400", 1908=>x"6100", 1909=>x"6000", 1910=>x"5900", 1911=>x"5600",
---- 1912=>x"6900", 1913=>x"9200", 1914=>x"6b00", 1915=>x"6700", 1916=>x"6300", 1917=>x"6000", 1918=>x"5900",
---- 1919=>x"5b00", 1920=>x"6b00", 1921=>x"6b00", 1922=>x"6c00", 1923=>x"6900", 1924=>x"6500", 1925=>x"6200",
---- 1926=>x"5d00", 1927=>x"5d00", 1928=>x"6900", 1929=>x"7000", 1930=>x"6e00", 1931=>x"6800", 1932=>x"6700",
---- 1933=>x"6200", 1934=>x"6100", 1935=>x"5f00", 1936=>x"6500", 1937=>x"6b00", 1938=>x"6b00", 1939=>x"6900",
---- 1940=>x"6900", 1941=>x"6100", 1942=>x"5f00", 1943=>x"6300", 1944=>x"6300", 1945=>x"6600", 1946=>x"6800",
---- 1947=>x"6500", 1948=>x"6a00", 1949=>x"6500", 1950=>x"6000", 1951=>x"6300", 1952=>x"6200", 1953=>x"6500",
---- 1954=>x"6300", 1955=>x"6600", 1956=>x"6800", 1957=>x"6700", 1958=>x"6200", 1959=>x"6400", 1960=>x"5e00",
---- 1961=>x"6300", 1962=>x"6200", 1963=>x"6600", 1964=>x"6a00", 1965=>x"6900", 1966=>x"6500", 1967=>x"6800",
---- 1968=>x"5800", 1969=>x"5f00", 1970=>x"6200", 1971=>x"6200", 1972=>x"6800", 1973=>x"6b00", 1974=>x"6800",
---- 1975=>x"6c00", 1976=>x"5600", 1977=>x"5c00", 1978=>x"6100", 1979=>x"6300", 1980=>x"6600", 1981=>x"6b00",
---- 1982=>x"6b00", 1983=>x"6e00", 1984=>x"5600", 1985=>x"5800", 1986=>x"5f00", 1987=>x"6100", 1988=>x"6300",
---- 1989=>x"6a00", 1990=>x"6d00", 1991=>x"9000", 1992=>x"5500", 1993=>x"5a00", 1994=>x"5e00", 1995=>x"6300",
---- 1996=>x"6500", 1997=>x"6b00", 1998=>x"6f00", 1999=>x"6e00", 2000=>x"5300", 2001=>x"5600", 2002=>x"5c00",
---- 2003=>x"6400", 2004=>x"6a00", 2005=>x"6a00", 2006=>x"6d00", 2007=>x"6e00", 2008=>x"5100", 2009=>x"5400",
---- 2010=>x"5a00", 2011=>x"5f00", 2012=>x"5d00", 2013=>x"6700", 2014=>x"6d00", 2015=>x"6900", 2016=>x"4a00",
---- 2017=>x"5200", 2018=>x"5e00", 2019=>x"6500", 2020=>x"6500", 2021=>x"6600", 2022=>x"6400", 2023=>x"6b00",
---- 2024=>x"4600", 2025=>x"5200", 2026=>x"5500", 2027=>x"5800", 2028=>x"6000", 2029=>x"6500", 2030=>x"6400",
---- 2031=>x"6800", 2032=>x"4a00", 2033=>x"5600", 2034=>x"5800", 2035=>x"5e00", 2036=>x"5a00", 2037=>x"5b00",
---- 2038=>x"5f00", 2039=>x"6900", 2040=>x"6800", 2041=>x"6400", 2042=>x"5a00", 2043=>x"5c00", 2044=>x"5a00",
---- 2045=>x"5b00", 2046=>x"6000", 2047=>x"6400"),
---- 25 => (0=>x"9900", 1=>x"a100", 2=>x"bf00", 3=>x"cc00", 4=>x"d400", 5=>x"d500", 6=>x"da00", 7=>x"da00",
---- 8=>x"9a00", 9=>x"a100", 10=>x"c000", 11=>x"cd00", 12=>x"d300", 13=>x"d500", 14=>x"2500",
---- 15=>x"da00", 16=>x"9800", 17=>x"a000", 18=>x"be00", 19=>x"cc00", 20=>x"d200", 21=>x"d600",
---- 22=>x"d900", 23=>x"da00", 24=>x"9800", 25=>x"9800", 26=>x"ae00", 27=>x"c700", 28=>x"d000",
---- 29=>x"d600", 30=>x"d800", 31=>x"da00", 32=>x"9a00", 33=>x"9600", 34=>x"9c00", 35=>x"ba00",
---- 36=>x"cc00", 37=>x"d300", 38=>x"d500", 39=>x"d900", 40=>x"9a00", 41=>x"9800", 42=>x"9500",
---- 43=>x"a700", 44=>x"c300", 45=>x"cf00", 46=>x"d600", 47=>x"d700", 48=>x"9a00", 49=>x"9600",
---- 50=>x"9500", 51=>x"9900", 52=>x"b400", 53=>x"c800", 54=>x"d200", 55=>x"d600", 56=>x"9800",
---- 57=>x"9800", 58=>x"9700", 59=>x"9400", 60=>x"a100", 61=>x"c100", 62=>x"cc00", 63=>x"d400",
---- 64=>x"9800", 65=>x"9600", 66=>x"9400", 67=>x"9600", 68=>x"9600", 69=>x"b200", 70=>x"c900",
---- 71=>x"d200", 72=>x"9700", 73=>x"9800", 74=>x"9700", 75=>x"9400", 76=>x"9200", 77=>x"9c00",
---- 78=>x"bb00", 79=>x"ce00", 80=>x"9600", 81=>x"9700", 82=>x"9800", 83=>x"9600", 84=>x"9600",
---- 85=>x"9200", 86=>x"a800", 87=>x"c500", 88=>x"9800", 89=>x"9500", 90=>x"9600", 91=>x"9500",
---- 92=>x"9200", 93=>x"7100", 94=>x"9800", 95=>x"b700", 96=>x"9800", 97=>x"9500", 98=>x"9600",
---- 99=>x"9600", 100=>x"9500", 101=>x"9100", 102=>x"9100", 103=>x"a500", 104=>x"9800", 105=>x"9700",
---- 106=>x"9600", 107=>x"9700", 108=>x"9400", 109=>x"9300", 110=>x"9100", 111=>x"9600", 112=>x"9800",
---- 113=>x"9700", 114=>x"9800", 115=>x"9700", 116=>x"9400", 117=>x"9300", 118=>x"9200", 119=>x"9000",
---- 120=>x"9800", 121=>x"9900", 122=>x"9600", 123=>x"9600", 124=>x"9500", 125=>x"9200", 126=>x"9100",
---- 127=>x"9000", 128=>x"9a00", 129=>x"9b00", 130=>x"9800", 131=>x"9800", 132=>x"9600", 133=>x"9500",
---- 134=>x"9400", 135=>x"8d00", 136=>x"9b00", 137=>x"9900", 138=>x"9800", 139=>x"9900", 140=>x"9800",
---- 141=>x"9400", 142=>x"9400", 143=>x"8f00", 144=>x"9c00", 145=>x"9900", 146=>x"9700", 147=>x"9800",
---- 148=>x"9700", 149=>x"9500", 150=>x"9500", 151=>x"9100", 152=>x"9b00", 153=>x"9900", 154=>x"9500",
---- 155=>x"9400", 156=>x"9700", 157=>x"9400", 158=>x"9400", 159=>x"9100", 160=>x"9700", 161=>x"9900",
---- 162=>x"9600", 163=>x"9400", 164=>x"9500", 165=>x"9400", 166=>x"9100", 167=>x"6d00", 168=>x"6800",
---- 169=>x"9300", 170=>x"9500", 171=>x"9400", 172=>x"9200", 173=>x"9200", 174=>x"9100", 175=>x"8f00",
---- 176=>x"9500", 177=>x"9400", 178=>x"9000", 179=>x"8f00", 180=>x"9000", 181=>x"9000", 182=>x"8f00",
---- 183=>x"9000", 184=>x"9300", 185=>x"9500", 186=>x"9200", 187=>x"8f00", 188=>x"9100", 189=>x"9000",
---- 190=>x"8f00", 191=>x"8f00", 192=>x"9300", 193=>x"9100", 194=>x"9300", 195=>x"9000", 196=>x"9200",
---- 197=>x"9000", 198=>x"8e00", 199=>x"8e00", 200=>x"9200", 201=>x"8f00", 202=>x"8e00", 203=>x"8d00",
---- 204=>x"8f00", 205=>x"8f00", 206=>x"8b00", 207=>x"8e00", 208=>x"9200", 209=>x"8c00", 210=>x"8c00",
---- 211=>x"8e00", 212=>x"8d00", 213=>x"8d00", 214=>x"8c00", 215=>x"8e00", 216=>x"9300", 217=>x"9100",
---- 218=>x"8c00", 219=>x"7200", 220=>x"8e00", 221=>x"8b00", 222=>x"7200", 223=>x"8c00", 224=>x"9000",
---- 225=>x"8d00", 226=>x"8e00", 227=>x"8b00", 228=>x"8c00", 229=>x"8c00", 230=>x"8a00", 231=>x"8d00",
---- 232=>x"8f00", 233=>x"8e00", 234=>x"8d00", 235=>x"8e00", 236=>x"8b00", 237=>x"8d00", 238=>x"8a00",
---- 239=>x"8a00", 240=>x"8e00", 241=>x"8f00", 242=>x"8d00", 243=>x"8d00", 244=>x"8d00", 245=>x"8b00",
---- 246=>x"8d00", 247=>x"8d00", 248=>x"9000", 249=>x"8e00", 250=>x"9000", 251=>x"8e00", 252=>x"8d00",
---- 253=>x"8d00", 254=>x"8d00", 255=>x"8e00", 256=>x"9000", 257=>x"8f00", 258=>x"9100", 259=>x"8f00",
---- 260=>x"8d00", 261=>x"8b00", 262=>x"8d00", 263=>x"8e00", 264=>x"8d00", 265=>x"8f00", 266=>x"8e00",
---- 267=>x"8d00", 268=>x"8e00", 269=>x"8c00", 270=>x"8e00", 271=>x"8e00", 272=>x"8e00", 273=>x"9000",
---- 274=>x"8e00", 275=>x"9000", 276=>x"8d00", 277=>x"8d00", 278=>x"8c00", 279=>x"8f00", 280=>x"8e00",
---- 281=>x"8e00", 282=>x"8e00", 283=>x"8e00", 284=>x"8e00", 285=>x"8d00", 286=>x"8f00", 287=>x"8f00",
---- 288=>x"8f00", 289=>x"8f00", 290=>x"8f00", 291=>x"8c00", 292=>x"8e00", 293=>x"8f00", 294=>x"9000",
---- 295=>x"9000", 296=>x"8c00", 297=>x"9100", 298=>x"8d00", 299=>x"8c00", 300=>x"9000", 301=>x"8e00",
---- 302=>x"9000", 303=>x"9100", 304=>x"8d00", 305=>x"8e00", 306=>x"8f00", 307=>x"8f00", 308=>x"8f00",
---- 309=>x"9000", 310=>x"9100", 311=>x"9100", 312=>x"8f00", 313=>x"9100", 314=>x"8f00", 315=>x"8f00",
---- 316=>x"8f00", 317=>x"8f00", 318=>x"9000", 319=>x"9000", 320=>x"8f00", 321=>x"8f00", 322=>x"8f00",
---- 323=>x"9000", 324=>x"9000", 325=>x"9200", 326=>x"9000", 327=>x"9100", 328=>x"8c00", 329=>x"8f00",
---- 330=>x"9000", 331=>x"8f00", 332=>x"9000", 333=>x"9100", 334=>x"9100", 335=>x"9200", 336=>x"8e00",
---- 337=>x"8f00", 338=>x"9000", 339=>x"8e00", 340=>x"8e00", 341=>x"8f00", 342=>x"9200", 343=>x"9300",
---- 344=>x"8e00", 345=>x"8e00", 346=>x"9200", 347=>x"9200", 348=>x"8e00", 349=>x"8f00", 350=>x"9100",
---- 351=>x"9000", 352=>x"9000", 353=>x"8e00", 354=>x"9000", 355=>x"9000", 356=>x"9000", 357=>x"8f00",
---- 358=>x"8f00", 359=>x"9100", 360=>x"9100", 361=>x"8e00", 362=>x"8e00", 363=>x"8e00", 364=>x"9100",
---- 365=>x"9100", 366=>x"9100", 367=>x"6c00", 368=>x"8f00", 369=>x"8f00", 370=>x"9000", 371=>x"8e00",
---- 372=>x"8f00", 373=>x"8f00", 374=>x"9200", 375=>x"9000", 376=>x"8c00", 377=>x"8e00", 378=>x"8e00",
---- 379=>x"9000", 380=>x"9100", 381=>x"9000", 382=>x"8f00", 383=>x"9000", 384=>x"8e00", 385=>x"8e00",
---- 386=>x"8d00", 387=>x"8d00", 388=>x"8f00", 389=>x"9100", 390=>x"9000", 391=>x"9200", 392=>x"8f00",
---- 393=>x"8f00", 394=>x"8d00", 395=>x"8d00", 396=>x"8d00", 397=>x"9000", 398=>x"6e00", 399=>x"9100",
---- 400=>x"9000", 401=>x"8e00", 402=>x"8b00", 403=>x"8e00", 404=>x"8f00", 405=>x"8f00", 406=>x"9100",
---- 407=>x"9200", 408=>x"9100", 409=>x"8d00", 410=>x"8c00", 411=>x"8d00", 412=>x"8f00", 413=>x"8e00",
---- 414=>x"9400", 415=>x"9400", 416=>x"9000", 417=>x"8c00", 418=>x"8c00", 419=>x"8b00", 420=>x"8b00",
---- 421=>x"6f00", 422=>x"9200", 423=>x"9300", 424=>x"6c00", 425=>x"8e00", 426=>x"8c00", 427=>x"8a00",
---- 428=>x"8c00", 429=>x"9000", 430=>x"9300", 431=>x"6900", 432=>x"8f00", 433=>x"8700", 434=>x"8700",
---- 435=>x"8a00", 436=>x"8e00", 437=>x"8f00", 438=>x"9300", 439=>x"9500", 440=>x"9f00", 441=>x"a300",
---- 442=>x"9b00", 443=>x"8600", 444=>x"8900", 445=>x"9300", 446=>x"9700", 447=>x"9500", 448=>x"d700",
---- 449=>x"da00", 450=>x"ce00", 451=>x"a800", 452=>x"a500", 453=>x"c200", 454=>x"ae00", 455=>x"8e00",
---- 456=>x"d200", 457=>x"c900", 458=>x"c800", 459=>x"cd00", 460=>x"d500", 461=>x"d900", 462=>x"d700",
---- 463=>x"ac00", 464=>x"bd00", 465=>x"c600", 466=>x"cf00", 467=>x"d800", 468=>x"da00", 469=>x"da00",
---- 470=>x"dc00", 471=>x"d400", 472=>x"d000", 473=>x"da00", 474=>x"df00", 475=>x"e200", 476=>x"e500",
---- 477=>x"e900", 478=>x"df00", 479=>x"e300", 480=>x"db00", 481=>x"e100", 482=>x"e200", 483=>x"df00",
---- 484=>x"e000", 485=>x"e400", 486=>x"e800", 487=>x"ed00", 488=>x"da00", 489=>x"db00", 490=>x"da00",
---- 491=>x"d900", 492=>x"de00", 493=>x"de00", 494=>x"e200", 495=>x"eb00", 496=>x"d600", 497=>x"d500",
---- 498=>x"d700", 499=>x"d700", 500=>x"d300", 501=>x"d600", 502=>x"df00", 503=>x"e800", 504=>x"d200",
---- 505=>x"d300", 506=>x"d500", 507=>x"ce00", 508=>x"c900", 509=>x"d200", 510=>x"dc00", 511=>x"e600",
---- 512=>x"c800", 513=>x"cb00", 514=>x"ce00", 515=>x"cb00", 516=>x"d100", 517=>x"d700", 518=>x"dc00",
---- 519=>x"e200", 520=>x"c600", 521=>x"ca00", 522=>x"ca00", 523=>x"3100", 524=>x"d400", 525=>x"db00",
---- 526=>x"de00", 527=>x"e300", 528=>x"ca00", 529=>x"cc00", 530=>x"cd00", 531=>x"d300", 532=>x"d700",
---- 533=>x"d900", 534=>x"dd00", 535=>x"e100", 536=>x"cb00", 537=>x"cc00", 538=>x"cf00", 539=>x"d300",
---- 540=>x"d900", 541=>x"dc00", 542=>x"de00", 543=>x"e000", 544=>x"cb00", 545=>x"cf00", 546=>x"d300",
---- 547=>x"d500", 548=>x"2700", 549=>x"da00", 550=>x"de00", 551=>x"e100", 552=>x"ce00", 553=>x"d200",
---- 554=>x"d500", 555=>x"d700", 556=>x"d800", 557=>x"db00", 558=>x"dd00", 559=>x"e200", 560=>x"cd00",
---- 561=>x"d200", 562=>x"d500", 563=>x"d500", 564=>x"da00", 565=>x"de00", 566=>x"dc00", 567=>x"e500",
---- 568=>x"cb00", 569=>x"ce00", 570=>x"d200", 571=>x"d500", 572=>x"db00", 573=>x"dd00", 574=>x"dc00",
---- 575=>x"e600", 576=>x"c700", 577=>x"ce00", 578=>x"d100", 579=>x"d400", 580=>x"da00", 581=>x"de00",
---- 582=>x"dd00", 583=>x"e600", 584=>x"c700", 585=>x"d300", 586=>x"d300", 587=>x"d400", 588=>x"db00",
---- 589=>x"de00", 590=>x"e000", 591=>x"e000", 592=>x"c900", 593=>x"d000", 594=>x"d100", 595=>x"d300",
---- 596=>x"db00", 597=>x"de00", 598=>x"e100", 599=>x"ca00", 600=>x"c800", 601=>x"cd00", 602=>x"d200",
---- 603=>x"d200", 604=>x"d800", 605=>x"d800", 606=>x"df00", 607=>x"a400", 608=>x"be00", 609=>x"ca00",
---- 610=>x"d000", 611=>x"cd00", 612=>x"d700", 613=>x"d800", 614=>x"dc00", 615=>x"7500", 616=>x"bc00",
---- 617=>x"cc00", 618=>x"c100", 619=>x"c400", 620=>x"d300", 621=>x"d700", 622=>x"c900", 623=>x"4100",
---- 624=>x"be00", 625=>x"a400", 626=>x"a800", 627=>x"be00", 628=>x"cb00", 629=>x"db00", 630=>x"9700",
---- 631=>x"2400", 632=>x"9600", 633=>x"7b00", 634=>x"a700", 635=>x"bd00", 636=>x"c600", 637=>x"d500",
---- 638=>x"5900", 639=>x"2500", 640=>x"7a00", 641=>x"9600", 642=>x"ad00", 643=>x"ba00", 644=>x"d300",
---- 645=>x"b600", 646=>x"2d00", 647=>x"2600", 648=>x"9100", 649=>x"a600", 650=>x"b000", 651=>x"b600",
---- 652=>x"de00", 653=>x"8f00", 654=>x"1d00", 655=>x"2900", 656=>x"a900", 657=>x"a600", 658=>x"a900",
---- 659=>x"c600", 660=>x"dc00", 661=>x"5600", 662=>x"2000", 663=>x"2d00", 664=>x"9b00", 665=>x"9000",
---- 666=>x"ad00", 667=>x"df00", 668=>x"b900", 669=>x"3000", 670=>x"2600", 671=>x"2c00", 672=>x"7d00",
---- 673=>x"9d00", 674=>x"c300", 675=>x"e500", 676=>x"7d00", 677=>x"1d00", 678=>x"2900", 679=>x"2a00",
---- 680=>x"8200", 681=>x"b100", 682=>x"d900", 683=>x"d600", 684=>x"4b00", 685=>x"1f00", 686=>x"d900",
---- 687=>x"2c00", 688=>x"9f00", 689=>x"c700", 690=>x"e700", 691=>x"a900", 692=>x"2500", 693=>x"2200",
---- 694=>x"2300", 695=>x"2a00", 696=>x"c400", 697=>x"d900", 698=>x"e000", 699=>x"6300", 700=>x"1c00",
---- 701=>x"2700", 702=>x"2600", 703=>x"2b00", 704=>x"2d00", 705=>x"e300", 706=>x"a300", 707=>x"2600",
---- 708=>x"2300", 709=>x"2c00", 710=>x"2e00", 711=>x"2e00", 712=>x"d700", 713=>x"cb00", 714=>x"4300",
---- 715=>x"2100", 716=>x"2700", 717=>x"d500", 718=>x"3200", 719=>x"3100", 720=>x"e300", 721=>x"7f00",
---- 722=>x"2a00", 723=>x"2a00", 724=>x"2a00", 725=>x"2f00", 726=>x"3000", 727=>x"3300", 728=>x"a100",
---- 729=>x"3000", 730=>x"3300", 731=>x"2b00", 732=>x"2b00", 733=>x"3100", 734=>x"3400", 735=>x"3200",
---- 736=>x"3300", 737=>x"2300", 738=>x"2800", 739=>x"2a00", 740=>x"3100", 741=>x"3400", 742=>x"3300",
---- 743=>x"3000", 744=>x"2900", 745=>x"d500", 746=>x"2d00", 747=>x"3000", 748=>x"3400", 749=>x"3200",
---- 750=>x"3000", 751=>x"2c00", 752=>x"2e00", 753=>x"2e00", 754=>x"2d00", 755=>x"3300", 756=>x"3300",
---- 757=>x"3500", 758=>x"2f00", 759=>x"2e00", 760=>x"3000", 761=>x"2f00", 762=>x"3400", 763=>x"3600",
---- 764=>x"3700", 765=>x"3500", 766=>x"2e00", 767=>x"2c00", 768=>x"2f00", 769=>x"3400", 770=>x"3800",
---- 771=>x"3500", 772=>x"3600", 773=>x"3800", 774=>x"2f00", 775=>x"2f00", 776=>x"3700", 777=>x"3b00",
---- 778=>x"3800", 779=>x"3400", 780=>x"3200", 781=>x"3000", 782=>x"3100", 783=>x"3200", 784=>x"3500",
---- 785=>x"3700", 786=>x"3600", 787=>x"3300", 788=>x"c700", 789=>x"3100", 790=>x"2d00", 791=>x"2d00",
---- 792=>x"3500", 793=>x"3400", 794=>x"3600", 795=>x"3400", 796=>x"3700", 797=>x"3100", 798=>x"2c00",
---- 799=>x"2f00", 800=>x"3500", 801=>x"3700", 802=>x"3500", 803=>x"3700", 804=>x"3500", 805=>x"3100",
---- 806=>x"2e00", 807=>x"2e00", 808=>x"3800", 809=>x"3900", 810=>x"3f00", 811=>x"3600", 812=>x"3300",
---- 813=>x"3200", 814=>x"2e00", 815=>x"2c00", 816=>x"3800", 817=>x"3b00", 818=>x"3700", 819=>x"2f00",
---- 820=>x"2c00", 821=>x"3000", 822=>x"2c00", 823=>x"2c00", 824=>x"3700", 825=>x"3800", 826=>x"3700",
---- 827=>x"3100", 828=>x"2e00", 829=>x"2e00", 830=>x"2f00", 831=>x"2e00", 832=>x"3600", 833=>x"3700",
---- 834=>x"3500", 835=>x"d000", 836=>x"2b00", 837=>x"2f00", 838=>x"2d00", 839=>x"3100", 840=>x"3700",
---- 841=>x"3a00", 842=>x"3300", 843=>x"2a00", 844=>x"2900", 845=>x"2f00", 846=>x"3000", 847=>x"3400",
---- 848=>x"3800", 849=>x"3500", 850=>x"3000", 851=>x"2900", 852=>x"2900", 853=>x"3000", 854=>x"3600",
---- 855=>x"3700", 856=>x"3900", 857=>x"3000", 858=>x"3000", 859=>x"2c00", 860=>x"2900", 861=>x"2c00",
---- 862=>x"3200", 863=>x"3500", 864=>x"3600", 865=>x"2f00", 866=>x"3500", 867=>x"2d00", 868=>x"2900",
---- 869=>x"2c00", 870=>x"3300", 871=>x"3300", 872=>x"3700", 873=>x"2f00", 874=>x"2d00", 875=>x"2e00",
---- 876=>x"2d00", 877=>x"3300", 878=>x"3400", 879=>x"d300", 880=>x"3200", 881=>x"3000", 882=>x"2e00",
---- 883=>x"2a00", 884=>x"2e00", 885=>x"3400", 886=>x"3100", 887=>x"2f00", 888=>x"2e00", 889=>x"2c00",
---- 890=>x"2d00", 891=>x"2d00", 892=>x"2e00", 893=>x"3600", 894=>x"2e00", 895=>x"3000", 896=>x"2f00",
---- 897=>x"2d00", 898=>x"2d00", 899=>x"2f00", 900=>x"3400", 901=>x"3600", 902=>x"2b00", 903=>x"2c00",
---- 904=>x"2e00", 905=>x"2c00", 906=>x"3000", 907=>x"3300", 908=>x"3800", 909=>x"3700", 910=>x"2d00",
---- 911=>x"2a00", 912=>x"2e00", 913=>x"d300", 914=>x"3000", 915=>x"3300", 916=>x"3700", 917=>x"3300",
---- 918=>x"2a00", 919=>x"2d00", 920=>x"2f00", 921=>x"2e00", 922=>x"2e00", 923=>x"3300", 924=>x"3500",
---- 925=>x"2e00", 926=>x"2b00", 927=>x"3a00", 928=>x"2e00", 929=>x"3300", 930=>x"3200", 931=>x"3600",
---- 932=>x"3900", 933=>x"2e00", 934=>x"2a00", 935=>x"4700", 936=>x"2d00", 937=>x"2e00", 938=>x"3700",
---- 939=>x"3700", 940=>x"3000", 941=>x"2b00", 942=>x"2d00", 943=>x"5600", 944=>x"3300", 945=>x"3300",
---- 946=>x"3800", 947=>x"3300", 948=>x"2a00", 949=>x"2c00", 950=>x"4300", 951=>x"6e00", 952=>x"3300",
---- 953=>x"3600", 954=>x"3600", 955=>x"3200", 956=>x"2a00", 957=>x"3100", 958=>x"5700", 959=>x"7e00",
---- 960=>x"3000", 961=>x"3400", 962=>x"3500", 963=>x"2e00", 964=>x"2b00", 965=>x"3600", 966=>x"6300",
---- 967=>x"8600", 968=>x"3300", 969=>x"3900", 970=>x"3400", 971=>x"2c00", 972=>x"3100", 973=>x"4b00",
---- 974=>x"7000", 975=>x"8900", 976=>x"3400", 977=>x"3800", 978=>x"3100", 979=>x"2d00", 980=>x"3400",
---- 981=>x"5800", 982=>x"7f00", 983=>x"8b00", 984=>x"3400", 985=>x"3600", 986=>x"2f00", 987=>x"2d00",
---- 988=>x"c200", 989=>x"6400", 990=>x"8500", 991=>x"8d00", 992=>x"3900", 993=>x"3400", 994=>x"3000",
---- 995=>x"2c00", 996=>x"4500", 997=>x"7000", 998=>x"8900", 999=>x"8a00", 1000=>x"3900", 1001=>x"3800",
---- 1002=>x"3300", 1003=>x"3000", 1004=>x"4e00", 1005=>x"7f00", 1006=>x"8e00", 1007=>x"8600", 1008=>x"3800",
---- 1009=>x"3a00", 1010=>x"3700", 1011=>x"3600", 1012=>x"5b00", 1013=>x"8400", 1014=>x"8d00", 1015=>x"8400",
---- 1016=>x"3600", 1017=>x"3100", 1018=>x"3700", 1019=>x"4400", 1020=>x"6c00", 1021=>x"8900", 1022=>x"8b00",
---- 1023=>x"8200", 1024=>x"3400", 1025=>x"2b00", 1026=>x"3200", 1027=>x"5000", 1028=>x"7d00", 1029=>x"8d00",
---- 1030=>x"8900", 1031=>x"7f00", 1032=>x"3400", 1033=>x"2800", 1034=>x"2c00", 1035=>x"5a00", 1036=>x"8700",
---- 1037=>x"8d00", 1038=>x"8600", 1039=>x"8100", 1040=>x"3400", 1041=>x"2700", 1042=>x"2e00", 1043=>x"6500",
---- 1044=>x"8e00", 1045=>x"8c00", 1046=>x"8500", 1047=>x"8600", 1048=>x"3100", 1049=>x"2c00", 1050=>x"4200",
---- 1051=>x"7700", 1052=>x"8e00", 1053=>x"8d00", 1054=>x"8700", 1055=>x"8b00", 1056=>x"2d00", 1057=>x"3100",
---- 1058=>x"5900", 1059=>x"8300", 1060=>x"9100", 1061=>x"8e00", 1062=>x"8700", 1063=>x"9100", 1064=>x"cd00",
---- 1065=>x"4000", 1066=>x"6900", 1067=>x"8c00", 1068=>x"8e00", 1069=>x"8b00", 1070=>x"8900", 1071=>x"9500",
---- 1072=>x"3300", 1073=>x"4800", 1074=>x"7800", 1075=>x"8e00", 1076=>x"8e00", 1077=>x"8800", 1078=>x"8a00",
---- 1079=>x"9600", 1080=>x"2e00", 1081=>x"5400", 1082=>x"8400", 1083=>x"9100", 1084=>x"8c00", 1085=>x"8900",
---- 1086=>x"8f00", 1087=>x"9a00", 1088=>x"3200", 1089=>x"6400", 1090=>x"8800", 1091=>x"8d00", 1092=>x"8a00",
---- 1093=>x"8a00", 1094=>x"9400", 1095=>x"a100", 1096=>x"4100", 1097=>x"7100", 1098=>x"8c00", 1099=>x"8b00",
---- 1100=>x"8700", 1101=>x"8b00", 1102=>x"9800", 1103=>x"9f00", 1104=>x"5f00", 1105=>x"7900", 1106=>x"8d00",
---- 1107=>x"8800", 1108=>x"8600", 1109=>x"8d00", 1110=>x"9c00", 1111=>x"9f00", 1112=>x"6a00", 1113=>x"8500",
---- 1114=>x"8a00", 1115=>x"8500", 1116=>x"8700", 1117=>x"9200", 1118=>x"a000", 1119=>x"a000", 1120=>x"7900",
---- 1121=>x"8b00", 1122=>x"8800", 1123=>x"8300", 1124=>x"8900", 1125=>x"9b00", 1126=>x"a000", 1127=>x"9d00",
---- 1128=>x"8100", 1129=>x"8900", 1130=>x"8500", 1131=>x"8100", 1132=>x"8d00", 1133=>x"9d00", 1134=>x"9e00",
---- 1135=>x"9d00", 1136=>x"8700", 1137=>x"8b00", 1138=>x"8500", 1139=>x"8500", 1140=>x"9100", 1141=>x"9c00",
---- 1142=>x"9d00", 1143=>x"9b00", 1144=>x"8700", 1145=>x"8700", 1146=>x"7b00", 1147=>x"8800", 1148=>x"9800",
---- 1149=>x"9d00", 1150=>x"9c00", 1151=>x"9c00", 1152=>x"8b00", 1153=>x"8800", 1154=>x"8400", 1155=>x"8b00",
---- 1156=>x"9c00", 1157=>x"9f00", 1158=>x"9e00", 1159=>x"9b00", 1160=>x"8d00", 1161=>x"8600", 1162=>x"8400",
---- 1163=>x"9300", 1164=>x"a000", 1165=>x"9e00", 1166=>x"9c00", 1167=>x"9b00", 1168=>x"8b00", 1169=>x"8500",
---- 1170=>x"8600", 1171=>x"9900", 1172=>x"9f00", 1173=>x"9e00", 1174=>x"9b00", 1175=>x"9b00", 1176=>x"8b00",
---- 1177=>x"8600", 1178=>x"8a00", 1179=>x"9b00", 1180=>x"a100", 1181=>x"a000", 1182=>x"9d00", 1183=>x"9c00",
---- 1184=>x"8c00", 1185=>x"8800", 1186=>x"9200", 1187=>x"9f00", 1188=>x"a100", 1189=>x"9d00", 1190=>x"9a00",
---- 1191=>x"9900", 1192=>x"8900", 1193=>x"8900", 1194=>x"9800", 1195=>x"a200", 1196=>x"a100", 1197=>x"9d00",
---- 1198=>x"9b00", 1199=>x"9800", 1200=>x"8900", 1201=>x"9000", 1202=>x"a300", 1203=>x"a700", 1204=>x"a000",
---- 1205=>x"9c00", 1206=>x"9c00", 1207=>x"9a00", 1208=>x"8500", 1209=>x"9200", 1210=>x"ae00", 1211=>x"ac00",
---- 1212=>x"9c00", 1213=>x"9d00", 1214=>x"9c00", 1215=>x"9a00", 1216=>x"8800", 1217=>x"9a00", 1218=>x"a000",
---- 1219=>x"a200", 1220=>x"9e00", 1221=>x"9c00", 1222=>x"9c00", 1223=>x"9a00", 1224=>x"8c00", 1225=>x"9e00",
---- 1226=>x"a200", 1227=>x"a000", 1228=>x"5e00", 1229=>x"9d00", 1230=>x"9c00", 1231=>x"9a00", 1232=>x"9100",
---- 1233=>x"a000", 1234=>x"a000", 1235=>x"9e00", 1236=>x"9d00", 1237=>x"9c00", 1238=>x"9a00", 1239=>x"9900",
---- 1240=>x"9700", 1241=>x"a000", 1242=>x"9f00", 1243=>x"9f00", 1244=>x"9e00", 1245=>x"9c00", 1246=>x"9500",
---- 1247=>x"9800", 1248=>x"9b00", 1249=>x"a000", 1250=>x"9d00", 1251=>x"9d00", 1252=>x"9d00", 1253=>x"9b00",
---- 1254=>x"9600", 1255=>x"9800", 1256=>x"9e00", 1257=>x"a100", 1258=>x"9c00", 1259=>x"9d00", 1260=>x"9b00",
---- 1261=>x"9800", 1262=>x"9b00", 1263=>x"9800", 1264=>x"a000", 1265=>x"9f00", 1266=>x"9c00", 1267=>x"9a00",
---- 1268=>x"9a00", 1269=>x"9a00", 1270=>x"9800", 1271=>x"9500", 1272=>x"a100", 1273=>x"9d00", 1274=>x"9c00",
---- 1275=>x"9c00", 1276=>x"9b00", 1277=>x"9b00", 1278=>x"9700", 1279=>x"9600", 1280=>x"a000", 1281=>x"9e00",
---- 1282=>x"9c00", 1283=>x"9a00", 1284=>x"9800", 1285=>x"9900", 1286=>x"9900", 1287=>x"9600", 1288=>x"a000",
---- 1289=>x"9d00", 1290=>x"9c00", 1291=>x"9a00", 1292=>x"9a00", 1293=>x"9900", 1294=>x"9600", 1295=>x"9500",
---- 1296=>x"9d00", 1297=>x"9d00", 1298=>x"9900", 1299=>x"9900", 1300=>x"9900", 1301=>x"9500", 1302=>x"9600",
---- 1303=>x"9700", 1304=>x"9d00", 1305=>x"9d00", 1306=>x"9b00", 1307=>x"9900", 1308=>x"9600", 1309=>x"9500",
---- 1310=>x"9700", 1311=>x"9600", 1312=>x"9e00", 1313=>x"9b00", 1314=>x"9900", 1315=>x"9b00", 1316=>x"9900",
---- 1317=>x"9600", 1318=>x"9800", 1319=>x"9700", 1320=>x"9b00", 1321=>x"9b00", 1322=>x"9b00", 1323=>x"9a00",
---- 1324=>x"9700", 1325=>x"9900", 1326=>x"9800", 1327=>x"9700", 1328=>x"9a00", 1329=>x"9900", 1330=>x"9a00",
---- 1331=>x"9a00", 1332=>x"9700", 1333=>x"9700", 1334=>x"9900", 1335=>x"9500", 1336=>x"9c00", 1337=>x"9b00",
---- 1338=>x"6500", 1339=>x"6600", 1340=>x"6900", 1341=>x"9600", 1342=>x"9700", 1343=>x"9800", 1344=>x"9900",
---- 1345=>x"9900", 1346=>x"9900", 1347=>x"9800", 1348=>x"9600", 1349=>x"9900", 1350=>x"9600", 1351=>x"9600",
---- 1352=>x"9a00", 1353=>x"9b00", 1354=>x"9700", 1355=>x"9800", 1356=>x"9600", 1357=>x"9600", 1358=>x"9600",
---- 1359=>x"9300", 1360=>x"9a00", 1361=>x"9a00", 1362=>x"9800", 1363=>x"9800", 1364=>x"9800", 1365=>x"9500",
---- 1366=>x"9400", 1367=>x"9800", 1368=>x"9b00", 1369=>x"9a00", 1370=>x"9800", 1371=>x"9800", 1372=>x"9800",
---- 1373=>x"9400", 1374=>x"9400", 1375=>x"9600", 1376=>x"9b00", 1377=>x"9900", 1378=>x"9800", 1379=>x"9700",
---- 1380=>x"9700", 1381=>x"9600", 1382=>x"9200", 1383=>x"6b00", 1384=>x"9a00", 1385=>x"9900", 1386=>x"9500",
---- 1387=>x"9700", 1388=>x"9600", 1389=>x"9400", 1390=>x"9300", 1391=>x"9200", 1392=>x"9900", 1393=>x"9600",
---- 1394=>x"9800", 1395=>x"9500", 1396=>x"9500", 1397=>x"9400", 1398=>x"9400", 1399=>x"9200", 1400=>x"9600",
---- 1401=>x"9800", 1402=>x"9900", 1403=>x"9800", 1404=>x"9700", 1405=>x"9600", 1406=>x"9500", 1407=>x"9300",
---- 1408=>x"9900", 1409=>x"9800", 1410=>x"9700", 1411=>x"9700", 1412=>x"9800", 1413=>x"9600", 1414=>x"9700",
---- 1415=>x"9400", 1416=>x"9700", 1417=>x"9800", 1418=>x"9a00", 1419=>x"9700", 1420=>x"9800", 1421=>x"9600",
---- 1422=>x"9a00", 1423=>x"6b00", 1424=>x"9600", 1425=>x"9800", 1426=>x"9a00", 1427=>x"9700", 1428=>x"9a00",
---- 1429=>x"9800", 1430=>x"9800", 1431=>x"9500", 1432=>x"9b00", 1433=>x"9c00", 1434=>x"9900", 1435=>x"9800",
---- 1436=>x"9800", 1437=>x"9900", 1438=>x"9500", 1439=>x"9900", 1440=>x"9900", 1441=>x"9a00", 1442=>x"9a00",
---- 1443=>x"9900", 1444=>x"9a00", 1445=>x"9800", 1446=>x"9900", 1447=>x"9800", 1448=>x"9900", 1449=>x"9700",
---- 1450=>x"9a00", 1451=>x"9a00", 1452=>x"9b00", 1453=>x"9800", 1454=>x"9600", 1455=>x"9700", 1456=>x"9900",
---- 1457=>x"9900", 1458=>x"9b00", 1459=>x"9900", 1460=>x"9b00", 1461=>x"9900", 1462=>x"9700", 1463=>x"9a00",
---- 1464=>x"9a00", 1465=>x"9b00", 1466=>x"9b00", 1467=>x"9800", 1468=>x"9c00", 1469=>x"9900", 1470=>x"9c00",
---- 1471=>x"9d00", 1472=>x"9a00", 1473=>x"6600", 1474=>x"9b00", 1475=>x"9a00", 1476=>x"9a00", 1477=>x"9a00",
---- 1478=>x"9b00", 1479=>x"9a00", 1480=>x"9900", 1481=>x"9700", 1482=>x"9c00", 1483=>x"9800", 1484=>x"9900",
---- 1485=>x"9800", 1486=>x"9700", 1487=>x"9800", 1488=>x"9a00", 1489=>x"9800", 1490=>x"9c00", 1491=>x"9700",
---- 1492=>x"9600", 1493=>x"9800", 1494=>x"9500", 1495=>x"9800", 1496=>x"9a00", 1497=>x"9a00", 1498=>x"9a00",
---- 1499=>x"9700", 1500=>x"9800", 1501=>x"9900", 1502=>x"9600", 1503=>x"9800", 1504=>x"9500", 1505=>x"9800",
---- 1506=>x"9700", 1507=>x"9600", 1508=>x"9600", 1509=>x"9500", 1510=>x"9500", 1511=>x"9700", 1512=>x"9500",
---- 1513=>x"9600", 1514=>x"9800", 1515=>x"9700", 1516=>x"9700", 1517=>x"9600", 1518=>x"9800", 1519=>x"6b00",
---- 1520=>x"9200", 1521=>x"9500", 1522=>x"9800", 1523=>x"9800", 1524=>x"9700", 1525=>x"9700", 1526=>x"9500",
---- 1527=>x"9400", 1528=>x"9500", 1529=>x"9800", 1530=>x"9400", 1531=>x"9600", 1532=>x"9600", 1533=>x"9600",
---- 1534=>x"9500", 1535=>x"9400", 1536=>x"9200", 1537=>x"9300", 1538=>x"9200", 1539=>x"9600", 1540=>x"9700",
---- 1541=>x"9400", 1542=>x"9800", 1543=>x"9500", 1544=>x"8900", 1545=>x"8b00", 1546=>x"8b00", 1547=>x"8c00",
---- 1548=>x"6e00", 1549=>x"9300", 1550=>x"9200", 1551=>x"9300", 1552=>x"7b00", 1553=>x"8400", 1554=>x"8100",
---- 1555=>x"8100", 1556=>x"8800", 1557=>x"8c00", 1558=>x"8c00", 1559=>x"8b00", 1560=>x"7500", 1561=>x"7a00",
---- 1562=>x"7500", 1563=>x"7a00", 1564=>x"7c00", 1565=>x"7d00", 1566=>x"8100", 1567=>x"8500", 1568=>x"7200",
---- 1569=>x"7100", 1570=>x"7200", 1571=>x"7400", 1572=>x"7200", 1573=>x"7500", 1574=>x"7600", 1575=>x"7600",
---- 1576=>x"7100", 1577=>x"6e00", 1578=>x"7000", 1579=>x"6f00", 1580=>x"6d00", 1581=>x"6d00", 1582=>x"6d00",
---- 1583=>x"6d00", 1584=>x"7500", 1585=>x"7100", 1586=>x"6f00", 1587=>x"6c00", 1588=>x"6a00", 1589=>x"6900",
---- 1590=>x"6b00", 1591=>x"6800", 1592=>x"7a00", 1593=>x"7b00", 1594=>x"7700", 1595=>x"7100", 1596=>x"6f00",
---- 1597=>x"6b00", 1598=>x"6900", 1599=>x"6500", 1600=>x"7c00", 1601=>x"8000", 1602=>x"7f00", 1603=>x"8500",
---- 1604=>x"7a00", 1605=>x"7400", 1606=>x"9300", 1607=>x"6b00", 1608=>x"8600", 1609=>x"8600", 1610=>x"8200",
---- 1611=>x"8300", 1612=>x"8000", 1613=>x"7b00", 1614=>x"7a00", 1615=>x"7500", 1616=>x"8800", 1617=>x"8900",
---- 1618=>x"8900", 1619=>x"8900", 1620=>x"8600", 1621=>x"8000", 1622=>x"7e00", 1623=>x"7900", 1624=>x"8b00",
---- 1625=>x"8a00", 1626=>x"8a00", 1627=>x"8700", 1628=>x"8800", 1629=>x"8500", 1630=>x"8200", 1631=>x"7f00",
---- 1632=>x"8e00", 1633=>x"8e00", 1634=>x"8c00", 1635=>x"8800", 1636=>x"8800", 1637=>x"8700", 1638=>x"8700",
---- 1639=>x"8200", 1640=>x"9000", 1641=>x"8f00", 1642=>x"8c00", 1643=>x"8b00", 1644=>x"8900", 1645=>x"8700",
---- 1646=>x"8a00", 1647=>x"8800", 1648=>x"8e00", 1649=>x"8d00", 1650=>x"8e00", 1651=>x"8d00", 1652=>x"8b00",
---- 1653=>x"8a00", 1654=>x"8900", 1655=>x"8900", 1656=>x"8f00", 1657=>x"8f00", 1658=>x"8e00", 1659=>x"8d00",
---- 1660=>x"8d00", 1661=>x"8a00", 1662=>x"8a00", 1663=>x"8600", 1664=>x"8c00", 1665=>x"8e00", 1666=>x"8d00",
---- 1667=>x"8d00", 1668=>x"8d00", 1669=>x"8c00", 1670=>x"8d00", 1671=>x"8700", 1672=>x"8f00", 1673=>x"9000",
---- 1674=>x"8f00", 1675=>x"8f00", 1676=>x"8d00", 1677=>x"8d00", 1678=>x"8b00", 1679=>x"8b00", 1680=>x"8d00",
---- 1681=>x"8f00", 1682=>x"8d00", 1683=>x"8c00", 1684=>x"8d00", 1685=>x"8b00", 1686=>x"8a00", 1687=>x"8a00",
---- 1688=>x"8a00", 1689=>x"8c00", 1690=>x"8d00", 1691=>x"8a00", 1692=>x"8d00", 1693=>x"8a00", 1694=>x"7300",
---- 1695=>x"8a00", 1696=>x"8b00", 1697=>x"8b00", 1698=>x"8d00", 1699=>x"8d00", 1700=>x"8a00", 1701=>x"8600",
---- 1702=>x"8900", 1703=>x"8b00", 1704=>x"8e00", 1705=>x"8d00", 1706=>x"8d00", 1707=>x"8b00", 1708=>x"8900",
---- 1709=>x"8800", 1710=>x"8600", 1711=>x"8900", 1712=>x"8f00", 1713=>x"8f00", 1714=>x"8a00", 1715=>x"8b00",
---- 1716=>x"8a00", 1717=>x"8800", 1718=>x"8700", 1719=>x"8600", 1720=>x"8e00", 1721=>x"8d00", 1722=>x"8b00",
---- 1723=>x"8a00", 1724=>x"8400", 1725=>x"8400", 1726=>x"8500", 1727=>x"8600", 1728=>x"8b00", 1729=>x"8c00",
---- 1730=>x"8c00", 1731=>x"8800", 1732=>x"8500", 1733=>x"8500", 1734=>x"8700", 1735=>x"8400", 1736=>x"8a00",
---- 1737=>x"8b00", 1738=>x"8c00", 1739=>x"8a00", 1740=>x"8900", 1741=>x"8600", 1742=>x"8500", 1743=>x"8500",
---- 1744=>x"8c00", 1745=>x"8d00", 1746=>x"8900", 1747=>x"8b00", 1748=>x"8700", 1749=>x"8400", 1750=>x"8700",
---- 1751=>x"8600", 1752=>x"8a00", 1753=>x"8d00", 1754=>x"8d00", 1755=>x"8900", 1756=>x"8900", 1757=>x"8500",
---- 1758=>x"8300", 1759=>x"8400", 1760=>x"8a00", 1761=>x"8c00", 1762=>x"8d00", 1763=>x"8a00", 1764=>x"8900",
---- 1765=>x"8700", 1766=>x"8500", 1767=>x"8400", 1768=>x"8b00", 1769=>x"8c00", 1770=>x"8a00", 1771=>x"8a00",
---- 1772=>x"8900", 1773=>x"8700", 1774=>x"8800", 1775=>x"8200", 1776=>x"8b00", 1777=>x"8e00", 1778=>x"8b00",
---- 1779=>x"8c00", 1780=>x"8d00", 1781=>x"8700", 1782=>x"8800", 1783=>x"8100", 1784=>x"8a00", 1785=>x"8b00",
---- 1786=>x"8c00", 1787=>x"8b00", 1788=>x"8a00", 1789=>x"8600", 1790=>x"8800", 1791=>x"8700", 1792=>x"8a00",
---- 1793=>x"8b00", 1794=>x"8d00", 1795=>x"8a00", 1796=>x"8a00", 1797=>x"8a00", 1798=>x"8600", 1799=>x"8300",
---- 1800=>x"8c00", 1801=>x"8c00", 1802=>x"8f00", 1803=>x"8b00", 1804=>x"8900", 1805=>x"8800", 1806=>x"8500",
---- 1807=>x"8200", 1808=>x"8d00", 1809=>x"8f00", 1810=>x"8d00", 1811=>x"8b00", 1812=>x"8c00", 1813=>x"8b00",
---- 1814=>x"8800", 1815=>x"8500", 1816=>x"8e00", 1817=>x"8e00", 1818=>x"8f00", 1819=>x"8d00", 1820=>x"8a00",
---- 1821=>x"8800", 1822=>x"8800", 1823=>x"8400", 1824=>x"8f00", 1825=>x"9000", 1826=>x"8f00", 1827=>x"9000",
---- 1828=>x"8e00", 1829=>x"8b00", 1830=>x"8b00", 1831=>x"8800", 1832=>x"9100", 1833=>x"9200", 1834=>x"9000",
---- 1835=>x"8f00", 1836=>x"8d00", 1837=>x"8c00", 1838=>x"8b00", 1839=>x"8c00", 1840=>x"8b00", 1841=>x"8e00",
---- 1842=>x"8e00", 1843=>x"8b00", 1844=>x"8c00", 1845=>x"8e00", 1846=>x"8e00", 1847=>x"8b00", 1848=>x"7b00",
---- 1849=>x"8000", 1850=>x"8600", 1851=>x"8500", 1852=>x"8800", 1853=>x"8a00", 1854=>x"8c00", 1855=>x"8e00",
---- 1856=>x"6800", 1857=>x"6b00", 1858=>x"7400", 1859=>x"7600", 1860=>x"7900", 1861=>x"7c00", 1862=>x"8600",
---- 1863=>x"8900", 1864=>x"5500", 1865=>x"5900", 1866=>x"5d00", 1867=>x"6200", 1868=>x"6500", 1869=>x"6900",
---- 1870=>x"7300", 1871=>x"7c00", 1872=>x"4700", 1873=>x"4800", 1874=>x"4a00", 1875=>x"4900", 1876=>x"4f00",
---- 1877=>x"4d00", 1878=>x"5a00", 1879=>x"6700", 1880=>x"3e00", 1881=>x"3900", 1882=>x"3800", 1883=>x"3700",
---- 1884=>x"3300", 1885=>x"3500", 1886=>x"3d00", 1887=>x"4800", 1888=>x"3f00", 1889=>x"3900", 1890=>x"3500",
---- 1891=>x"3100", 1892=>x"2b00", 1893=>x"2f00", 1894=>x"2900", 1895=>x"3000", 1896=>x"b500", 1897=>x"3e00",
---- 1898=>x"3700", 1899=>x"3300", 1900=>x"2e00", 1901=>x"2900", 1902=>x"2300", 1903=>x"2700", 1904=>x"5000",
---- 1905=>x"4700", 1906=>x"3f00", 1907=>x"3600", 1908=>x"2d00", 1909=>x"2d00", 1910=>x"2800", 1911=>x"2600",
---- 1912=>x"5400", 1913=>x"4d00", 1914=>x"4900", 1915=>x"4100", 1916=>x"3900", 1917=>x"2f00", 1918=>x"2a00",
---- 1919=>x"2900", 1920=>x"5500", 1921=>x"5100", 1922=>x"5200", 1923=>x"4600", 1924=>x"4200", 1925=>x"3600",
---- 1926=>x"2e00", 1927=>x"2e00", 1928=>x"5b00", 1929=>x"5800", 1930=>x"5200", 1931=>x"4b00", 1932=>x"4800",
---- 1933=>x"4200", 1934=>x"3c00", 1935=>x"3800", 1936=>x"5f00", 1937=>x"5e00", 1938=>x"5500", 1939=>x"4f00",
---- 1940=>x"5100", 1941=>x"4b00", 1942=>x"4a00", 1943=>x"4d00", 1944=>x"9e00", 1945=>x"6200", 1946=>x"5c00",
---- 1947=>x"5500", 1948=>x"5400", 1949=>x"5400", 1950=>x"5700", 1951=>x"5900", 1952=>x"6200", 1953=>x"6600",
---- 1954=>x"5f00", 1955=>x"5900", 1956=>x"5800", 1957=>x"5e00", 1958=>x"5f00", 1959=>x"5e00", 1960=>x"6700",
---- 1961=>x"6500", 1962=>x"6100", 1963=>x"6000", 1964=>x"6500", 1965=>x"6600", 1966=>x"6a00", 1967=>x"6600",
---- 1968=>x"6800", 1969=>x"6400", 1970=>x"6400", 1971=>x"6400", 1972=>x"6800", 1973=>x"6d00", 1974=>x"6f00",
---- 1975=>x"6f00", 1976=>x"6d00", 1977=>x"6700", 1978=>x"6700", 1979=>x"6900", 1980=>x"7000", 1981=>x"7400",
---- 1982=>x"7400", 1983=>x"7100", 1984=>x"6e00", 1985=>x"6b00", 1986=>x"6a00", 1987=>x"7000", 1988=>x"7500",
---- 1989=>x"7400", 1990=>x"7400", 1991=>x"7200", 1992=>x"6d00", 1993=>x"7100", 1994=>x"7300", 1995=>x"7500",
---- 1996=>x"7600", 1997=>x"7900", 1998=>x"7600", 1999=>x"7200", 2000=>x"6f00", 2001=>x"7300", 2002=>x"7900",
---- 2003=>x"7800", 2004=>x"7600", 2005=>x"7700", 2006=>x"7200", 2007=>x"7300", 2008=>x"6e00", 2009=>x"7500",
---- 2010=>x"7800", 2011=>x"7800", 2012=>x"7c00", 2013=>x"7300", 2014=>x"7600", 2015=>x"7400", 2016=>x"7000",
---- 2017=>x"7500", 2018=>x"7600", 2019=>x"7800", 2020=>x"7600", 2021=>x"7900", 2022=>x"8700", 2023=>x"7500",
---- 2024=>x"6e00", 2025=>x"7300", 2026=>x"7600", 2027=>x"7500", 2028=>x"7700", 2029=>x"7c00", 2030=>x"7c00",
---- 2031=>x"7a00", 2032=>x"6d00", 2033=>x"7200", 2034=>x"7100", 2035=>x"7300", 2036=>x"7d00", 2037=>x"8200",
---- 2038=>x"7f00", 2039=>x"7b00", 2040=>x"6900", 2041=>x"6700", 2042=>x"7400", 2043=>x"7d00", 2044=>x"8200",
---- 2045=>x"8700", 2046=>x"8300", 2047=>x"7d00"),
---- 26 => (0=>x"da00", 1=>x"d300", 2=>x"c000", 3=>x"9600", 4=>x"6c00", 5=>x"6500", 6=>x"6900", 7=>x"6c00",
---- 8=>x"da00", 9=>x"d300", 10=>x"c000", 11=>x"9500", 12=>x"6a00", 13=>x"6600", 14=>x"6900",
---- 15=>x"6c00", 16=>x"db00", 17=>x"d400", 18=>x"c100", 19=>x"9800", 20=>x"6c00", 21=>x"6500",
---- 22=>x"9600", 23=>x"6d00", 24=>x"db00", 25=>x"d900", 26=>x"ce00", 27=>x"b100", 28=>x"7f00",
---- 29=>x"6400", 30=>x"6600", 31=>x"6c00", 32=>x"d900", 33=>x"d900", 34=>x"2a00", 35=>x"c200",
---- 36=>x"9d00", 37=>x"6f00", 38=>x"6700", 39=>x"6b00", 40=>x"d900", 41=>x"db00", 42=>x"d900",
---- 43=>x"d000", 44=>x"b600", 45=>x"8900", 46=>x"6800", 47=>x"6700", 48=>x"db00", 49=>x"db00",
---- 50=>x"da00", 51=>x"d800", 52=>x"c800", 53=>x"a600", 54=>x"8a00", 55=>x"6700", 56=>x"d800",
---- 57=>x"d900", 58=>x"db00", 59=>x"db00", 60=>x"d300", 61=>x"c000", 62=>x"9400", 63=>x"6a00",
---- 64=>x"d800", 65=>x"d900", 66=>x"dc00", 67=>x"dc00", 68=>x"d900", 69=>x"ce00", 70=>x"b300",
---- 71=>x"8000", 72=>x"d500", 73=>x"d900", 74=>x"da00", 75=>x"db00", 76=>x"db00", 77=>x"d600",
---- 78=>x"c400", 79=>x"9c00", 80=>x"d000", 81=>x"d600", 82=>x"d900", 83=>x"dc00", 84=>x"dc00",
---- 85=>x"da00", 86=>x"d100", 87=>x"b900", 88=>x"cc00", 89=>x"d300", 90=>x"d700", 91=>x"d900",
---- 92=>x"db00", 93=>x"de00", 94=>x"da00", 95=>x"c900", 96=>x"c300", 97=>x"cf00", 98=>x"d600",
---- 99=>x"d800", 100=>x"db00", 101=>x"dc00", 102=>x"db00", 103=>x"d300", 104=>x"b500", 105=>x"cc00",
---- 106=>x"d300", 107=>x"d700", 108=>x"da00", 109=>x"dc00", 110=>x"de00", 111=>x"d900", 112=>x"a100",
---- 113=>x"c200", 114=>x"d000", 115=>x"d700", 116=>x"2600", 117=>x"db00", 118=>x"dd00", 119=>x"de00",
---- 120=>x"9000", 121=>x"b000", 122=>x"ca00", 123=>x"d200", 124=>x"d800", 125=>x"da00", 126=>x"dd00",
---- 127=>x"de00", 128=>x"8a00", 129=>x"9800", 130=>x"b800", 131=>x"3700", 132=>x"cf00", 133=>x"d600",
---- 134=>x"2400", 135=>x"2200", 136=>x"8c00", 137=>x"8f00", 138=>x"aa00", 139=>x"c800", 140=>x"d200",
---- 141=>x"d700", 142=>x"db00", 143=>x"df00", 144=>x"9000", 145=>x"8e00", 146=>x"9700", 147=>x"b900",
---- 148=>x"ce00", 149=>x"d700", 150=>x"db00", 151=>x"dd00", 152=>x"8e00", 153=>x"8d00", 154=>x"8c00",
---- 155=>x"a300", 156=>x"c600", 157=>x"d200", 158=>x"d800", 159=>x"dd00", 160=>x"8f00", 161=>x"8e00",
---- 162=>x"8c00", 163=>x"9200", 164=>x"b700", 165=>x"ce00", 166=>x"d600", 167=>x"db00", 168=>x"8e00",
---- 169=>x"8c00", 170=>x"8c00", 171=>x"8b00", 172=>x"a200", 173=>x"c500", 174=>x"d200", 175=>x"d900",
---- 176=>x"8d00", 177=>x"8e00", 178=>x"8c00", 179=>x"8e00", 180=>x"9100", 181=>x"b400", 182=>x"ce00",
---- 183=>x"d500", 184=>x"8e00", 185=>x"9000", 186=>x"9000", 187=>x"8e00", 188=>x"8c00", 189=>x"9e00",
---- 190=>x"c200", 191=>x"d000", 192=>x"8f00", 193=>x"8e00", 194=>x"8f00", 195=>x"8c00", 196=>x"8e00",
---- 197=>x"9200", 198=>x"ae00", 199=>x"cb00", 200=>x"8e00", 201=>x"8b00", 202=>x"8d00", 203=>x"8c00",
---- 204=>x"8e00", 205=>x"8f00", 206=>x"9a00", 207=>x"bc00", 208=>x"8c00", 209=>x"8e00", 210=>x"8e00",
---- 211=>x"8c00", 212=>x"8c00", 213=>x"8d00", 214=>x"8f00", 215=>x"a700", 216=>x"8d00", 217=>x"8c00",
---- 218=>x"8e00", 219=>x"8d00", 220=>x"8b00", 221=>x"8d00", 222=>x"8a00", 223=>x"8d00", 224=>x"8d00",
---- 225=>x"8e00", 226=>x"8e00", 227=>x"8c00", 228=>x"8b00", 229=>x"8d00", 230=>x"8a00", 231=>x"8700",
---- 232=>x"8b00", 233=>x"8a00", 234=>x"8e00", 235=>x"8c00", 236=>x"8d00", 237=>x"8d00", 238=>x"8b00",
---- 239=>x"8800", 240=>x"8d00", 241=>x"8c00", 242=>x"8d00", 243=>x"8e00", 244=>x"8e00", 245=>x"8f00",
---- 246=>x"8d00", 247=>x"8a00", 248=>x"8e00", 249=>x"8e00", 250=>x"8f00", 251=>x"8e00", 252=>x"9000",
---- 253=>x"8f00", 254=>x"8c00", 255=>x"8c00", 256=>x"8a00", 257=>x"8b00", 258=>x"9200", 259=>x"9000",
---- 260=>x"9000", 261=>x"9100", 262=>x"8e00", 263=>x"8d00", 264=>x"8c00", 265=>x"8d00", 266=>x"9000",
---- 267=>x"9100", 268=>x"8f00", 269=>x"8f00", 270=>x"9100", 271=>x"8e00", 272=>x"8e00", 273=>x"8f00",
---- 274=>x"8f00", 275=>x"9200", 276=>x"7200", 277=>x"8f00", 278=>x"9100", 279=>x"9100", 280=>x"9000",
---- 281=>x"9000", 282=>x"8e00", 283=>x"9000", 284=>x"9100", 285=>x"9000", 286=>x"6e00", 287=>x"9200",
---- 288=>x"9100", 289=>x"9000", 290=>x"6f00", 291=>x"9000", 292=>x"9200", 293=>x"9200", 294=>x"9400",
---- 295=>x"9500", 296=>x"9000", 297=>x"9000", 298=>x"9100", 299=>x"9400", 300=>x"9200", 301=>x"9100",
---- 302=>x"9600", 303=>x"9400", 304=>x"9000", 305=>x"9200", 306=>x"9200", 307=>x"9300", 308=>x"9000",
---- 309=>x"9200", 310=>x"9400", 311=>x"9700", 312=>x"9000", 313=>x"8c00", 314=>x"9300", 315=>x"9100",
---- 316=>x"9100", 317=>x"9600", 318=>x"9500", 319=>x"9800", 320=>x"8f00", 321=>x"9000", 322=>x"6c00",
---- 323=>x"9000", 324=>x"9400", 325=>x"9400", 326=>x"9600", 327=>x"9400", 328=>x"9200", 329=>x"9100",
---- 330=>x"9100", 331=>x"9400", 332=>x"9300", 333=>x"9400", 334=>x"9400", 335=>x"9a00", 336=>x"9000",
---- 337=>x"9100", 338=>x"9100", 339=>x"9200", 340=>x"9400", 341=>x"9500", 342=>x"9600", 343=>x"9c00",
---- 344=>x"8e00", 345=>x"8f00", 346=>x"9000", 347=>x"9100", 348=>x"9300", 349=>x"9600", 350=>x"9a00",
---- 351=>x"9d00", 352=>x"8d00", 353=>x"8f00", 354=>x"9000", 355=>x"9100", 356=>x"9400", 357=>x"9600",
---- 358=>x"9c00", 359=>x"9900", 360=>x"9000", 361=>x"9200", 362=>x"9400", 363=>x"9300", 364=>x"9700",
---- 365=>x"9b00", 366=>x"9900", 367=>x"7e00", 368=>x"9100", 369=>x"9100", 370=>x"9300", 371=>x"9600",
---- 372=>x"9900", 373=>x"a000", 374=>x"8f00", 375=>x"5600", 376=>x"9100", 377=>x"9100", 378=>x"9300",
---- 379=>x"9500", 380=>x"9b00", 381=>x"9a00", 382=>x"7400", 383=>x"3500", 384=>x"9200", 385=>x"9300",
---- 386=>x"9700", 387=>x"9900", 388=>x"6400", 389=>x"8400", 390=>x"4a00", 391=>x"2e00", 392=>x"9200",
---- 393=>x"9600", 394=>x"9a00", 395=>x"9a00", 396=>x"8f00", 397=>x"6200", 398=>x"2c00", 399=>x"2900",
---- 400=>x"9300", 401=>x"6800", 402=>x"9b00", 403=>x"9700", 404=>x"7300", 405=>x"3800", 406=>x"2600",
---- 407=>x"2900", 408=>x"9500", 409=>x"9b00", 410=>x"9900", 411=>x"8700", 412=>x"4900", 413=>x"2900",
---- 414=>x"2500", 415=>x"2800", 416=>x"9800", 417=>x"9a00", 418=>x"9200", 419=>x"6200", 420=>x"2d00",
---- 421=>x"2a00", 422=>x"2900", 423=>x"2e00", 424=>x"9900", 425=>x"9700", 426=>x"7500", 427=>x"3c00",
---- 428=>x"2800", 429=>x"2c00", 430=>x"2800", 431=>x"2a00", 432=>x"9b00", 433=>x"8b00", 434=>x"4d00",
---- 435=>x"2900", 436=>x"2b00", 437=>x"2b00", 438=>x"2b00", 439=>x"2c00", 440=>x"9200", 441=>x"6200",
---- 442=>x"3000", 443=>x"2a00", 444=>x"2b00", 445=>x"2d00", 446=>x"2c00", 447=>x"2f00", 448=>x"7400",
---- 449=>x"3a00", 450=>x"2900", 451=>x"2a00", 452=>x"2d00", 453=>x"3000", 454=>x"3200", 455=>x"2f00",
---- 456=>x"b600", 457=>x"2900", 458=>x"2b00", 459=>x"2d00", 460=>x"2a00", 461=>x"3500", 462=>x"2d00",
---- 463=>x"3100", 464=>x"5b00", 465=>x"1d00", 466=>x"2c00", 467=>x"2d00", 468=>x"2d00", 469=>x"2f00",
---- 470=>x"2e00", 471=>x"3100", 472=>x"9100", 473=>x"2000", 474=>x"2b00", 475=>x"2c00", 476=>x"2f00",
---- 477=>x"2e00", 478=>x"3100", 479=>x"3a00", 480=>x"c600", 481=>x"3800", 482=>x"2700", 483=>x"2c00",
---- 484=>x"2e00", 485=>x"2d00", 486=>x"2f00", 487=>x"3400", 488=>x"de00", 489=>x"5700", 490=>x"2200",
---- 491=>x"2c00", 492=>x"2c00", 493=>x"2e00", 494=>x"3200", 495=>x"3200", 496=>x"e400", 497=>x"7700",
---- 498=>x"2300", 499=>x"2c00", 500=>x"2c00", 501=>x"d000", 502=>x"3200", 503=>x"3400", 504=>x"eb00",
---- 505=>x"7500", 506=>x"2200", 507=>x"2c00", 508=>x"2b00", 509=>x"2c00", 510=>x"2e00", 511=>x"3200",
---- 512=>x"ec00", 513=>x"8800", 514=>x"1f00", 515=>x"2a00", 516=>x"2c00", 517=>x"2e00", 518=>x"3400",
---- 519=>x"3700", 520=>x"e900", 521=>x"8600", 522=>x"1c00", 523=>x"2900", 524=>x"2e00", 525=>x"3100",
---- 526=>x"3500", 527=>x"3c00", 528=>x"e400", 529=>x"7b00", 530=>x"2000", 531=>x"2d00", 532=>x"2f00",
---- 533=>x"3200", 534=>x"3300", 535=>x"3600", 536=>x"e200", 537=>x"6800", 538=>x"2500", 539=>x"2a00",
---- 540=>x"2d00", 541=>x"3000", 542=>x"2f00", 543=>x"3100", 544=>x"d800", 545=>x"4c00", 546=>x"2700",
---- 547=>x"3000", 548=>x"3100", 549=>x"3400", 550=>x"2f00", 551=>x"3100", 552=>x"c700", 553=>x"3a00",
---- 554=>x"2600", 555=>x"2c00", 556=>x"3300", 557=>x"3200", 558=>x"3200", 559=>x"2e00", 560=>x"b100",
---- 561=>x"2c00", 562=>x"d400", 563=>x"3300", 564=>x"3600", 565=>x"3300", 566=>x"3400", 567=>x"3200",
---- 568=>x"9400", 569=>x"2700", 570=>x"3100", 571=>x"3100", 572=>x"3300", 573=>x"3500", 574=>x"3500",
---- 575=>x"3300", 576=>x"7d00", 577=>x"2000", 578=>x"3100", 579=>x"3300", 580=>x"3300", 581=>x"3800",
---- 582=>x"3300", 583=>x"3300", 584=>x"5d00", 585=>x"1e00", 586=>x"2f00", 587=>x"2c00", 588=>x"2e00",
---- 589=>x"2e00", 590=>x"3100", 591=>x"3900", 592=>x"3c00", 593=>x"2100", 594=>x"2c00", 595=>x"2b00",
---- 596=>x"3200", 597=>x"2d00", 598=>x"2e00", 599=>x"3400", 600=>x"2800", 601=>x"2400", 602=>x"2c00",
---- 603=>x"2e00", 604=>x"2e00", 605=>x"3000", 606=>x"3100", 607=>x"3400", 608=>x"2300", 609=>x"2800",
---- 610=>x"2b00", 611=>x"2a00", 612=>x"2c00", 613=>x"3300", 614=>x"3100", 615=>x"3800", 616=>x"2500",
---- 617=>x"2b00", 618=>x"2b00", 619=>x"2d00", 620=>x"3000", 621=>x"3200", 622=>x"2e00", 623=>x"3400",
---- 624=>x"2a00", 625=>x"3400", 626=>x"3500", 627=>x"3100", 628=>x"2f00", 629=>x"3500", 630=>x"3500",
---- 631=>x"3300", 632=>x"2800", 633=>x"3300", 634=>x"3b00", 635=>x"3200", 636=>x"3500", 637=>x"3500",
---- 638=>x"3200", 639=>x"2d00", 640=>x"2800", 641=>x"2800", 642=>x"3100", 643=>x"3a00", 644=>x"4200",
---- 645=>x"3100", 646=>x"2d00", 647=>x"2800", 648=>x"2800", 649=>x"2a00", 650=>x"3200", 651=>x"3400",
---- 652=>x"3400", 653=>x"d100", 654=>x"2b00", 655=>x"2a00", 656=>x"2b00", 657=>x"2c00", 658=>x"3000",
---- 659=>x"3100", 660=>x"3100", 661=>x"3800", 662=>x"2900", 663=>x"2900", 664=>x"3100", 665=>x"2f00",
---- 666=>x"3000", 667=>x"3200", 668=>x"3000", 669=>x"2e00", 670=>x"3400", 671=>x"3300", 672=>x"2f00",
---- 673=>x"3500", 674=>x"3500", 675=>x"3100", 676=>x"3a00", 677=>x"3000", 678=>x"3700", 679=>x"4200",
---- 680=>x"3100", 681=>x"3600", 682=>x"3700", 683=>x"3100", 684=>x"3400", 685=>x"3000", 686=>x"3100",
---- 687=>x"4200", 688=>x"2f00", 689=>x"2e00", 690=>x"3000", 691=>x"2d00", 692=>x"2e00", 693=>x"2d00",
---- 694=>x"3300", 695=>x"3a00", 696=>x"3100", 697=>x"3100", 698=>x"3200", 699=>x"2c00", 700=>x"2c00",
---- 701=>x"3200", 702=>x"3500", 703=>x"3800", 704=>x"3000", 705=>x"2f00", 706=>x"3200", 707=>x"2b00",
---- 708=>x"2a00", 709=>x"3100", 710=>x"3600", 711=>x"3800", 712=>x"2f00", 713=>x"3000", 714=>x"2e00",
---- 715=>x"2a00", 716=>x"2b00", 717=>x"3100", 718=>x"3800", 719=>x"3300", 720=>x"3000", 721=>x"3000",
---- 722=>x"2d00", 723=>x"3100", 724=>x"3300", 725=>x"3600", 726=>x"3600", 727=>x"2e00", 728=>x"3400",
---- 729=>x"3300", 730=>x"3100", 731=>x"2a00", 732=>x"3300", 733=>x"3900", 734=>x"2f00", 735=>x"2d00",
---- 736=>x"3000", 737=>x"3200", 738=>x"3400", 739=>x"3200", 740=>x"3700", 741=>x"3900", 742=>x"2f00",
---- 743=>x"2800", 744=>x"3000", 745=>x"2b00", 746=>x"3100", 747=>x"3300", 748=>x"3800", 749=>x"3700",
---- 750=>x"3100", 751=>x"2c00", 752=>x"2e00", 753=>x"2d00", 754=>x"3200", 755=>x"3500", 756=>x"3c00",
---- 757=>x"3c00", 758=>x"3300", 759=>x"3000", 760=>x"2c00", 761=>x"2b00", 762=>x"3300", 763=>x"3b00",
---- 764=>x"3700", 765=>x"3d00", 766=>x"3c00", 767=>x"3400", 768=>x"2a00", 769=>x"2a00", 770=>x"3400",
---- 771=>x"4000", 772=>x"3e00", 773=>x"3500", 774=>x"3200", 775=>x"3f00", 776=>x"3200", 777=>x"2e00",
---- 778=>x"3600", 779=>x"3500", 780=>x"2a00", 781=>x"2e00", 782=>x"2f00", 783=>x"5200", 784=>x"3000",
---- 785=>x"3300", 786=>x"3600", 787=>x"3500", 788=>x"2b00", 789=>x"3100", 790=>x"3500", 791=>x"6800",
---- 792=>x"2f00", 793=>x"3400", 794=>x"3600", 795=>x"3400", 796=>x"3300", 797=>x"3200", 798=>x"4900",
---- 799=>x"7900", 800=>x"3100", 801=>x"3400", 802=>x"3300", 803=>x"3100", 804=>x"3300", 805=>x"3800",
---- 806=>x"6000", 807=>x"8400", 808=>x"3000", 809=>x"3300", 810=>x"3500", 811=>x"2f00", 812=>x"3400",
---- 813=>x"4500", 814=>x"6b00", 815=>x"8700", 816=>x"ce00", 817=>x"3500", 818=>x"3400", 819=>x"3600",
---- 820=>x"4200", 821=>x"5000", 822=>x"7800", 823=>x"8a00", 824=>x"3700", 825=>x"3900", 826=>x"3200",
---- 827=>x"3b00", 828=>x"4700", 829=>x"6200", 830=>x"8200", 831=>x"8900", 832=>x"3800", 833=>x"3300",
---- 834=>x"3400", 835=>x"3d00", 836=>x"4c00", 837=>x"7400", 838=>x"8600", 839=>x"8500", 840=>x"3600",
---- 841=>x"2f00", 842=>x"3600", 843=>x"4400", 844=>x"5900", 845=>x"7c00", 846=>x"8500", 847=>x"8000",
---- 848=>x"3000", 849=>x"3300", 850=>x"3e00", 851=>x"4a00", 852=>x"7000", 853=>x"8700", 854=>x"8500",
---- 855=>x"7a00", 856=>x"3000", 857=>x"3400", 858=>x"3e00", 859=>x"5800", 860=>x"7b00", 861=>x"8800",
---- 862=>x"8100", 863=>x"7a00", 864=>x"2e00", 865=>x"3100", 866=>x"b800", 867=>x"6c00", 868=>x"8400",
---- 869=>x"8900", 870=>x"8100", 871=>x"7a00", 872=>x"2e00", 873=>x"3500", 874=>x"5300", 875=>x"7b00",
---- 876=>x"8d00", 877=>x"8800", 878=>x"7e00", 879=>x"7e00", 880=>x"3200", 881=>x"3f00", 882=>x"6300",
---- 883=>x"8400", 884=>x"8e00", 885=>x"8600", 886=>x"7f00", 887=>x"8800", 888=>x"3700", 889=>x"4c00",
---- 890=>x"7700", 891=>x"8b00", 892=>x"8b00", 893=>x"8200", 894=>x"8100", 895=>x"9300", 896=>x"3900",
---- 897=>x"5f00", 898=>x"8400", 899=>x"9200", 900=>x"8900", 901=>x"7e00", 902=>x"8800", 903=>x"9900",
---- 904=>x"3b00", 905=>x"6e00", 906=>x"8c00", 907=>x"8f00", 908=>x"8600", 909=>x"8100", 910=>x"9000",
---- 911=>x"a000", 912=>x"4a00", 913=>x"7900", 914=>x"8e00", 915=>x"8c00", 916=>x"8300", 917=>x"8900",
---- 918=>x"9900", 919=>x"a300", 920=>x"6100", 921=>x"8600", 922=>x"9000", 923=>x"8c00", 924=>x"8200",
---- 925=>x"8e00", 926=>x"9e00", 927=>x"a700", 928=>x"7a00", 929=>x"9100", 930=>x"8f00", 931=>x"8700",
---- 932=>x"8400", 933=>x"6c00", 934=>x"a200", 935=>x"a500", 936=>x"8500", 937=>x"9200", 938=>x"8e00",
---- 939=>x"8400", 940=>x"8900", 941=>x"9a00", 942=>x"a500", 943=>x"a700", 944=>x"8900", 945=>x"9000",
---- 946=>x"8800", 947=>x"8500", 948=>x"8f00", 949=>x"9f00", 950=>x"a600", 951=>x"a300", 952=>x"8b00",
---- 953=>x"8b00", 954=>x"8600", 955=>x"7600", 956=>x"9400", 957=>x"a000", 958=>x"a500", 959=>x"a400",
---- 960=>x"8d00", 961=>x"8700", 962=>x"8000", 963=>x"8a00", 964=>x"9a00", 965=>x"a300", 966=>x"a200",
---- 967=>x"a400", 968=>x"8d00", 969=>x"8500", 970=>x"8100", 971=>x"9000", 972=>x"9d00", 973=>x"a200",
---- 974=>x"a300", 975=>x"a400", 976=>x"8900", 977=>x"8200", 978=>x"8400", 979=>x"9500", 980=>x"a000",
---- 981=>x"a000", 982=>x"a000", 983=>x"a000", 984=>x"8700", 985=>x"8100", 986=>x"8900", 987=>x"9a00",
---- 988=>x"a200", 989=>x"a100", 990=>x"a000", 991=>x"9f00", 992=>x"8500", 993=>x"7e00", 994=>x"9000",
---- 995=>x"9f00", 996=>x"a500", 997=>x"a400", 998=>x"9f00", 999=>x"9f00", 1000=>x"7f00", 1001=>x"8400",
---- 1002=>x"9600", 1003=>x"a200", 1004=>x"a100", 1005=>x"a200", 1006=>x"9f00", 1007=>x"9f00", 1008=>x"8000",
---- 1009=>x"8d00", 1010=>x"9c00", 1011=>x"a100", 1012=>x"a300", 1013=>x"a100", 1014=>x"9f00", 1015=>x"a000",
---- 1016=>x"8000", 1017=>x"8f00", 1018=>x"9e00", 1019=>x"a000", 1020=>x"a100", 1021=>x"9f00", 1022=>x"9e00",
---- 1023=>x"9e00", 1024=>x"8300", 1025=>x"9600", 1026=>x"a000", 1027=>x"a000", 1028=>x"9f00", 1029=>x"9f00",
---- 1030=>x"9e00", 1031=>x"9b00", 1032=>x"8a00", 1033=>x"9900", 1034=>x"a000", 1035=>x"a000", 1036=>x"9f00",
---- 1037=>x"9f00", 1038=>x"9d00", 1039=>x"9c00", 1040=>x"9500", 1041=>x"a100", 1042=>x"a100", 1043=>x"a000",
---- 1044=>x"9d00", 1045=>x"9c00", 1046=>x"9d00", 1047=>x"9a00", 1048=>x"9900", 1049=>x"a300", 1050=>x"9e00",
---- 1051=>x"9e00", 1052=>x"9d00", 1053=>x"9c00", 1054=>x"9b00", 1055=>x"6500", 1056=>x"9d00", 1057=>x"a000",
---- 1058=>x"9f00", 1059=>x"9e00", 1060=>x"9d00", 1061=>x"9c00", 1062=>x"9c00", 1063=>x"6600", 1064=>x"9f00",
---- 1065=>x"9e00", 1066=>x"9f00", 1067=>x"9c00", 1068=>x"9d00", 1069=>x"9e00", 1070=>x"9c00", 1071=>x"9800",
---- 1072=>x"9e00", 1073=>x"9e00", 1074=>x"9f00", 1075=>x"9d00", 1076=>x"9c00", 1077=>x"9f00", 1078=>x"9b00",
---- 1079=>x"9900", 1080=>x"9e00", 1081=>x"9d00", 1082=>x"9c00", 1083=>x"9c00", 1084=>x"9b00", 1085=>x"9c00",
---- 1086=>x"9800", 1087=>x"9900", 1088=>x"9f00", 1089=>x"9d00", 1090=>x"9b00", 1091=>x"9b00", 1092=>x"9b00",
---- 1093=>x"9a00", 1094=>x"9a00", 1095=>x"9900", 1096=>x"9d00", 1097=>x"9a00", 1098=>x"9d00", 1099=>x"9a00",
---- 1100=>x"9800", 1101=>x"9800", 1102=>x"9900", 1103=>x"9800", 1104=>x"9b00", 1105=>x"9b00", 1106=>x"9c00",
---- 1107=>x"9d00", 1108=>x"9800", 1109=>x"9700", 1110=>x"9900", 1111=>x"9400", 1112=>x"9e00", 1113=>x"9b00",
---- 1114=>x"9b00", 1115=>x"9a00", 1116=>x"9900", 1117=>x"9900", 1118=>x"9900", 1119=>x"9800", 1120=>x"9e00",
---- 1121=>x"9900", 1122=>x"9a00", 1123=>x"9900", 1124=>x"9a00", 1125=>x"9700", 1126=>x"9800", 1127=>x"9800",
---- 1128=>x"9b00", 1129=>x"9700", 1130=>x"9a00", 1131=>x"9b00", 1132=>x"9800", 1133=>x"9500", 1134=>x"9600",
---- 1135=>x"9600", 1136=>x"9a00", 1137=>x"9b00", 1138=>x"9800", 1139=>x"9900", 1140=>x"9800", 1141=>x"9700",
---- 1142=>x"9500", 1143=>x"6600", 1144=>x"9d00", 1145=>x"9b00", 1146=>x"9800", 1147=>x"9700", 1148=>x"9800",
---- 1149=>x"9700", 1150=>x"9600", 1151=>x"9600", 1152=>x"6400", 1153=>x"9900", 1154=>x"9a00", 1155=>x"9600",
---- 1156=>x"9500", 1157=>x"9700", 1158=>x"9700", 1159=>x"9700", 1160=>x"9c00", 1161=>x"9800", 1162=>x"9900",
---- 1163=>x"9900", 1164=>x"9900", 1165=>x"9a00", 1166=>x"9800", 1167=>x"9500", 1168=>x"9900", 1169=>x"9800",
---- 1170=>x"9a00", 1171=>x"9700", 1172=>x"9700", 1173=>x"9700", 1174=>x"9600", 1175=>x"9600", 1176=>x"9b00",
---- 1177=>x"9b00", 1178=>x"9b00", 1179=>x"9a00", 1180=>x"9500", 1181=>x"9800", 1182=>x"9900", 1183=>x"9700",
---- 1184=>x"9a00", 1185=>x"9c00", 1186=>x"9a00", 1187=>x"9800", 1188=>x"9600", 1189=>x"9700", 1190=>x"9700",
---- 1191=>x"9600", 1192=>x"9900", 1193=>x"9a00", 1194=>x"9900", 1195=>x"9900", 1196=>x"9800", 1197=>x"6a00",
---- 1198=>x"9300", 1199=>x"9700", 1200=>x"9b00", 1201=>x"9b00", 1202=>x"9a00", 1203=>x"9700", 1204=>x"9700",
---- 1205=>x"9700", 1206=>x"9700", 1207=>x"9400", 1208=>x"9d00", 1209=>x"9900", 1210=>x"9900", 1211=>x"9800",
---- 1212=>x"9800", 1213=>x"9500", 1214=>x"9400", 1215=>x"9500", 1216=>x"9800", 1217=>x"9900", 1218=>x"9900",
---- 1219=>x"9700", 1220=>x"9600", 1221=>x"9500", 1222=>x"9400", 1223=>x"9500", 1224=>x"9b00", 1225=>x"9a00",
---- 1226=>x"9a00", 1227=>x"9800", 1228=>x"9800", 1229=>x"9700", 1230=>x"9500", 1231=>x"9600", 1232=>x"9900",
---- 1233=>x"9a00", 1234=>x"9b00", 1235=>x"9700", 1236=>x"9700", 1237=>x"9900", 1238=>x"9600", 1239=>x"9600",
---- 1240=>x"9b00", 1241=>x"9b00", 1242=>x"9b00", 1243=>x"9900", 1244=>x"9600", 1245=>x"9700", 1246=>x"9800",
---- 1247=>x"9600", 1248=>x"9700", 1249=>x"9900", 1250=>x"9700", 1251=>x"9a00", 1252=>x"9900", 1253=>x"9700",
---- 1254=>x"9700", 1255=>x"9500", 1256=>x"9700", 1257=>x"9700", 1258=>x"9400", 1259=>x"9700", 1260=>x"9800",
---- 1261=>x"9800", 1262=>x"9600", 1263=>x"9400", 1264=>x"9700", 1265=>x"9700", 1266=>x"9600", 1267=>x"9300",
---- 1268=>x"9600", 1269=>x"9500", 1270=>x"9600", 1271=>x"9900", 1272=>x"9600", 1273=>x"9500", 1274=>x"9700",
---- 1275=>x"6a00", 1276=>x"9700", 1277=>x"9600", 1278=>x"9300", 1279=>x"9400", 1280=>x"9600", 1281=>x"9700",
---- 1282=>x"9700", 1283=>x"6900", 1284=>x"9700", 1285=>x"9500", 1286=>x"9500", 1287=>x"9500", 1288=>x"9700",
---- 1289=>x"9700", 1290=>x"9600", 1291=>x"9600", 1292=>x"9700", 1293=>x"9600", 1294=>x"9400", 1295=>x"9000",
---- 1296=>x"9500", 1297=>x"9400", 1298=>x"9400", 1299=>x"9600", 1300=>x"9500", 1301=>x"9500", 1302=>x"9300",
---- 1303=>x"9400", 1304=>x"9600", 1305=>x"9500", 1306=>x"9700", 1307=>x"9800", 1308=>x"9600", 1309=>x"9400",
---- 1310=>x"9400", 1311=>x"9500", 1312=>x"9500", 1313=>x"9500", 1314=>x"9800", 1315=>x"9500", 1316=>x"9500",
---- 1317=>x"9700", 1318=>x"9500", 1319=>x"9400", 1320=>x"9400", 1321=>x"9600", 1322=>x"6b00", 1323=>x"9400",
---- 1324=>x"9300", 1325=>x"9400", 1326=>x"9600", 1327=>x"9300", 1328=>x"9400", 1329=>x"9500", 1330=>x"9500",
---- 1331=>x"9200", 1332=>x"9500", 1333=>x"9600", 1334=>x"9300", 1335=>x"9200", 1336=>x"9200", 1337=>x"9400",
---- 1338=>x"9600", 1339=>x"9600", 1340=>x"9500", 1341=>x"9300", 1342=>x"9000", 1343=>x"9400", 1344=>x"9400",
---- 1345=>x"9500", 1346=>x"9400", 1347=>x"9300", 1348=>x"9200", 1349=>x"9100", 1350=>x"9100", 1351=>x"9100",
---- 1352=>x"9300", 1353=>x"9500", 1354=>x"9400", 1355=>x"9500", 1356=>x"9300", 1357=>x"8e00", 1358=>x"9000",
---- 1359=>x"9200", 1360=>x"9300", 1361=>x"9400", 1362=>x"9600", 1363=>x"9400", 1364=>x"9100", 1365=>x"9100",
---- 1366=>x"9000", 1367=>x"9200", 1368=>x"9200", 1369=>x"9300", 1370=>x"9500", 1371=>x"9400", 1372=>x"9000",
---- 1373=>x"9300", 1374=>x"9400", 1375=>x"9000", 1376=>x"9400", 1377=>x"9600", 1378=>x"9500", 1379=>x"9300",
---- 1380=>x"9300", 1381=>x"9400", 1382=>x"9000", 1383=>x"9200", 1384=>x"9300", 1385=>x"9800", 1386=>x"9300",
---- 1387=>x"9200", 1388=>x"9500", 1389=>x"9400", 1390=>x"9000", 1391=>x"9100", 1392=>x"9300", 1393=>x"9400",
---- 1394=>x"9400", 1395=>x"9400", 1396=>x"9400", 1397=>x"9300", 1398=>x"9300", 1399=>x"9100", 1400=>x"9400",
---- 1401=>x"9500", 1402=>x"9400", 1403=>x"9100", 1404=>x"9200", 1405=>x"9400", 1406=>x"9500", 1407=>x"6e00",
---- 1408=>x"9200", 1409=>x"9500", 1410=>x"9300", 1411=>x"9200", 1412=>x"9400", 1413=>x"9500", 1414=>x"9200",
---- 1415=>x"9100", 1416=>x"9100", 1417=>x"9300", 1418=>x"9200", 1419=>x"9000", 1420=>x"9400", 1421=>x"9300",
---- 1422=>x"9200", 1423=>x"9200", 1424=>x"9500", 1425=>x"9700", 1426=>x"6b00", 1427=>x"9300", 1428=>x"9400",
---- 1429=>x"9300", 1430=>x"9100", 1431=>x"9000", 1432=>x"9800", 1433=>x"9600", 1434=>x"9500", 1435=>x"9700",
---- 1436=>x"9300", 1437=>x"9200", 1438=>x"9100", 1439=>x"9000", 1440=>x"9700", 1441=>x"9500", 1442=>x"9500",
---- 1443=>x"9800", 1444=>x"9500", 1445=>x"9300", 1446=>x"9100", 1447=>x"9200", 1448=>x"9500", 1449=>x"9500",
---- 1450=>x"9500", 1451=>x"9400", 1452=>x"9600", 1453=>x"9200", 1454=>x"9100", 1455=>x"9100", 1456=>x"9900",
---- 1457=>x"9700", 1458=>x"9500", 1459=>x"9500", 1460=>x"9500", 1461=>x"9500", 1462=>x"9200", 1463=>x"9200",
---- 1464=>x"9d00", 1465=>x"9a00", 1466=>x"9800", 1467=>x"9700", 1468=>x"9500", 1469=>x"9400", 1470=>x"9200",
---- 1471=>x"9100", 1472=>x"9a00", 1473=>x"9600", 1474=>x"9700", 1475=>x"9600", 1476=>x"9500", 1477=>x"9400",
---- 1478=>x"9200", 1479=>x"9200", 1480=>x"9700", 1481=>x"9900", 1482=>x"9500", 1483=>x"9500", 1484=>x"9400",
---- 1485=>x"9400", 1486=>x"9400", 1487=>x"9100", 1488=>x"9900", 1489=>x"9b00", 1490=>x"9600", 1491=>x"9400",
---- 1492=>x"9600", 1493=>x"9500", 1494=>x"9000", 1495=>x"9000", 1496=>x"9900", 1497=>x"9700", 1498=>x"9600",
---- 1499=>x"9800", 1500=>x"9600", 1501=>x"9500", 1502=>x"6e00", 1503=>x"8f00", 1504=>x"9800", 1505=>x"9800",
---- 1506=>x"9800", 1507=>x"9700", 1508=>x"9400", 1509=>x"9300", 1510=>x"9000", 1511=>x"8e00", 1512=>x"9500",
---- 1513=>x"9700", 1514=>x"9500", 1515=>x"9400", 1516=>x"9500", 1517=>x"9300", 1518=>x"9000", 1519=>x"8e00",
---- 1520=>x"9700", 1521=>x"9500", 1522=>x"9500", 1523=>x"9400", 1524=>x"9100", 1525=>x"8f00", 1526=>x"8e00",
---- 1527=>x"8d00", 1528=>x"9400", 1529=>x"9600", 1530=>x"9500", 1531=>x"9200", 1532=>x"9100", 1533=>x"8f00",
---- 1534=>x"8f00", 1535=>x"8c00", 1536=>x"9700", 1537=>x"9300", 1538=>x"9400", 1539=>x"9300", 1540=>x"9200",
---- 1541=>x"9000", 1542=>x"8f00", 1543=>x"8d00", 1544=>x"9400", 1545=>x"9500", 1546=>x"9200", 1547=>x"9100",
---- 1548=>x"9000", 1549=>x"9100", 1550=>x"8d00", 1551=>x"7300", 1552=>x"8f00", 1553=>x"9600", 1554=>x"9500",
---- 1555=>x"9300", 1556=>x"6f00", 1557=>x"8f00", 1558=>x"8f00", 1559=>x"8c00", 1560=>x"8700", 1561=>x"8b00",
---- 1562=>x"7200", 1563=>x"8f00", 1564=>x"8e00", 1565=>x"8c00", 1566=>x"8c00", 1567=>x"8c00", 1568=>x"7c00",
---- 1569=>x"8000", 1570=>x"8100", 1571=>x"8400", 1572=>x"8500", 1573=>x"8600", 1574=>x"8800", 1575=>x"8900",
---- 1576=>x"6f00", 1577=>x"7200", 1578=>x"7500", 1579=>x"7900", 1580=>x"7800", 1581=>x"7a00", 1582=>x"7b00",
---- 1583=>x"7d00", 1584=>x"6600", 1585=>x"6600", 1586=>x"6900", 1587=>x"7000", 1588=>x"7000", 1589=>x"7300",
---- 1590=>x"7000", 1591=>x"7000", 1592=>x"6500", 1593=>x"6400", 1594=>x"6400", 1595=>x"6200", 1596=>x"6400",
---- 1597=>x"6900", 1598=>x"6600", 1599=>x"9b00", 1600=>x"6a00", 1601=>x"6400", 1602=>x"6400", 1603=>x"6100",
---- 1604=>x"5f00", 1605=>x"6100", 1606=>x"6000", 1607=>x"5c00", 1608=>x"7100", 1609=>x"6e00", 1610=>x"6900",
---- 1611=>x"6500", 1612=>x"6100", 1613=>x"5f00", 1614=>x"5e00", 1615=>x"5700", 1616=>x"7a00", 1617=>x"7600",
---- 1618=>x"7200", 1619=>x"6b00", 1620=>x"6800", 1621=>x"6b00", 1622=>x"5f00", 1623=>x"5800", 1624=>x"7e00",
---- 1625=>x"7a00", 1626=>x"7500", 1627=>x"7500", 1628=>x"7200", 1629=>x"6d00", 1630=>x"6800", 1631=>x"6100",
---- 1632=>x"8100", 1633=>x"7d00", 1634=>x"7b00", 1635=>x"7900", 1636=>x"7600", 1637=>x"7500", 1638=>x"7400",
---- 1639=>x"9600", 1640=>x"8200", 1641=>x"7f00", 1642=>x"8300", 1643=>x"8100", 1644=>x"7b00", 1645=>x"7c00",
---- 1646=>x"7700", 1647=>x"7100", 1648=>x"8700", 1649=>x"8200", 1650=>x"8200", 1651=>x"8000", 1652=>x"7f00",
---- 1653=>x"7f00", 1654=>x"7800", 1655=>x"7700", 1656=>x"8600", 1657=>x"8600", 1658=>x"8200", 1659=>x"8400",
---- 1660=>x"7f00", 1661=>x"7e00", 1662=>x"7a00", 1663=>x"7b00", 1664=>x"8500", 1665=>x"8600", 1666=>x"8500",
---- 1667=>x"8400", 1668=>x"7f00", 1669=>x"8000", 1670=>x"7c00", 1671=>x"7e00", 1672=>x"8600", 1673=>x"8700",
---- 1674=>x"8600", 1675=>x"8200", 1676=>x"8100", 1677=>x"7e00", 1678=>x"8100", 1679=>x"7f00", 1680=>x"8700",
---- 1681=>x"8a00", 1682=>x"8400", 1683=>x"8500", 1684=>x"8100", 1685=>x"7e00", 1686=>x"8200", 1687=>x"7f00",
---- 1688=>x"8900", 1689=>x"8900", 1690=>x"8600", 1691=>x"8300", 1692=>x"8200", 1693=>x"8200", 1694=>x"7e00",
---- 1695=>x"7b00", 1696=>x"8900", 1697=>x"8300", 1698=>x"8700", 1699=>x"8300", 1700=>x"7f00", 1701=>x"7e00",
---- 1702=>x"7d00", 1703=>x"7a00", 1704=>x"8600", 1705=>x"8500", 1706=>x"8500", 1707=>x"8100", 1708=>x"7d00",
---- 1709=>x"7b00", 1710=>x"7b00", 1711=>x"7900", 1712=>x"8700", 1713=>x"8400", 1714=>x"8200", 1715=>x"8000",
---- 1716=>x"7c00", 1717=>x"7e00", 1718=>x"7a00", 1719=>x"7f00", 1720=>x"8600", 1721=>x"8200", 1722=>x"8000",
---- 1723=>x"7d00", 1724=>x"7a00", 1725=>x"7b00", 1726=>x"7900", 1727=>x"8b00", 1728=>x"8100", 1729=>x"8100",
---- 1730=>x"8200", 1731=>x"7e00", 1732=>x"8000", 1733=>x"7800", 1734=>x"7b00", 1735=>x"9d00", 1736=>x"7f00",
---- 1737=>x"7f00", 1738=>x"8000", 1739=>x"7e00", 1740=>x"7f00", 1741=>x"7700", 1742=>x"8000", 1743=>x"ae00",
---- 1744=>x"8200", 1745=>x"7f00", 1746=>x"8200", 1747=>x"7c00", 1748=>x"7900", 1749=>x"7700", 1750=>x"8500",
---- 1751=>x"ba00", 1752=>x"8200", 1753=>x"7e00", 1754=>x"7c00", 1755=>x"7900", 1756=>x"7800", 1757=>x"7800",
---- 1758=>x"6f00", 1759=>x"c100", 1760=>x"8300", 1761=>x"7d00", 1762=>x"7f00", 1763=>x"7d00", 1764=>x"7a00",
---- 1765=>x"7c00", 1766=>x"9600", 1767=>x"c400", 1768=>x"8000", 1769=>x"8100", 1770=>x"7b00", 1771=>x"7a00",
---- 1772=>x"7b00", 1773=>x"8200", 1774=>x"9c00", 1775=>x"c700", 1776=>x"7e00", 1777=>x"7c00", 1778=>x"7b00",
---- 1779=>x"7d00", 1780=>x"7f00", 1781=>x"8300", 1782=>x"a300", 1783=>x"ca00", 1784=>x"7f00", 1785=>x"7f00",
---- 1786=>x"7f00", 1787=>x"7f00", 1788=>x"7f00", 1789=>x"8200", 1790=>x"a800", 1791=>x"cb00", 1792=>x"8200",
---- 1793=>x"7e00", 1794=>x"8000", 1795=>x"8200", 1796=>x"7e00", 1797=>x"8400", 1798=>x"a200", 1799=>x"c200",
---- 1800=>x"7e00", 1801=>x"8200", 1802=>x"8500", 1803=>x"8400", 1804=>x"8100", 1805=>x"8400", 1806=>x"9600",
---- 1807=>x"b800", 1808=>x"8000", 1809=>x"8300", 1810=>x"8400", 1811=>x"8500", 1812=>x"8800", 1813=>x"8600",
---- 1814=>x"8a00", 1815=>x"9d00", 1816=>x"8300", 1817=>x"8600", 1818=>x"8800", 1819=>x"8700", 1820=>x"8c00",
---- 1821=>x"8a00", 1822=>x"8a00", 1823=>x"8b00", 1824=>x"8800", 1825=>x"8800", 1826=>x"8d00", 1827=>x"8d00",
---- 1828=>x"8e00", 1829=>x"8d00", 1830=>x"8c00", 1831=>x"8a00", 1832=>x"8800", 1833=>x"6f00", 1834=>x"9100",
---- 1835=>x"9300", 1836=>x"9400", 1837=>x"9200", 1838=>x"8f00", 1839=>x"8c00", 1840=>x"8a00", 1841=>x"8d00",
---- 1842=>x"9600", 1843=>x"9800", 1844=>x"9600", 1845=>x"9100", 1846=>x"9000", 1847=>x"8c00", 1848=>x"9200",
---- 1849=>x"9500", 1850=>x"9900", 1851=>x"9b00", 1852=>x"9400", 1853=>x"8d00", 1854=>x"8700", 1855=>x"8300",
---- 1856=>x"9000", 1857=>x"9900", 1858=>x"a000", 1859=>x"9e00", 1860=>x"9700", 1861=>x"8e00", 1862=>x"7c00",
---- 1863=>x"7d00", 1864=>x"8900", 1865=>x"9100", 1866=>x"9d00", 1867=>x"a100", 1868=>x"9600", 1869=>x"8f00",
---- 1870=>x"9100", 1871=>x"9200", 1872=>x"7700", 1873=>x"8600", 1874=>x"8e00", 1875=>x"9200", 1876=>x"9400",
---- 1877=>x"a200", 1878=>x"a700", 1879=>x"9b00", 1880=>x"5b00", 1881=>x"6c00", 1882=>x"7100", 1883=>x"8900",
---- 1884=>x"ad00", 1885=>x"bc00", 1886=>x"b400", 1887=>x"a000", 1888=>x"3c00", 1889=>x"5000", 1890=>x"6d00",
---- 1891=>x"a200", 1892=>x"c300", 1893=>x"c300", 1894=>x"bd00", 1895=>x"a800", 1896=>x"2b00", 1897=>x"4300",
---- 1898=>x"8a00", 1899=>x"bd00", 1900=>x"ca00", 1901=>x"ca00", 1902=>x"bb00", 1903=>x"9f00", 1904=>x"2000",
---- 1905=>x"4500", 1906=>x"9b00", 1907=>x"c800", 1908=>x"ce00", 1909=>x"d000", 1910=>x"b100", 1911=>x"9400",
---- 1912=>x"2700", 1913=>x"4500", 1914=>x"9800", 1915=>x"c400", 1916=>x"cc00", 1917=>x"cb00", 1918=>x"ae00",
---- 1919=>x"9f00", 1920=>x"3100", 1921=>x"4a00", 1922=>x"8d00", 1923=>x"b900", 1924=>x"ca00", 1925=>x"c900",
---- 1926=>x"bd00", 1927=>x"b800", 1928=>x"3d00", 1929=>x"4800", 1930=>x"7e00", 1931=>x"b500", 1932=>x"c900",
---- 1933=>x"ca00", 1934=>x"ca00", 1935=>x"c500", 1936=>x"4d00", 1937=>x"5700", 1938=>x"8300", 1939=>x"b700",
---- 1940=>x"cd00", 1941=>x"d200", 1942=>x"d100", 1943=>x"c800", 1944=>x"5200", 1945=>x"5f00", 1946=>x"8c00",
---- 1947=>x"b500", 1948=>x"cd00", 1949=>x"d500", 1950=>x"d000", 1951=>x"bf00", 1952=>x"5900", 1953=>x"5e00",
---- 1954=>x"8800", 1955=>x"b200", 1956=>x"ca00", 1957=>x"ce00", 1958=>x"c300", 1959=>x"ab00", 1960=>x"6100",
---- 1961=>x"6100", 1962=>x"7b00", 1963=>x"a200", 1964=>x"b700", 1965=>x"b600", 1966=>x"a700", 1967=>x"7b00",
---- 1968=>x"6900", 1969=>x"6800", 1970=>x"7000", 1971=>x"8900", 1972=>x"9400", 1973=>x"8c00", 1974=>x"7300",
---- 1975=>x"5800", 1976=>x"7000", 1977=>x"7000", 1978=>x"6d00", 1979=>x"7100", 1980=>x"7500", 1981=>x"6e00",
---- 1982=>x"6000", 1983=>x"5700", 1984=>x"7300", 1985=>x"7200", 1986=>x"6e00", 1987=>x"6b00", 1988=>x"6900",
---- 1989=>x"6500", 1990=>x"5f00", 1991=>x"5b00", 1992=>x"7200", 1993=>x"7100", 1994=>x"8f00", 1995=>x"6800",
---- 1996=>x"6700", 1997=>x"6600", 1998=>x"6200", 1999=>x"6000", 2000=>x"7400", 2001=>x"7200", 2002=>x"7000",
---- 2003=>x"6d00", 2004=>x"6a00", 2005=>x"6800", 2006=>x"6500", 2007=>x"6200", 2008=>x"7200", 2009=>x"7400",
---- 2010=>x"7100", 2011=>x"7000", 2012=>x"6b00", 2013=>x"6b00", 2014=>x"6a00", 2015=>x"6e00", 2016=>x"7300",
---- 2017=>x"7400", 2018=>x"7100", 2019=>x"6e00", 2020=>x"6e00", 2021=>x"7100", 2022=>x"7300", 2023=>x"7800",
---- 2024=>x"7500", 2025=>x"7500", 2026=>x"7100", 2027=>x"7500", 2028=>x"7600", 2029=>x"7500", 2030=>x"7b00",
---- 2031=>x"7f00", 2032=>x"7a00", 2033=>x"7700", 2034=>x"7600", 2035=>x"7900", 2036=>x"7d00", 2037=>x"8200",
---- 2038=>x"8700", 2039=>x"8500", 2040=>x"7b00", 2041=>x"7d00", 2042=>x"7d00", 2043=>x"8400", 2044=>x"8400",
---- 2045=>x"8a00", 2046=>x"8b00", 2047=>x"8600"),
---- 27 => (0=>x"7300", 1=>x"7600", 2=>x"7600", 3=>x"7900", 4=>x"8100", 5=>x"7600", 6=>x"7900", 7=>x"7900",
---- 8=>x"7300", 9=>x"7600", 10=>x"7600", 11=>x"7900", 12=>x"7d00", 13=>x"7600", 14=>x"7900",
---- 15=>x"7900", 16=>x"7300", 17=>x"7600", 18=>x"7600", 19=>x"7800", 20=>x"7d00", 21=>x"7600",
---- 22=>x"7800", 23=>x"7b00", 24=>x"7100", 25=>x"7400", 26=>x"7700", 27=>x"7600", 28=>x"7700",
---- 29=>x"7900", 30=>x"8800", 31=>x"7b00", 32=>x"6f00", 33=>x"8f00", 34=>x"7500", 35=>x"7700",
---- 36=>x"7700", 37=>x"7800", 38=>x"7700", 39=>x"7a00", 40=>x"6a00", 41=>x"6e00", 42=>x"7100",
---- 43=>x"7300", 44=>x"7a00", 45=>x"8800", 46=>x"7700", 47=>x"7900", 48=>x"6800", 49=>x"6e00",
---- 50=>x"7000", 51=>x"7300", 52=>x"7500", 53=>x"7a00", 54=>x"7700", 55=>x"7800", 56=>x"6a00",
---- 57=>x"6d00", 58=>x"6e00", 59=>x"7000", 60=>x"7500", 61=>x"7500", 62=>x"7400", 63=>x"7600",
---- 64=>x"6800", 65=>x"6800", 66=>x"6c00", 67=>x"6e00", 68=>x"7600", 69=>x"7400", 70=>x"7400",
---- 71=>x"7800", 72=>x"6d00", 73=>x"6700", 74=>x"6900", 75=>x"9300", 76=>x"7100", 77=>x"7400",
---- 78=>x"7500", 79=>x"7700", 80=>x"8600", 81=>x"6600", 82=>x"6d00", 83=>x"6a00", 84=>x"7000",
---- 85=>x"7000", 86=>x"7200", 87=>x"7600", 88=>x"a300", 89=>x"7100", 90=>x"6900", 91=>x"6a00",
---- 92=>x"6f00", 93=>x"7100", 94=>x"7300", 95=>x"7500", 96=>x"c000", 97=>x"9100", 98=>x"6700",
---- 99=>x"6900", 100=>x"6d00", 101=>x"6f00", 102=>x"7400", 103=>x"7800", 104=>x"ce00", 105=>x"b100",
---- 106=>x"7800", 107=>x"6400", 108=>x"6b00", 109=>x"6f00", 110=>x"7300", 111=>x"7200", 112=>x"d500",
---- 113=>x"c700", 114=>x"9a00", 115=>x"6900", 116=>x"6900", 117=>x"6d00", 118=>x"7200", 119=>x"7200",
---- 120=>x"dc00", 121=>x"d500", 122=>x"ba00", 123=>x"7f00", 124=>x"6500", 125=>x"6d00", 126=>x"6f00",
---- 127=>x"7400", 128=>x"de00", 129=>x"dc00", 130=>x"d100", 131=>x"b100", 132=>x"7c00", 133=>x"6d00",
---- 134=>x"6e00", 135=>x"7000", 136=>x"df00", 137=>x"de00", 138=>x"d800", 139=>x"c300", 140=>x"9000",
---- 141=>x"6800", 142=>x"6900", 143=>x"6b00", 144=>x"de00", 145=>x"e100", 146=>x"db00", 147=>x"cf00",
---- 148=>x"b300", 149=>x"7a00", 150=>x"6400", 151=>x"6800", 152=>x"de00", 153=>x"df00", 154=>x"e100",
---- 155=>x"d900", 156=>x"ca00", 157=>x"9c00", 158=>x"6700", 159=>x"6000", 160=>x"df00", 161=>x"de00",
---- 162=>x"e100", 163=>x"de00", 164=>x"d400", 165=>x"bc00", 166=>x"8400", 167=>x"6200", 168=>x"dc00",
---- 169=>x"de00", 170=>x"2000", 171=>x"df00", 172=>x"db00", 173=>x"ca00", 174=>x"a300", 175=>x"6c00",
---- 176=>x"da00", 177=>x"dd00", 178=>x"df00", 179=>x"e100", 180=>x"df00", 181=>x"d400", 182=>x"bf00",
---- 183=>x"8600", 184=>x"d900", 185=>x"dc00", 186=>x"e000", 187=>x"e000", 188=>x"e000", 189=>x"db00",
---- 190=>x"cf00", 191=>x"ab00", 192=>x"d300", 193=>x"da00", 194=>x"dc00", 195=>x"dc00", 196=>x"df00",
---- 197=>x"2000", 198=>x"d800", 199=>x"c600", 200=>x"d000", 201=>x"d700", 202=>x"d900", 203=>x"de00",
---- 204=>x"e000", 205=>x"e200", 206=>x"df00", 207=>x"d300", 208=>x"c500", 209=>x"d300", 210=>x"2700",
---- 211=>x"db00", 212=>x"df00", 213=>x"e200", 214=>x"e300", 215=>x"dd00", 216=>x"b400", 217=>x"cd00",
---- 218=>x"d600", 219=>x"dc00", 220=>x"df00", 221=>x"e000", 222=>x"1c00", 223=>x"e200", 224=>x"9b00",
---- 225=>x"c200", 226=>x"d200", 227=>x"db00", 228=>x"df00", 229=>x"e000", 230=>x"e200", 231=>x"e400",
---- 232=>x"8a00", 233=>x"ac00", 234=>x"cd00", 235=>x"d700", 236=>x"dd00", 237=>x"df00", 238=>x"e200",
---- 239=>x"e300", 240=>x"7700", 241=>x"9300", 242=>x"bd00", 243=>x"d000", 244=>x"d900", 245=>x"dd00",
---- 246=>x"e200", 247=>x"e400", 248=>x"8c00", 249=>x"8b00", 250=>x"a500", 251=>x"c600", 252=>x"d500",
---- 253=>x"dc00", 254=>x"e100", 255=>x"e500", 256=>x"8d00", 257=>x"8c00", 258=>x"9200", 259=>x"b300",
---- 260=>x"d300", 261=>x"dc00", 262=>x"e400", 263=>x"e600", 264=>x"8f00", 265=>x"8f00", 266=>x"8e00",
---- 267=>x"9900", 268=>x"c500", 269=>x"da00", 270=>x"e100", 271=>x"e000", 272=>x"9100", 273=>x"9300",
---- 274=>x"9300", 275=>x"9100", 276=>x"ae00", 277=>x"d200", 278=>x"db00", 279=>x"d100", 280=>x"9200",
---- 281=>x"9400", 282=>x"9800", 283=>x"9600", 284=>x"a300", 285=>x"c900", 286=>x"c400", 287=>x"8500",
---- 288=>x"9400", 289=>x"6b00", 290=>x"9900", 291=>x"9a00", 292=>x"a000", 293=>x"a300", 294=>x"7500",
---- 295=>x"3600", 296=>x"9600", 297=>x"9600", 298=>x"9900", 299=>x"9e00", 300=>x"9900", 301=>x"6f00",
---- 302=>x"3900", 303=>x"2d00", 304=>x"9600", 305=>x"9900", 306=>x"9c00", 307=>x"9d00", 308=>x"8300",
---- 309=>x"4700", 310=>x"2900", 311=>x"2d00", 312=>x"9900", 313=>x"9b00", 314=>x"9e00", 315=>x"8b00",
---- 316=>x"5800", 317=>x"3200", 318=>x"2a00", 319=>x"2b00", 320=>x"9a00", 321=>x"9d00", 322=>x"9100",
---- 323=>x"6700", 324=>x"3000", 325=>x"2e00", 326=>x"2c00", 327=>x"2e00", 328=>x"9d00", 329=>x"9800",
---- 330=>x"7500", 331=>x"3d00", 332=>x"2900", 333=>x"2c00", 334=>x"2800", 335=>x"2b00", 336=>x"9b00",
---- 337=>x"8400", 338=>x"4e00", 339=>x"2c00", 340=>x"2b00", 341=>x"2600", 342=>x"2500", 343=>x"2a00",
---- 344=>x"9200", 345=>x"5d00", 346=>x"2d00", 347=>x"2500", 348=>x"2700", 349=>x"2900", 350=>x"2800",
---- 351=>x"d600", 352=>x"7100", 353=>x"3700", 354=>x"2800", 355=>x"2700", 356=>x"2b00", 357=>x"2a00",
---- 358=>x"2b00", 359=>x"2d00", 360=>x"4500", 361=>x"2900", 362=>x"3c00", 363=>x"4100", 364=>x"3700",
---- 365=>x"2c00", 366=>x"2a00", 367=>x"3300", 368=>x"2e00", 369=>x"2e00", 370=>x"3500", 371=>x"3500",
---- 372=>x"2f00", 373=>x"d200", 374=>x"2c00", 375=>x"3300", 376=>x"2700", 377=>x"2600", 378=>x"2900",
---- 379=>x"2b00", 380=>x"2a00", 381=>x"2f00", 382=>x"3200", 383=>x"3600", 384=>x"2700", 385=>x"2400",
---- 386=>x"2c00", 387=>x"2b00", 388=>x"3000", 389=>x"3400", 390=>x"3900", 391=>x"3800", 392=>x"2700",
---- 393=>x"2700", 394=>x"2800", 395=>x"2e00", 396=>x"3200", 397=>x"3b00", 398=>x"3a00", 399=>x"3800",
---- 400=>x"2600", 401=>x"2800", 402=>x"2b00", 403=>x"2d00", 404=>x"3500", 405=>x"3600", 406=>x"3900",
---- 407=>x"3a00", 408=>x"2900", 409=>x"2900", 410=>x"2f00", 411=>x"2f00", 412=>x"3600", 413=>x"3a00",
---- 414=>x"3500", 415=>x"3400", 416=>x"2d00", 417=>x"2f00", 418=>x"3000", 419=>x"3200", 420=>x"3600",
---- 421=>x"3700", 422=>x"3300", 423=>x"3300", 424=>x"2c00", 425=>x"2e00", 426=>x"3300", 427=>x"3700",
---- 428=>x"3600", 429=>x"3500", 430=>x"3b00", 431=>x"3500", 432=>x"ce00", 433=>x"2f00", 434=>x"3500",
---- 435=>x"3400", 436=>x"3400", 437=>x"3700", 438=>x"3700", 439=>x"3300", 440=>x"3300", 441=>x"3500",
---- 442=>x"3c00", 443=>x"3600", 444=>x"2e00", 445=>x"3600", 446=>x"3600", 447=>x"3600", 448=>x"3400",
---- 449=>x"3500", 450=>x"3900", 451=>x"3600", 452=>x"3200", 453=>x"3700", 454=>x"3a00", 455=>x"3b00",
---- 456=>x"3a00", 457=>x"3500", 458=>x"3500", 459=>x"3400", 460=>x"3400", 461=>x"3800", 462=>x"3f00",
---- 463=>x"c700", 464=>x"3a00", 465=>x"3900", 466=>x"3400", 467=>x"c500", 468=>x"3900", 469=>x"3200",
---- 470=>x"3200", 471=>x"3300", 472=>x"3700", 473=>x"3400", 474=>x"3200", 475=>x"3b00", 476=>x"3e00",
---- 477=>x"3600", 478=>x"3400", 479=>x"3200", 480=>x"3800", 481=>x"3600", 482=>x"3700", 483=>x"3600",
---- 484=>x"3300", 485=>x"3100", 486=>x"2e00", 487=>x"3000", 488=>x"3600", 489=>x"3800", 490=>x"3a00",
---- 491=>x"3100", 492=>x"3300", 493=>x"2f00", 494=>x"3000", 495=>x"3600", 496=>x"3500", 497=>x"3500",
---- 498=>x"3500", 499=>x"3300", 500=>x"3200", 501=>x"3100", 502=>x"3200", 503=>x"3100", 504=>x"3400",
---- 505=>x"3400", 506=>x"3800", 507=>x"3100", 508=>x"2c00", 509=>x"3000", 510=>x"3100", 511=>x"2e00",
---- 512=>x"3400", 513=>x"3100", 514=>x"2f00", 515=>x"2b00", 516=>x"2c00", 517=>x"3200", 518=>x"2f00",
---- 519=>x"2c00", 520=>x"3a00", 521=>x"2f00", 522=>x"2f00", 523=>x"2d00", 524=>x"2b00", 525=>x"2d00",
---- 526=>x"2c00", 527=>x"2e00", 528=>x"3a00", 529=>x"2f00", 530=>x"3200", 531=>x"3000", 532=>x"2f00",
---- 533=>x"2f00", 534=>x"2b00", 535=>x"2e00", 536=>x"3900", 537=>x"3700", 538=>x"3900", 539=>x"3200",
---- 540=>x"2f00", 541=>x"2f00", 542=>x"3100", 543=>x"3500", 544=>x"3300", 545=>x"3400", 546=>x"3500",
---- 547=>x"3000", 548=>x"2b00", 549=>x"2b00", 550=>x"2b00", 551=>x"3300", 552=>x"3200", 553=>x"3200",
---- 554=>x"3500", 555=>x"3000", 556=>x"2c00", 557=>x"2e00", 558=>x"2900", 559=>x"3000", 560=>x"3300",
---- 561=>x"3200", 562=>x"2e00", 563=>x"2f00", 564=>x"2900", 565=>x"2a00", 566=>x"2c00", 567=>x"3200",
---- 568=>x"3400", 569=>x"3100", 570=>x"2e00", 571=>x"2800", 572=>x"2900", 573=>x"3100", 574=>x"3100",
---- 575=>x"3400", 576=>x"3800", 577=>x"3100", 578=>x"2f00", 579=>x"2c00", 580=>x"2e00", 581=>x"3200",
---- 582=>x"2f00", 583=>x"3200", 584=>x"3800", 585=>x"3200", 586=>x"2e00", 587=>x"2800", 588=>x"2e00",
---- 589=>x"3100", 590=>x"2e00", 591=>x"3400", 592=>x"2f00", 593=>x"2d00", 594=>x"2b00", 595=>x"2d00",
---- 596=>x"2e00", 597=>x"3500", 598=>x"3700", 599=>x"3600", 600=>x"3300", 601=>x"2e00", 602=>x"2a00",
---- 603=>x"3000", 604=>x"2d00", 605=>x"3700", 606=>x"3900", 607=>x"3100", 608=>x"3f00", 609=>x"2d00",
---- 610=>x"2e00", 611=>x"2f00", 612=>x"3300", 613=>x"3800", 614=>x"3900", 615=>x"2d00", 616=>x"3200",
---- 617=>x"2d00", 618=>x"2e00", 619=>x"3000", 620=>x"3100", 621=>x"3100", 622=>x"3500", 623=>x"3100",
---- 624=>x"2d00", 625=>x"2a00", 626=>x"d100", 627=>x"d000", 628=>x"2a00", 629=>x"2d00", 630=>x"3900",
---- 631=>x"4300", 632=>x"2c00", 633=>x"2b00", 634=>x"3200", 635=>x"2f00", 636=>x"2c00", 637=>x"3200",
---- 638=>x"4400", 639=>x"5100", 640=>x"2d00", 641=>x"3200", 642=>x"3300", 643=>x"2d00", 644=>x"2f00",
---- 645=>x"3900", 646=>x"4700", 647=>x"5b00", 648=>x"3100", 649=>x"3500", 650=>x"3200", 651=>x"2e00",
---- 652=>x"3100", 653=>x"4200", 654=>x"4b00", 655=>x"6a00", 656=>x"3000", 657=>x"3500", 658=>x"2f00",
---- 659=>x"2e00", 660=>x"3800", 661=>x"4400", 662=>x"5b00", 663=>x"7f00", 664=>x"3400", 665=>x"3600",
---- 666=>x"3000", 667=>x"3400", 668=>x"4000", 669=>x"4700", 670=>x"6c00", 671=>x"9000", 672=>x"3a00",
---- 673=>x"3500", 674=>x"3200", 675=>x"3300", 676=>x"3d00", 677=>x"5800", 678=>x"8100", 679=>x"9800",
---- 680=>x"3a00", 681=>x"3400", 682=>x"3500", 683=>x"3800", 684=>x"4200", 685=>x"6b00", 686=>x"9000",
---- 687=>x"9b00", 688=>x"3200", 689=>x"3500", 690=>x"3800", 691=>x"3b00", 692=>x"5600", 693=>x"7f00",
---- 694=>x"9800", 695=>x"9a00", 696=>x"3400", 697=>x"3200", 698=>x"3600", 699=>x"4100", 700=>x"6900",
---- 701=>x"8d00", 702=>x"9700", 703=>x"9800", 704=>x"3500", 705=>x"3000", 706=>x"3900", 707=>x"5600",
---- 708=>x"7c00", 709=>x"9600", 710=>x"9700", 711=>x"9300", 712=>x"2d00", 713=>x"2e00", 714=>x"4300",
---- 715=>x"6b00", 716=>x"8e00", 717=>x"9900", 718=>x"9600", 719=>x"9100", 720=>x"2900", 721=>x"2c00",
---- 722=>x"5100", 723=>x"8000", 724=>x"9500", 725=>x"9500", 726=>x"9100", 727=>x"8e00", 728=>x"2900",
---- 729=>x"3400", 730=>x"6200", 731=>x"8c00", 732=>x"9500", 733=>x"9300", 734=>x"8f00", 735=>x"8f00",
---- 736=>x"2500", 737=>x"4400", 738=>x"7900", 739=>x"6b00", 740=>x"6800", 741=>x"9100", 742=>x"9000",
---- 743=>x"9300", 744=>x"3200", 745=>x"5d00", 746=>x"8700", 747=>x"9500", 748=>x"9700", 749=>x"8f00",
---- 750=>x"8e00", 751=>x"9700", 752=>x"4300", 753=>x"7300", 754=>x"9000", 755=>x"9600", 756=>x"9500",
---- 757=>x"8e00", 758=>x"9300", 759=>x"9e00", 760=>x"5800", 761=>x"8600", 762=>x"9500", 763=>x"9600",
---- 764=>x"9300", 765=>x"8e00", 766=>x"9700", 767=>x"a100", 768=>x"7100", 769=>x"8f00", 770=>x"9600",
---- 771=>x"9400", 772=>x"9000", 773=>x"9000", 774=>x"9d00", 775=>x"a400", 776=>x"8000", 777=>x"9400",
---- 778=>x"9300", 779=>x"9300", 780=>x"8b00", 781=>x"9200", 782=>x"a200", 783=>x"a500", 784=>x"8f00",
---- 785=>x"9700", 786=>x"9200", 787=>x"9100", 788=>x"8f00", 789=>x"9b00", 790=>x"a400", 791=>x"a700",
---- 792=>x"9200", 793=>x"9300", 794=>x"8f00", 795=>x"8e00", 796=>x"9400", 797=>x"a000", 798=>x"a500",
---- 799=>x"a400", 800=>x"9000", 801=>x"9100", 802=>x"8c00", 803=>x"8d00", 804=>x"9a00", 805=>x"a400",
---- 806=>x"a600", 807=>x"a800", 808=>x"8a00", 809=>x"8a00", 810=>x"8700", 811=>x"8f00", 812=>x"a000",
---- 813=>x"a600", 814=>x"a600", 815=>x"a700", 816=>x"8400", 817=>x"8400", 818=>x"8200", 819=>x"9600",
---- 820=>x"a500", 821=>x"a600", 822=>x"a500", 823=>x"a700", 824=>x"7f00", 825=>x"7b00", 826=>x"8600",
---- 827=>x"9d00", 828=>x"a700", 829=>x"a700", 830=>x"a700", 831=>x"a700", 832=>x"7c00", 833=>x"7c00",
---- 834=>x"8e00", 835=>x"a300", 836=>x"a800", 837=>x"a900", 838=>x"a800", 839=>x"a700", 840=>x"7b00",
---- 841=>x"8000", 842=>x"9400", 843=>x"a500", 844=>x"a900", 845=>x"a700", 846=>x"a700", 847=>x"a700",
---- 848=>x"7a00", 849=>x"8600", 850=>x"9900", 851=>x"a500", 852=>x"a700", 853=>x"a500", 854=>x"a700",
---- 855=>x"a500", 856=>x"7c00", 857=>x"8e00", 858=>x"9b00", 859=>x"a200", 860=>x"a600", 861=>x"a700",
---- 862=>x"a600", 863=>x"a500", 864=>x"8100", 865=>x"9600", 866=>x"a000", 867=>x"a100", 868=>x"a300",
---- 869=>x"a600", 870=>x"a400", 871=>x"a500", 872=>x"8c00", 873=>x"9a00", 874=>x"9b00", 875=>x"9e00",
---- 876=>x"a100", 877=>x"a500", 878=>x"a700", 879=>x"a500", 880=>x"6c00", 881=>x"6600", 882=>x"9600",
---- 883=>x"9600", 884=>x"9b00", 885=>x"a000", 886=>x"a400", 887=>x"a400", 888=>x"9a00", 889=>x"9800",
---- 890=>x"9700", 891=>x"9600", 892=>x"9800", 893=>x"9800", 894=>x"9b00", 895=>x"a000", 896=>x"a100",
---- 897=>x"9b00", 898=>x"9800", 899=>x"9700", 900=>x"9800", 901=>x"9600", 902=>x"9500", 903=>x"9900",
---- 904=>x"a200", 905=>x"9d00", 906=>x"9900", 907=>x"9800", 908=>x"9800", 909=>x"9600", 910=>x"9600",
---- 911=>x"9500", 912=>x"a300", 913=>x"9e00", 914=>x"9a00", 915=>x"9a00", 916=>x"9b00", 917=>x"9700",
---- 918=>x"9900", 919=>x"6700", 920=>x"a500", 921=>x"a100", 922=>x"9f00", 923=>x"9c00", 924=>x"9b00",
---- 925=>x"9900", 926=>x"9800", 927=>x"9800", 928=>x"a400", 929=>x"a300", 930=>x"a400", 931=>x"a200",
---- 932=>x"a000", 933=>x"9d00", 934=>x"9900", 935=>x"9800", 936=>x"a500", 937=>x"a200", 938=>x"a300",
---- 939=>x"a200", 940=>x"a100", 941=>x"9f00", 942=>x"9d00", 943=>x"a000", 944=>x"a000", 945=>x"a200",
---- 946=>x"a200", 947=>x"a400", 948=>x"a000", 949=>x"9e00", 950=>x"a300", 951=>x"a500", 952=>x"a100",
---- 953=>x"a200", 954=>x"a100", 955=>x"a000", 956=>x"9f00", 957=>x"a000", 958=>x"a200", 959=>x"a400",
---- 960=>x"a200", 961=>x"a300", 962=>x"a200", 963=>x"a100", 964=>x"a100", 965=>x"a000", 966=>x"a100",
---- 967=>x"a500", 968=>x"a300", 969=>x"a200", 970=>x"a100", 971=>x"9f00", 972=>x"9f00", 973=>x"a000",
---- 974=>x"a100", 975=>x"a200", 976=>x"a000", 977=>x"a100", 978=>x"a000", 979=>x"a000", 980=>x"9f00",
---- 981=>x"a000", 982=>x"a000", 983=>x"a000", 984=>x"6000", 985=>x"9d00", 986=>x"9e00", 987=>x"9f00",
---- 988=>x"9f00", 989=>x"9d00", 990=>x"9d00", 991=>x"9f00", 992=>x"9e00", 993=>x"9d00", 994=>x"9e00",
---- 995=>x"9f00", 996=>x"9c00", 997=>x"9d00", 998=>x"9c00", 999=>x"a000", 1000=>x"9d00", 1001=>x"9d00",
---- 1002=>x"9e00", 1003=>x"9e00", 1004=>x"9e00", 1005=>x"9e00", 1006=>x"6400", 1007=>x"9b00", 1008=>x"9e00",
---- 1009=>x"9c00", 1010=>x"9c00", 1011=>x"9d00", 1012=>x"9d00", 1013=>x"6400", 1014=>x"9b00", 1015=>x"9c00",
---- 1016=>x"9d00", 1017=>x"9b00", 1018=>x"9c00", 1019=>x"9d00", 1020=>x"9c00", 1021=>x"9c00", 1022=>x"9b00",
---- 1023=>x"9a00", 1024=>x"9c00", 1025=>x"9c00", 1026=>x"9d00", 1027=>x"9c00", 1028=>x"9d00", 1029=>x"9b00",
---- 1030=>x"9a00", 1031=>x"9a00", 1032=>x"9b00", 1033=>x"9b00", 1034=>x"9b00", 1035=>x"9b00", 1036=>x"9d00",
---- 1037=>x"9c00", 1038=>x"9a00", 1039=>x"9b00", 1040=>x"9b00", 1041=>x"6500", 1042=>x"9900", 1043=>x"9800",
---- 1044=>x"9b00", 1045=>x"9b00", 1046=>x"9b00", 1047=>x"9e00", 1048=>x"9900", 1049=>x"9800", 1050=>x"9800",
---- 1051=>x"9a00", 1052=>x"9b00", 1053=>x"9700", 1054=>x"9800", 1055=>x"9d00", 1056=>x"9a00", 1057=>x"9d00",
---- 1058=>x"9800", 1059=>x"9900", 1060=>x"9800", 1061=>x"9900", 1062=>x"9900", 1063=>x"9b00", 1064=>x"9800",
---- 1065=>x"9900", 1066=>x"9900", 1067=>x"9800", 1068=>x"9a00", 1069=>x"9b00", 1070=>x"9800", 1071=>x"9a00",
---- 1072=>x"6600", 1073=>x"6800", 1074=>x"9800", 1075=>x"9700", 1076=>x"9600", 1077=>x"9700", 1078=>x"9700",
---- 1079=>x"9900", 1080=>x"9800", 1081=>x"9700", 1082=>x"9900", 1083=>x"9700", 1084=>x"9900", 1085=>x"9600",
---- 1086=>x"9700", 1087=>x"9a00", 1088=>x"9700", 1089=>x"9900", 1090=>x"9800", 1091=>x"9800", 1092=>x"9f00",
---- 1093=>x"9a00", 1094=>x"9600", 1095=>x"9900", 1096=>x"6a00", 1097=>x"9700", 1098=>x"9800", 1099=>x"9900",
---- 1100=>x"9e00", 1101=>x"a400", 1102=>x"9800", 1103=>x"9a00", 1104=>x"9300", 1105=>x"9700", 1106=>x"9800",
---- 1107=>x"9800", 1108=>x"9f00", 1109=>x"a900", 1110=>x"9900", 1111=>x"9800", 1112=>x"9600", 1113=>x"9500",
---- 1114=>x"9600", 1115=>x"9700", 1116=>x"9a00", 1117=>x"9700", 1118=>x"9500", 1119=>x"9900", 1120=>x"9800",
---- 1121=>x"9700", 1122=>x"9700", 1123=>x"9800", 1124=>x"9600", 1125=>x"9600", 1126=>x"9700", 1127=>x"9800",
---- 1128=>x"9800", 1129=>x"9600", 1130=>x"9700", 1131=>x"9700", 1132=>x"9700", 1133=>x"9400", 1134=>x"9600",
---- 1135=>x"9500", 1136=>x"9800", 1137=>x"9700", 1138=>x"9800", 1139=>x"9700", 1140=>x"9800", 1141=>x"9700",
---- 1142=>x"9600", 1143=>x"9700", 1144=>x"9600", 1145=>x"9800", 1146=>x"9800", 1147=>x"9600", 1148=>x"9700",
---- 1149=>x"9500", 1150=>x"9400", 1151=>x"9700", 1152=>x"9500", 1153=>x"9800", 1154=>x"9900", 1155=>x"9700",
---- 1156=>x"9600", 1157=>x"6c00", 1158=>x"9500", 1159=>x"9700", 1160=>x"9900", 1161=>x"9900", 1162=>x"9700",
---- 1163=>x"9800", 1164=>x"9800", 1165=>x"9400", 1166=>x"9300", 1167=>x"9300", 1168=>x"9600", 1169=>x"9600",
---- 1170=>x"9900", 1171=>x"9900", 1172=>x"9600", 1173=>x"9200", 1174=>x"9300", 1175=>x"9300", 1176=>x"9600",
---- 1177=>x"9600", 1178=>x"9700", 1179=>x"9500", 1180=>x"9500", 1181=>x"9400", 1182=>x"9200", 1183=>x"9200",
---- 1184=>x"9500", 1185=>x"9500", 1186=>x"9600", 1187=>x"9500", 1188=>x"9500", 1189=>x"9300", 1190=>x"9300",
---- 1191=>x"9300", 1192=>x"9600", 1193=>x"6900", 1194=>x"9300", 1195=>x"9200", 1196=>x"9400", 1197=>x"9300",
---- 1198=>x"9400", 1199=>x"9400", 1200=>x"9300", 1201=>x"9600", 1202=>x"9300", 1203=>x"9100", 1204=>x"9500",
---- 1205=>x"9200", 1206=>x"9200", 1207=>x"9400", 1208=>x"9400", 1209=>x"9300", 1210=>x"9200", 1211=>x"9300",
---- 1212=>x"9200", 1213=>x"6f00", 1214=>x"9000", 1215=>x"8e00", 1216=>x"9400", 1217=>x"9000", 1218=>x"9200",
---- 1219=>x"9200", 1220=>x"9200", 1221=>x"9000", 1222=>x"9000", 1223=>x"9300", 1224=>x"9300", 1225=>x"9200",
---- 1226=>x"9300", 1227=>x"9100", 1228=>x"9200", 1229=>x"9000", 1230=>x"8e00", 1231=>x"8f00", 1232=>x"9400",
---- 1233=>x"9400", 1234=>x"9300", 1235=>x"9400", 1236=>x"9300", 1237=>x"9100", 1238=>x"8f00", 1239=>x"9000",
---- 1240=>x"9300", 1241=>x"9300", 1242=>x"9400", 1243=>x"9300", 1244=>x"9200", 1245=>x"9200", 1246=>x"9000",
---- 1247=>x"9000", 1248=>x"9600", 1249=>x"9400", 1250=>x"9600", 1251=>x"9300", 1252=>x"9100", 1253=>x"9100",
---- 1254=>x"8f00", 1255=>x"9100", 1256=>x"9400", 1257=>x"9200", 1258=>x"9400", 1259=>x"9400", 1260=>x"9400",
---- 1261=>x"9300", 1262=>x"9100", 1263=>x"8e00", 1264=>x"9700", 1265=>x"9500", 1266=>x"9400", 1267=>x"9400",
---- 1268=>x"9400", 1269=>x"9200", 1270=>x"9500", 1271=>x"9000", 1272=>x"9600", 1273=>x"9500", 1274=>x"9200",
---- 1275=>x"9400", 1276=>x"9300", 1277=>x"9100", 1278=>x"9300", 1279=>x"9100", 1280=>x"9300", 1281=>x"9500",
---- 1282=>x"9500", 1283=>x"6a00", 1284=>x"6c00", 1285=>x"9000", 1286=>x"9000", 1287=>x"8e00", 1288=>x"9300",
---- 1289=>x"9300", 1290=>x"9400", 1291=>x"9000", 1292=>x"9000", 1293=>x"9100", 1294=>x"9000", 1295=>x"8e00",
---- 1296=>x"9400", 1297=>x"9100", 1298=>x"9100", 1299=>x"9000", 1300=>x"9000", 1301=>x"9200", 1302=>x"9000",
---- 1303=>x"8d00", 1304=>x"9300", 1305=>x"9100", 1306=>x"6d00", 1307=>x"8f00", 1308=>x"9200", 1309=>x"9000",
---- 1310=>x"8c00", 1311=>x"8e00", 1312=>x"9200", 1313=>x"9100", 1314=>x"9300", 1315=>x"9000", 1316=>x"8f00",
---- 1317=>x"8e00", 1318=>x"8f00", 1319=>x"9100", 1320=>x"9200", 1321=>x"9400", 1322=>x"9100", 1323=>x"9100",
---- 1324=>x"9200", 1325=>x"8e00", 1326=>x"8d00", 1327=>x"8d00", 1328=>x"9200", 1329=>x"9300", 1330=>x"9200",
---- 1331=>x"9100", 1332=>x"9000", 1333=>x"9000", 1334=>x"8e00", 1335=>x"8d00", 1336=>x"9300", 1337=>x"9300",
---- 1338=>x"9400", 1339=>x"9100", 1340=>x"8e00", 1341=>x"8d00", 1342=>x"8c00", 1343=>x"8e00", 1344=>x"9300",
---- 1345=>x"9100", 1346=>x"9000", 1347=>x"9300", 1348=>x"9000", 1349=>x"8e00", 1350=>x"8c00", 1351=>x"8d00",
---- 1352=>x"8f00", 1353=>x"9100", 1354=>x"9200", 1355=>x"9000", 1356=>x"9000", 1357=>x"8d00", 1358=>x"8d00",
---- 1359=>x"8d00", 1360=>x"9100", 1361=>x"6e00", 1362=>x"9200", 1363=>x"9000", 1364=>x"8f00", 1365=>x"8f00",
---- 1366=>x"8a00", 1367=>x"8500", 1368=>x"9100", 1369=>x"9200", 1370=>x"9000", 1371=>x"9100", 1372=>x"9000",
---- 1373=>x"8e00", 1374=>x"8900", 1375=>x"8500", 1376=>x"8f00", 1377=>x"9200", 1378=>x"9100", 1379=>x"9000",
---- 1380=>x"8e00", 1381=>x"8c00", 1382=>x"8b00", 1383=>x"8a00", 1384=>x"9200", 1385=>x"9000", 1386=>x"9000",
---- 1387=>x"8f00", 1388=>x"8d00", 1389=>x"8b00", 1390=>x"8b00", 1391=>x"8800", 1392=>x"9100", 1393=>x"9000",
---- 1394=>x"9000", 1395=>x"8f00", 1396=>x"9000", 1397=>x"8d00", 1398=>x"8b00", 1399=>x"7700", 1400=>x"8f00",
---- 1401=>x"8f00", 1402=>x"9000", 1403=>x"9000", 1404=>x"9100", 1405=>x"8f00", 1406=>x"8a00", 1407=>x"8500",
---- 1408=>x"8f00", 1409=>x"9100", 1410=>x"9100", 1411=>x"9000", 1412=>x"8f00", 1413=>x"8d00", 1414=>x"8900",
---- 1415=>x"8600", 1416=>x"9000", 1417=>x"9200", 1418=>x"9000", 1419=>x"6d00", 1420=>x"9100", 1421=>x"8b00",
---- 1422=>x"8a00", 1423=>x"8500", 1424=>x"9200", 1425=>x"9400", 1426=>x"8f00", 1427=>x"9100", 1428=>x"8e00",
---- 1429=>x"8d00", 1430=>x"8700", 1431=>x"8400", 1432=>x"9300", 1433=>x"9200", 1434=>x"8d00", 1435=>x"9000",
---- 1436=>x"8f00", 1437=>x"8c00", 1438=>x"8700", 1439=>x"8300", 1440=>x"9300", 1441=>x"9000", 1442=>x"9100",
---- 1443=>x"9100", 1444=>x"9200", 1445=>x"8c00", 1446=>x"8600", 1447=>x"8400", 1448=>x"6e00", 1449=>x"8f00",
---- 1450=>x"8e00", 1451=>x"8c00", 1452=>x"8e00", 1453=>x"8a00", 1454=>x"8300", 1455=>x"8400", 1456=>x"9000",
---- 1457=>x"8f00", 1458=>x"8d00", 1459=>x"8d00", 1460=>x"8b00", 1461=>x"8900", 1462=>x"8300", 1463=>x"7f00",
---- 1464=>x"8f00", 1465=>x"9000", 1466=>x"8f00", 1467=>x"8e00", 1468=>x"8e00", 1469=>x"8700", 1470=>x"8300",
---- 1471=>x"7e00", 1472=>x"9000", 1473=>x"8d00", 1474=>x"8e00", 1475=>x"8d00", 1476=>x"8c00", 1477=>x"8700",
---- 1478=>x"8000", 1479=>x"7e00", 1480=>x"9300", 1481=>x"8f00", 1482=>x"8e00", 1483=>x"8c00", 1484=>x"8900",
---- 1485=>x"7a00", 1486=>x"7f00", 1487=>x"7a00", 1488=>x"8f00", 1489=>x"8e00", 1490=>x"8c00", 1491=>x"8b00",
---- 1492=>x"8a00", 1493=>x"8700", 1494=>x"7f00", 1495=>x"7800", 1496=>x"8e00", 1497=>x"8d00", 1498=>x"8c00",
---- 1499=>x"8d00", 1500=>x"8900", 1501=>x"8800", 1502=>x"8000", 1503=>x"7b00", 1504=>x"8e00", 1505=>x"8c00",
---- 1506=>x"8c00", 1507=>x"8800", 1508=>x"8600", 1509=>x"8500", 1510=>x"8100", 1511=>x"7d00", 1512=>x"8d00",
---- 1513=>x"8b00", 1514=>x"8c00", 1515=>x"8b00", 1516=>x"8800", 1517=>x"8400", 1518=>x"8000", 1519=>x"7900",
---- 1520=>x"8c00", 1521=>x"8800", 1522=>x"8a00", 1523=>x"8900", 1524=>x"8600", 1525=>x"8200", 1526=>x"7e00",
---- 1527=>x"7700", 1528=>x"8a00", 1529=>x"8b00", 1530=>x"8900", 1531=>x"8900", 1532=>x"8700", 1533=>x"8100",
---- 1534=>x"7e00", 1535=>x"7800", 1536=>x"8d00", 1537=>x"8b00", 1538=>x"8700", 1539=>x"8700", 1540=>x"8800",
---- 1541=>x"8000", 1542=>x"7a00", 1543=>x"7400", 1544=>x"8d00", 1545=>x"8800", 1546=>x"8500", 1547=>x"8500",
---- 1548=>x"8200", 1549=>x"7c00", 1550=>x"8700", 1551=>x"7200", 1552=>x"8900", 1553=>x"8700", 1554=>x"8700",
---- 1555=>x"8300", 1556=>x"8000", 1557=>x"7d00", 1558=>x"7500", 1559=>x"7000", 1560=>x"8900", 1561=>x"8a00",
---- 1562=>x"8700", 1563=>x"8100", 1564=>x"7d00", 1565=>x"7900", 1566=>x"7500", 1567=>x"7100", 1568=>x"8700",
---- 1569=>x"8700", 1570=>x"8600", 1571=>x"8200", 1572=>x"7e00", 1573=>x"7a00", 1574=>x"7500", 1575=>x"8c00",
---- 1576=>x"8100", 1577=>x"8000", 1578=>x"8100", 1579=>x"7f00", 1580=>x"7d00", 1581=>x"7a00", 1582=>x"7400",
---- 1583=>x"7300", 1584=>x"7300", 1585=>x"7300", 1586=>x"7400", 1587=>x"7300", 1588=>x"7500", 1589=>x"8e00",
---- 1590=>x"6d00", 1591=>x"7100", 1592=>x"9900", 1593=>x"6800", 1594=>x"6a00", 1595=>x"6d00", 1596=>x"6c00",
---- 1597=>x"6300", 1598=>x"6000", 1599=>x"6600", 1600=>x"5f00", 1601=>x"6000", 1602=>x"6c00", 1603=>x"6f00",
---- 1604=>x"6b00", 1605=>x"5d00", 1606=>x"4e00", 1607=>x"5600", 1608=>x"5b00", 1609=>x"6400", 1610=>x"7600",
---- 1611=>x"7700", 1612=>x"7200", 1613=>x"6100", 1614=>x"4c00", 1615=>x"4e00", 1616=>x"6200", 1617=>x"6d00",
---- 1618=>x"7f00", 1619=>x"8000", 1620=>x"7400", 1621=>x"6500", 1622=>x"4b00", 1623=>x"5000", 1624=>x"6400",
---- 1625=>x"7400", 1626=>x"8100", 1627=>x"8600", 1628=>x"7600", 1629=>x"6300", 1630=>x"4d00", 1631=>x"5f00",
---- 1632=>x"6b00", 1633=>x"7600", 1634=>x"8300", 1635=>x"8700", 1636=>x"8700", 1637=>x"6500", 1638=>x"5500",
---- 1639=>x"7900", 1640=>x"7100", 1641=>x"7c00", 1642=>x"8100", 1643=>x"8300", 1644=>x"7800", 1645=>x"6c00",
---- 1646=>x"6200", 1647=>x"8d00", 1648=>x"7500", 1649=>x"7c00", 1650=>x"7e00", 1651=>x"8500", 1652=>x"8000",
---- 1653=>x"7100", 1654=>x"6f00", 1655=>x"9d00", 1656=>x"7900", 1657=>x"7c00", 1658=>x"8500", 1659=>x"8400",
---- 1660=>x"8000", 1661=>x"7600", 1662=>x"7e00", 1663=>x"af00", 1664=>x"7d00", 1665=>x"8300", 1666=>x"8900",
---- 1667=>x"8900", 1668=>x"8300", 1669=>x"7900", 1670=>x"8b00", 1671=>x"bd00", 1672=>x"7e00", 1673=>x"8700",
---- 1674=>x"8a00", 1675=>x"8b00", 1676=>x"8900", 1677=>x"7f00", 1678=>x"9600", 1679=>x"c200", 1680=>x"7d00",
---- 1681=>x"8400", 1682=>x"8700", 1683=>x"8900", 1684=>x"8b00", 1685=>x"8700", 1686=>x"a300", 1687=>x"c600",
---- 1688=>x"7900", 1689=>x"7d00", 1690=>x"8b00", 1691=>x"9700", 1692=>x"9e00", 1693=>x"a400", 1694=>x"b500",
---- 1695=>x"c700", 1696=>x"7a00", 1697=>x"8600", 1698=>x"9800", 1699=>x"a500", 1700=>x"b300", 1701=>x"bc00",
---- 1702=>x"c700", 1703=>x"cd00", 1704=>x"8200", 1705=>x"9900", 1706=>x"aa00", 1707=>x"b800", 1708=>x"c000",
---- 1709=>x"c400", 1710=>x"ca00", 1711=>x"d100", 1712=>x"9600", 1713=>x"ad00", 1714=>x"bc00", 1715=>x"c600",
---- 1716=>x"c700", 1717=>x"ca00", 1718=>x"cf00", 1719=>x"d600", 1720=>x"ae00", 1721=>x"c300", 1722=>x"ca00",
---- 1723=>x"cb00", 1724=>x"c900", 1725=>x"cb00", 1726=>x"cf00", 1727=>x"d600", 1728=>x"c100", 1729=>x"2f00",
---- 1730=>x"d400", 1731=>x"d200", 1732=>x"ce00", 1733=>x"cb00", 1734=>x"cd00", 1735=>x"d500", 1736=>x"ce00",
---- 1737=>x"d600", 1738=>x"d900", 1739=>x"d800", 1740=>x"d100", 1741=>x"cf00", 1742=>x"d100", 1743=>x"d400",
---- 1744=>x"d300", 1745=>x"d900", 1746=>x"db00", 1747=>x"d700", 1748=>x"d200", 1749=>x"d200", 1750=>x"d400",
---- 1751=>x"d700", 1752=>x"d300", 1753=>x"da00", 1754=>x"d900", 1755=>x"d500", 1756=>x"d000", 1757=>x"d000",
---- 1758=>x"d500", 1759=>x"d800", 1760=>x"d500", 1761=>x"d800", 1762=>x"d600", 1763=>x"d000", 1764=>x"ce00",
---- 1765=>x"d100", 1766=>x"d500", 1767=>x"da00", 1768=>x"d400", 1769=>x"d700", 1770=>x"d300", 1771=>x"cd00",
---- 1772=>x"cc00", 1773=>x"d100", 1774=>x"d500", 1775=>x"2400", 1776=>x"d400", 1777=>x"d700", 1778=>x"d300",
---- 1779=>x"cd00", 1780=>x"cc00", 1781=>x"d100", 1782=>x"2900", 1783=>x"da00", 1784=>x"d300", 1785=>x"d900",
---- 1786=>x"d200", 1787=>x"ca00", 1788=>x"cc00", 1789=>x"d000", 1790=>x"d800", 1791=>x"dc00", 1792=>x"d000",
---- 1793=>x"d500", 1794=>x"d100", 1795=>x"cb00", 1796=>x"ca00", 1797=>x"d100", 1798=>x"d800", 1799=>x"db00",
---- 1800=>x"c900", 1801=>x"cd00", 1802=>x"cc00", 1803=>x"ca00", 1804=>x"ca00", 1805=>x"d200", 1806=>x"da00",
---- 1807=>x"db00", 1808=>x"b600", 1809=>x"bf00", 1810=>x"bf00", 1811=>x"c100", 1812=>x"c900", 1813=>x"d600",
---- 1814=>x"db00", 1815=>x"d900", 1816=>x"9700", 1817=>x"a600", 1818=>x"a900", 1819=>x"b300", 1820=>x"c900",
---- 1821=>x"d400", 1822=>x"db00", 1823=>x"d700", 1824=>x"8500", 1825=>x"8c00", 1826=>x"9500", 1827=>x"b100",
---- 1828=>x"cc00", 1829=>x"d800", 1830=>x"dc00", 1831=>x"d800", 1832=>x"8400", 1833=>x"8700", 1834=>x"9400",
---- 1835=>x"b600", 1836=>x"cf00", 1837=>x"dc00", 1838=>x"dc00", 1839=>x"d700", 1840=>x"8700", 1841=>x"8b00",
---- 1842=>x"9900", 1843=>x"be00", 1844=>x"d300", 1845=>x"dd00", 1846=>x"dc00", 1847=>x"d500", 1848=>x"8500",
---- 1849=>x"8d00", 1850=>x"a600", 1851=>x"3700", 1852=>x"d500", 1853=>x"dc00", 1854=>x"da00", 1855=>x"d100",
---- 1856=>x"8100", 1857=>x"9200", 1858=>x"b600", 1859=>x"cf00", 1860=>x"d800", 1861=>x"de00", 1862=>x"2700",
---- 1863=>x"ce00", 1864=>x"8c00", 1865=>x"9600", 1866=>x"bc00", 1867=>x"d300", 1868=>x"da00", 1869=>x"dc00",
---- 1870=>x"d500", 1871=>x"c500", 1872=>x"9500", 1873=>x"a400", 1874=>x"c400", 1875=>x"d500", 1876=>x"dc00",
---- 1877=>x"da00", 1878=>x"3000", 1879=>x"b800", 1880=>x"9700", 1881=>x"b300", 1882=>x"cb00", 1883=>x"d700",
---- 1884=>x"2500", 1885=>x"d500", 1886=>x"c900", 1887=>x"ad00", 1888=>x"a000", 1889=>x"4700", 1890=>x"ce00",
---- 1891=>x"d600", 1892=>x"d900", 1893=>x"d200", 1894=>x"c100", 1895=>x"a100", 1896=>x"a000", 1897=>x"c100",
---- 1898=>x"d100", 1899=>x"d800", 1900=>x"d600", 1901=>x"cd00", 1902=>x"b500", 1903=>x"8c00", 1904=>x"ab00",
---- 1905=>x"c800", 1906=>x"d300", 1907=>x"d600", 1908=>x"d200", 1909=>x"c300", 1910=>x"a000", 1911=>x"6400",
---- 1912=>x"b600", 1913=>x"c800", 1914=>x"cf00", 1915=>x"cf00", 1916=>x"c500", 1917=>x"a800", 1918=>x"7300",
---- 1919=>x"4200", 1920=>x"be00", 1921=>x"c800", 1922=>x"c800", 1923=>x"bf00", 1924=>x"a700", 1925=>x"7700",
---- 1926=>x"4400", 1927=>x"3700", 1928=>x"bf00", 1929=>x"ba00", 1930=>x"b200", 1931=>x"9f00", 1932=>x"7900",
---- 1933=>x"5000", 1934=>x"3800", 1935=>x"3400", 1936=>x"b800", 1937=>x"a200", 1938=>x"8f00", 1939=>x"7200",
---- 1940=>x"5100", 1941=>x"4300", 1942=>x"3500", 1943=>x"3400", 1944=>x"a100", 1945=>x"8000", 1946=>x"5d00",
---- 1947=>x"4b00", 1948=>x"4300", 1949=>x"3b00", 1950=>x"3600", 1951=>x"3c00", 1952=>x"7a00", 1953=>x"a800",
---- 1954=>x"4c00", 1955=>x"4700", 1956=>x"4200", 1957=>x"3e00", 1958=>x"4100", 1959=>x"4800", 1960=>x"5700",
---- 1961=>x"5000", 1962=>x"5500", 1963=>x"5000", 1964=>x"4800", 1965=>x"4700", 1966=>x"4d00", 1967=>x"4b00",
---- 1968=>x"5200", 1969=>x"4c00", 1970=>x"4c00", 1971=>x"4c00", 1972=>x"4f00", 1973=>x"5400", 1974=>x"5100",
---- 1975=>x"4f00", 1976=>x"5500", 1977=>x"5500", 1978=>x"5400", 1979=>x"5900", 1980=>x"5b00", 1981=>x"5600",
---- 1982=>x"aa00", 1983=>x"4e00", 1984=>x"5b00", 1985=>x"9f00", 1986=>x"6000", 1987=>x"6400", 1988=>x"5f00",
---- 1989=>x"5600", 1990=>x"5500", 1991=>x"4c00", 1992=>x"6000", 1993=>x"6900", 1994=>x"9300", 1995=>x"6800",
---- 1996=>x"6100", 1997=>x"5a00", 1998=>x"5300", 1999=>x"4f00", 2000=>x"6b00", 2001=>x"7100", 2002=>x"7100",
---- 2003=>x"6a00", 2004=>x"6100", 2005=>x"5c00", 2006=>x"5300", 2007=>x"5400", 2008=>x"7400", 2009=>x"7600",
---- 2010=>x"7200", 2011=>x"6b00", 2012=>x"6200", 2013=>x"5c00", 2014=>x"5700", 2015=>x"5e00", 2016=>x"7d00",
---- 2017=>x"7a00", 2018=>x"7200", 2019=>x"9600", 2020=>x"6000", 2021=>x"5e00", 2022=>x"5f00", 2023=>x"6600",
---- 2024=>x"8100", 2025=>x"7b00", 2026=>x"7000", 2027=>x"6600", 2028=>x"5d00", 2029=>x"5d00", 2030=>x"a100",
---- 2031=>x"6300", 2032=>x"7d00", 2033=>x"7700", 2034=>x"6f00", 2035=>x"6100", 2036=>x"6000", 2037=>x"a200",
---- 2038=>x"5900", 2039=>x"5900", 2040=>x"7d00", 2041=>x"7400", 2042=>x"6500", 2043=>x"5900", 2044=>x"5c00",
---- 2045=>x"5700", 2046=>x"4f00", 2047=>x"4c00"),
---- 28 => (0=>x"7900", 1=>x"7e00", 2=>x"7a00", 3=>x"7800", 4=>x"7800", 5=>x"7a00", 6=>x"7900", 7=>x"7a00",
---- 8=>x"7900", 9=>x"7f00", 10=>x"7a00", 11=>x"7800", 12=>x"7800", 13=>x"7a00", 14=>x"7900",
---- 15=>x"7a00", 16=>x"7b00", 17=>x"7c00", 18=>x"7a00", 19=>x"7700", 20=>x"7800", 21=>x"7a00",
---- 22=>x"7800", 23=>x"7a00", 24=>x"7a00", 25=>x"7c00", 26=>x"7a00", 27=>x"7800", 28=>x"7a00",
---- 29=>x"7900", 30=>x"7900", 31=>x"7c00", 32=>x"7700", 33=>x"7900", 34=>x"7b00", 35=>x"7a00",
---- 36=>x"7800", 37=>x"7800", 38=>x"7b00", 39=>x"7c00", 40=>x"7900", 41=>x"7a00", 42=>x"7800",
---- 43=>x"7900", 44=>x"7700", 45=>x"7800", 46=>x"7800", 47=>x"7800", 48=>x"7900", 49=>x"7a00",
---- 50=>x"7800", 51=>x"7900", 52=>x"7a00", 53=>x"7500", 54=>x"7800", 55=>x"7900", 56=>x"7700",
---- 57=>x"7700", 58=>x"7c00", 59=>x"7a00", 60=>x"7800", 61=>x"7800", 62=>x"7900", 63=>x"7a00",
---- 64=>x"7800", 65=>x"7700", 66=>x"7a00", 67=>x"7800", 68=>x"7700", 69=>x"7c00", 70=>x"7900",
---- 71=>x"7b00", 72=>x"7700", 73=>x"7a00", 74=>x"7c00", 75=>x"8500", 76=>x"7c00", 77=>x"7f00",
---- 78=>x"7a00", 79=>x"7b00", 80=>x"7600", 81=>x"7a00", 82=>x"7900", 83=>x"7b00", 84=>x"7a00",
---- 85=>x"7900", 86=>x"7900", 87=>x"7b00", 88=>x"7500", 89=>x"7400", 90=>x"7200", 91=>x"7a00",
---- 92=>x"7a00", 93=>x"7900", 94=>x"7900", 95=>x"7800", 96=>x"7700", 97=>x"7900", 98=>x"7800",
---- 99=>x"7800", 100=>x"7a00", 101=>x"7a00", 102=>x"7a00", 103=>x"7800", 104=>x"7a00", 105=>x"7b00",
---- 106=>x"7c00", 107=>x"7b00", 108=>x"8400", 109=>x"7c00", 110=>x"7a00", 111=>x"7900", 112=>x"7700",
---- 113=>x"7900", 114=>x"7900", 115=>x"7a00", 116=>x"7b00", 117=>x"7a00", 118=>x"7900", 119=>x"7a00",
---- 120=>x"7300", 121=>x"7400", 122=>x"7500", 123=>x"7a00", 124=>x"7b00", 125=>x"7700", 126=>x"7a00",
---- 127=>x"7800", 128=>x"7300", 129=>x"7700", 130=>x"7500", 131=>x"7800", 132=>x"7900", 133=>x"7a00",
---- 134=>x"7900", 135=>x"7900", 136=>x"7000", 137=>x"7200", 138=>x"7400", 139=>x"7500", 140=>x"7800",
---- 141=>x"7b00", 142=>x"7b00", 143=>x"7900", 144=>x"6c00", 145=>x"7200", 146=>x"7300", 147=>x"7300",
---- 148=>x"7700", 149=>x"7b00", 150=>x"7b00", 151=>x"7d00", 152=>x"6b00", 153=>x"6e00", 154=>x"7000",
---- 155=>x"7200", 156=>x"7400", 157=>x"7900", 158=>x"7700", 159=>x"7d00", 160=>x"6a00", 161=>x"6e00",
---- 162=>x"6b00", 163=>x"7200", 164=>x"7300", 165=>x"7300", 166=>x"7600", 167=>x"7b00", 168=>x"6300",
---- 169=>x"6b00", 170=>x"6b00", 171=>x"6e00", 172=>x"6f00", 173=>x"7000", 174=>x"7400", 175=>x"7900",
---- 176=>x"6200", 177=>x"6800", 178=>x"6a00", 179=>x"6c00", 180=>x"7200", 181=>x"7100", 182=>x"7700",
---- 183=>x"7c00", 184=>x"6e00", 185=>x"6a00", 186=>x"6f00", 187=>x"6d00", 188=>x"7500", 189=>x"7300",
---- 190=>x"7b00", 191=>x"7d00", 192=>x"9200", 193=>x"6c00", 194=>x"6c00", 195=>x"6e00", 196=>x"7300",
---- 197=>x"7900", 198=>x"7a00", 199=>x"6d00", 200=>x"b600", 201=>x"7f00", 202=>x"6a00", 203=>x"7300",
---- 204=>x"7800", 205=>x"7b00", 206=>x"6a00", 207=>x"4800", 208=>x"cd00", 209=>x"a400", 210=>x"7600",
---- 211=>x"7400", 212=>x"7900", 213=>x"7200", 214=>x"4b00", 215=>x"d000", 216=>x"da00", 217=>x"c600",
---- 218=>x"9000", 219=>x"7800", 220=>x"7200", 221=>x"5200", 222=>x"3200", 223=>x"2900", 224=>x"e100",
---- 225=>x"d800", 226=>x"b500", 227=>x"7a00", 228=>x"5300", 229=>x"3000", 230=>x"2b00", 231=>x"2a00",
---- 232=>x"e400", 233=>x"df00", 234=>x"d100", 235=>x"8100", 236=>x"3100", 237=>x"2a00", 238=>x"2900",
---- 239=>x"2900", 240=>x"e400", 241=>x"e400", 242=>x"db00", 243=>x"7700", 244=>x"2000", 245=>x"2800",
---- 246=>x"2800", 247=>x"2900", 248=>x"e600", 249=>x"e400", 250=>x"c100", 251=>x"4600", 252=>x"2100",
---- 253=>x"2900", 254=>x"2a00", 255=>x"2c00", 256=>x"e100", 257=>x"d300", 258=>x"7600", 259=>x"2000",
---- 260=>x"2a00", 261=>x"2700", 262=>x"2800", 263=>x"2b00", 264=>x"d500", 265=>x"9000", 266=>x"3100",
---- 267=>x"2300", 268=>x"2800", 269=>x"2b00", 270=>x"2a00", 271=>x"2900", 272=>x"9400", 273=>x"3700",
---- 274=>x"2600", 275=>x"2900", 276=>x"2c00", 277=>x"2c00", 278=>x"2d00", 279=>x"2c00", 280=>x"3700",
---- 281=>x"2800", 282=>x"2f00", 283=>x"2c00", 284=>x"2c00", 285=>x"2b00", 286=>x"2c00", 287=>x"2e00",
---- 288=>x"2a00", 289=>x"2e00", 290=>x"3000", 291=>x"2a00", 292=>x"2b00", 293=>x"2e00", 294=>x"3100",
---- 295=>x"3100", 296=>x"2e00", 297=>x"2c00", 298=>x"2a00", 299=>x"2c00", 300=>x"d600", 301=>x"2c00",
---- 302=>x"3100", 303=>x"3900", 304=>x"2a00", 305=>x"2b00", 306=>x"2e00", 307=>x"2900", 308=>x"2900",
---- 309=>x"3100", 310=>x"3400", 311=>x"3500", 312=>x"3000", 313=>x"2700", 314=>x"2d00", 315=>x"2d00",
---- 316=>x"2c00", 317=>x"3300", 318=>x"3300", 319=>x"3400", 320=>x"2b00", 321=>x"2a00", 322=>x"3200",
---- 323=>x"3000", 324=>x"2f00", 325=>x"3700", 326=>x"3200", 327=>x"3400", 328=>x"2b00", 329=>x"2c00",
---- 330=>x"2e00", 331=>x"3000", 332=>x"3300", 333=>x"3600", 334=>x"3500", 335=>x"3300", 336=>x"2f00",
---- 337=>x"2d00", 338=>x"3300", 339=>x"3400", 340=>x"3700", 341=>x"3400", 342=>x"3600", 343=>x"3400",
---- 344=>x"2b00", 345=>x"3000", 346=>x"3700", 347=>x"3800", 348=>x"3700", 349=>x"3700", 350=>x"3500",
---- 351=>x"3500", 352=>x"3300", 353=>x"3b00", 354=>x"3900", 355=>x"3500", 356=>x"3500", 357=>x"3600",
---- 358=>x"3400", 359=>x"3200", 360=>x"3a00", 361=>x"3800", 362=>x"3400", 363=>x"3700", 364=>x"3800",
---- 365=>x"3500", 366=>x"3100", 367=>x"2e00", 368=>x"3400", 369=>x"3400", 370=>x"3200", 371=>x"3400",
---- 372=>x"3600", 373=>x"3400", 374=>x"2e00", 375=>x"2d00", 376=>x"ca00", 377=>x"3400", 378=>x"3800",
---- 379=>x"3700", 380=>x"3100", 381=>x"2c00", 382=>x"2800", 383=>x"2a00", 384=>x"3900", 385=>x"3200",
---- 386=>x"3600", 387=>x"3100", 388=>x"2e00", 389=>x"2900", 390=>x"2800", 391=>x"3200", 392=>x"3600",
---- 393=>x"3400", 394=>x"3400", 395=>x"2f00", 396=>x"2b00", 397=>x"2d00", 398=>x"2e00", 399=>x"3a00",
---- 400=>x"3800", 401=>x"3500", 402=>x"3400", 403=>x"3200", 404=>x"2700", 405=>x"2b00", 406=>x"3600",
---- 407=>x"3a00", 408=>x"3500", 409=>x"3800", 410=>x"ce00", 411=>x"2e00", 412=>x"d200", 413=>x"3100",
---- 414=>x"3900", 415=>x"3c00", 416=>x"3b00", 417=>x"3700", 418=>x"2f00", 419=>x"2c00", 420=>x"3200",
---- 421=>x"3800", 422=>x"3500", 423=>x"2d00", 424=>x"3700", 425=>x"3300", 426=>x"2f00", 427=>x"2d00",
---- 428=>x"3400", 429=>x"3900", 430=>x"3200", 431=>x"2d00", 432=>x"3600", 433=>x"2e00", 434=>x"2e00",
---- 435=>x"3500", 436=>x"c800", 437=>x"3700", 438=>x"3100", 439=>x"2f00", 440=>x"3300", 441=>x"3000",
---- 442=>x"3300", 443=>x"3600", 444=>x"3700", 445=>x"3300", 446=>x"2f00", 447=>x"3100", 448=>x"3400",
---- 449=>x"3500", 450=>x"3200", 451=>x"3600", 452=>x"3300", 453=>x"2d00", 454=>x"3100", 455=>x"3800",
---- 456=>x"3200", 457=>x"3800", 458=>x"3600", 459=>x"3200", 460=>x"2f00", 461=>x"2f00", 462=>x"3200",
---- 463=>x"3700", 464=>x"3600", 465=>x"3500", 466=>x"3800", 467=>x"3400", 468=>x"2f00", 469=>x"3200",
---- 470=>x"3900", 471=>x"4000", 472=>x"3400", 473=>x"3500", 474=>x"3500", 475=>x"3200", 476=>x"3100",
---- 477=>x"3400", 478=>x"3800", 479=>x"3800", 480=>x"3300", 481=>x"3400", 482=>x"2e00", 483=>x"2e00",
---- 484=>x"3600", 485=>x"3700", 486=>x"3500", 487=>x"3600", 488=>x"3700", 489=>x"d000", 490=>x"2f00",
---- 491=>x"3000", 492=>x"3200", 493=>x"3500", 494=>x"3600", 495=>x"3400", 496=>x"2a00", 497=>x"2800",
---- 498=>x"3300", 499=>x"3100", 500=>x"3700", 501=>x"3800", 502=>x"3700", 503=>x"3600", 504=>x"2800",
---- 505=>x"2e00", 506=>x"3300", 507=>x"3000", 508=>x"3700", 509=>x"3800", 510=>x"3500", 511=>x"3000",
---- 512=>x"d200", 513=>x"2e00", 514=>x"3100", 515=>x"3300", 516=>x"3500", 517=>x"3200", 518=>x"2e00",
---- 519=>x"2c00", 520=>x"3200", 521=>x"3300", 522=>x"3400", 523=>x"3300", 524=>x"3200", 525=>x"2700",
---- 526=>x"2300", 527=>x"3000", 528=>x"3500", 529=>x"3700", 530=>x"3600", 531=>x"3700", 532=>x"2a00",
---- 533=>x"2100", 534=>x"2200", 535=>x"3b00", 536=>x"3300", 537=>x"3400", 538=>x"3600", 539=>x"3400",
---- 540=>x"2600", 541=>x"1f00", 542=>x"2a00", 543=>x"5b00", 544=>x"3300", 545=>x"3500", 546=>x"3500",
---- 547=>x"3000", 548=>x"2300", 549=>x"2400", 550=>x"4100", 551=>x"7400", 552=>x"3400", 553=>x"3200",
---- 554=>x"3000", 555=>x"2d00", 556=>x"2c00", 557=>x"3b00", 558=>x"6300", 559=>x"8a00", 560=>x"3400",
---- 561=>x"3500", 562=>x"3600", 563=>x"ca00", 564=>x"c500", 565=>x"5500", 566=>x"7d00", 567=>x"9400",
---- 568=>x"3300", 569=>x"3700", 570=>x"3c00", 571=>x"4100", 572=>x"4900", 573=>x"6800", 574=>x"8e00",
---- 575=>x"9600", 576=>x"3200", 577=>x"3600", 578=>x"3f00", 579=>x"4400", 580=>x"5d00", 581=>x"8100",
---- 582=>x"9500", 583=>x"9800", 584=>x"3b00", 585=>x"4000", 586=>x"4600", 587=>x"5700", 588=>x"7700",
---- 589=>x"9000", 590=>x"9900", 591=>x"9500", 592=>x"3500", 593=>x"3900", 594=>x"4c00", 595=>x"6900",
---- 596=>x"8700", 597=>x"9800", 598=>x"9800", 599=>x"9400", 600=>x"2c00", 601=>x"3b00", 602=>x"5c00",
---- 603=>x"7f00", 604=>x"9300", 605=>x"9800", 606=>x"9600", 607=>x"9000", 608=>x"2700", 609=>x"4000",
---- 610=>x"6d00", 611=>x"8e00", 612=>x"9a00", 613=>x"6800", 614=>x"9100", 615=>x"9100", 616=>x"3000",
---- 617=>x"5400", 618=>x"8000", 619=>x"9700", 620=>x"9b00", 621=>x"9400", 622=>x"9000", 623=>x"9300",
---- 624=>x"4700", 625=>x"6e00", 626=>x"8e00", 627=>x"9900", 628=>x"9700", 629=>x"9300", 630=>x"9100",
---- 631=>x"9800", 632=>x"6300", 633=>x"7b00", 634=>x"9500", 635=>x"9700", 636=>x"9300", 637=>x"8e00",
---- 638=>x"9300", 639=>x"9b00", 640=>x"7b00", 641=>x"9200", 642=>x"9700", 643=>x"9500", 644=>x"9100",
---- 645=>x"9200", 646=>x"9600", 647=>x"9f00", 648=>x"8c00", 649=>x"9c00", 650=>x"9800", 651=>x"9200",
---- 652=>x"9100", 653=>x"9400", 654=>x"9d00", 655=>x"a000", 656=>x"9600", 657=>x"9b00", 658=>x"9400",
---- 659=>x"9100", 660=>x"9100", 661=>x"9600", 662=>x"9c00", 663=>x"9f00", 664=>x"9a00", 665=>x"9800",
---- 666=>x"9100", 667=>x"8e00", 668=>x"9500", 669=>x"6200", 670=>x"9e00", 671=>x"9f00", 672=>x"9900",
---- 673=>x"9400", 674=>x"9400", 675=>x"8e00", 676=>x"9800", 677=>x"9d00", 678=>x"9e00", 679=>x"9f00",
---- 680=>x"9500", 681=>x"9300", 682=>x"9100", 683=>x"9400", 684=>x"9c00", 685=>x"9f00", 686=>x"a000",
---- 687=>x"a100", 688=>x"9200", 689=>x"9100", 690=>x"9300", 691=>x"9900", 692=>x"9c00", 693=>x"a000",
---- 694=>x"9e00", 695=>x"a200", 696=>x"9300", 697=>x"9100", 698=>x"9600", 699=>x"9e00", 700=>x"a100",
---- 701=>x"9f00", 702=>x"9f00", 703=>x"a100", 704=>x"9000", 705=>x"9300", 706=>x"9900", 707=>x"9f00",
---- 708=>x"a200", 709=>x"a100", 710=>x"9f00", 711=>x"9e00", 712=>x"8e00", 713=>x"9700", 714=>x"a000",
---- 715=>x"a100", 716=>x"a100", 717=>x"a000", 718=>x"a200", 719=>x"a000", 720=>x"6f00", 721=>x"9c00",
---- 722=>x"a000", 723=>x"a100", 724=>x"a100", 725=>x"a000", 726=>x"a000", 727=>x"9f00", 728=>x"9800",
---- 729=>x"a000", 730=>x"a300", 731=>x"a100", 732=>x"9f00", 733=>x"a100", 734=>x"a000", 735=>x"9f00",
---- 736=>x"9b00", 737=>x"a300", 738=>x"a300", 739=>x"a100", 740=>x"a400", 741=>x"a100", 742=>x"9f00",
---- 743=>x"a300", 744=>x"9f00", 745=>x"a400", 746=>x"a400", 747=>x"a200", 748=>x"a200", 749=>x"a100",
---- 750=>x"9e00", 751=>x"9f00", 752=>x"a500", 753=>x"a600", 754=>x"a400", 755=>x"a300", 756=>x"a200",
---- 757=>x"a300", 758=>x"9f00", 759=>x"a000", 760=>x"a400", 761=>x"a500", 762=>x"a400", 763=>x"a200",
---- 764=>x"a000", 765=>x"a200", 766=>x"a100", 767=>x"a200", 768=>x"a500", 769=>x"a400", 770=>x"a400",
---- 771=>x"a300", 772=>x"a200", 773=>x"5b00", 774=>x"a300", 775=>x"a100", 776=>x"a300", 777=>x"a400",
---- 778=>x"a600", 779=>x"a500", 780=>x"a700", 781=>x"a500", 782=>x"a200", 783=>x"a100", 784=>x"a400",
---- 785=>x"a400", 786=>x"a400", 787=>x"a500", 788=>x"a600", 789=>x"a300", 790=>x"a200", 791=>x"a200",
---- 792=>x"a700", 793=>x"a600", 794=>x"a400", 795=>x"a600", 796=>x"a800", 797=>x"a300", 798=>x"a300",
---- 799=>x"a300", 800=>x"a400", 801=>x"a600", 802=>x"a500", 803=>x"a500", 804=>x"a500", 805=>x"a500",
---- 806=>x"a400", 807=>x"a300", 808=>x"a400", 809=>x"a400", 810=>x"5900", 811=>x"a600", 812=>x"a400",
---- 813=>x"a100", 814=>x"a100", 815=>x"a400", 816=>x"a600", 817=>x"a500", 818=>x"a100", 819=>x"a500",
---- 820=>x"a400", 821=>x"a200", 822=>x"a000", 823=>x"a400", 824=>x"a400", 825=>x"a400", 826=>x"a200",
---- 827=>x"a300", 828=>x"a400", 829=>x"a200", 830=>x"a100", 831=>x"a400", 832=>x"a300", 833=>x"a200",
---- 834=>x"a200", 835=>x"a300", 836=>x"a400", 837=>x"a300", 838=>x"a300", 839=>x"a400", 840=>x"a600",
---- 841=>x"a200", 842=>x"a400", 843=>x"a300", 844=>x"a200", 845=>x"a400", 846=>x"a400", 847=>x"a400",
---- 848=>x"a600", 849=>x"a400", 850=>x"a600", 851=>x"a300", 852=>x"a200", 853=>x"a300", 854=>x"a300",
---- 855=>x"a400", 856=>x"a500", 857=>x"a700", 858=>x"a500", 859=>x"a200", 860=>x"a400", 861=>x"a300",
---- 862=>x"a200", 863=>x"a400", 864=>x"a200", 865=>x"a500", 866=>x"a300", 867=>x"a300", 868=>x"a200",
---- 869=>x"a100", 870=>x"a300", 871=>x"a300", 872=>x"a400", 873=>x"a500", 874=>x"a600", 875=>x"a500",
---- 876=>x"a200", 877=>x"a100", 878=>x"9e00", 879=>x"a100", 880=>x"a600", 881=>x"a700", 882=>x"a600",
---- 883=>x"a500", 884=>x"a400", 885=>x"a300", 886=>x"a100", 887=>x"a200", 888=>x"9f00", 889=>x"a300",
---- 890=>x"a500", 891=>x"a200", 892=>x"a200", 893=>x"a300", 894=>x"a300", 895=>x"a300", 896=>x"9a00",
---- 897=>x"9a00", 898=>x"9e00", 899=>x"9e00", 900=>x"a100", 901=>x"9f00", 902=>x"9f00", 903=>x"a100",
---- 904=>x"9500", 905=>x"9700", 906=>x"9600", 907=>x"9800", 908=>x"9a00", 909=>x"9b00", 910=>x"9e00",
---- 911=>x"a000", 912=>x"9700", 913=>x"9600", 914=>x"9400", 915=>x"9600", 916=>x"9800", 917=>x"9700",
---- 918=>x"9600", 919=>x"9900", 920=>x"9700", 921=>x"9500", 922=>x"9400", 923=>x"9300", 924=>x"9400",
---- 925=>x"9700", 926=>x"9600", 927=>x"9600", 928=>x"9600", 929=>x"9800", 930=>x"9700", 931=>x"9600",
---- 932=>x"9600", 933=>x"9700", 934=>x"9400", 935=>x"9300", 936=>x"9e00", 937=>x"9c00", 938=>x"9a00",
---- 939=>x"9a00", 940=>x"9900", 941=>x"9900", 942=>x"9900", 943=>x"9500", 944=>x"a200", 945=>x"9f00",
---- 946=>x"a100", 947=>x"9e00", 948=>x"9d00", 949=>x"9c00", 950=>x"9900", 951=>x"9b00", 952=>x"a300",
---- 953=>x"a300", 954=>x"a400", 955=>x"a400", 956=>x"a000", 957=>x"9e00", 958=>x"9b00", 959=>x"9c00",
---- 960=>x"a500", 961=>x"a600", 962=>x"5a00", 963=>x"a500", 964=>x"a500", 965=>x"a000", 966=>x"9e00",
---- 967=>x"9d00", 968=>x"a400", 969=>x"a300", 970=>x"a800", 971=>x"a600", 972=>x"a400", 973=>x"a300",
---- 974=>x"a000", 975=>x"9e00", 976=>x"a300", 977=>x"a300", 978=>x"a200", 979=>x"a400", 980=>x"a400",
---- 981=>x"a300", 982=>x"9f00", 983=>x"9d00", 984=>x"9e00", 985=>x"9f00", 986=>x"a200", 987=>x"a100",
---- 988=>x"a200", 989=>x"a200", 990=>x"a200", 991=>x"9d00", 992=>x"9d00", 993=>x"9e00", 994=>x"9f00",
---- 995=>x"9f00", 996=>x"9e00", 997=>x"a100", 998=>x"a100", 999=>x"9c00", 1000=>x"9b00", 1001=>x"9e00",
---- 1002=>x"9c00", 1003=>x"9e00", 1004=>x"9f00", 1005=>x"9f00", 1006=>x"9f00", 1007=>x"9b00", 1008=>x"9c00",
---- 1009=>x"9c00", 1010=>x"9c00", 1011=>x"9e00", 1012=>x"9d00", 1013=>x"9e00", 1014=>x"9e00", 1015=>x"9c00",
---- 1016=>x"9a00", 1017=>x"9a00", 1018=>x"9d00", 1019=>x"9e00", 1020=>x"9f00", 1021=>x"a000", 1022=>x"6200",
---- 1023=>x"9b00", 1024=>x"9c00", 1025=>x"9c00", 1026=>x"9c00", 1027=>x"9d00", 1028=>x"9e00", 1029=>x"9d00",
---- 1030=>x"9b00", 1031=>x"9b00", 1032=>x"9b00", 1033=>x"9c00", 1034=>x"9c00", 1035=>x"9c00", 1036=>x"9d00",
---- 1037=>x"9d00", 1038=>x"9e00", 1039=>x"9a00", 1040=>x"9a00", 1041=>x"9a00", 1042=>x"9c00", 1043=>x"9a00",
---- 1044=>x"9c00", 1045=>x"9b00", 1046=>x"9a00", 1047=>x"9a00", 1048=>x"9b00", 1049=>x"9900", 1050=>x"9a00",
---- 1051=>x"9d00", 1052=>x"9d00", 1053=>x"9a00", 1054=>x"9a00", 1055=>x"9800", 1056=>x"9900", 1057=>x"9a00",
---- 1058=>x"9b00", 1059=>x"9800", 1060=>x"6600", 1061=>x"9900", 1062=>x"9a00", 1063=>x"9a00", 1064=>x"9800",
---- 1065=>x"9900", 1066=>x"9800", 1067=>x"9600", 1068=>x"9800", 1069=>x"9800", 1070=>x"9800", 1071=>x"9a00",
---- 1072=>x"9900", 1073=>x"9b00", 1074=>x"9800", 1075=>x"9800", 1076=>x"9a00", 1077=>x"6500", 1078=>x"9800",
---- 1079=>x"9700", 1080=>x"9700", 1081=>x"9b00", 1082=>x"9b00", 1083=>x"9600", 1084=>x"9a00", 1085=>x"9800",
---- 1086=>x"9900", 1087=>x"9a00", 1088=>x"9900", 1089=>x"9800", 1090=>x"9a00", 1091=>x"9a00", 1092=>x"9900",
---- 1093=>x"9800", 1094=>x"9800", 1095=>x"9700", 1096=>x"9700", 1097=>x"9800", 1098=>x"9b00", 1099=>x"9900",
---- 1100=>x"9700", 1101=>x"9600", 1102=>x"9500", 1103=>x"9600", 1104=>x"9700", 1105=>x"9a00", 1106=>x"9a00",
---- 1107=>x"9a00", 1108=>x"9b00", 1109=>x"9800", 1110=>x"9700", 1111=>x"9500", 1112=>x"9700", 1113=>x"9500",
---- 1114=>x"9600", 1115=>x"9b00", 1116=>x"9900", 1117=>x"9700", 1118=>x"9700", 1119=>x"9400", 1120=>x"9700",
---- 1121=>x"9600", 1122=>x"9600", 1123=>x"9600", 1124=>x"9700", 1125=>x"9500", 1126=>x"9500", 1127=>x"9400",
---- 1128=>x"9600", 1129=>x"9800", 1130=>x"9600", 1131=>x"9700", 1132=>x"9600", 1133=>x"9300", 1134=>x"9200",
---- 1135=>x"9200", 1136=>x"9500", 1137=>x"9500", 1138=>x"9600", 1139=>x"9600", 1140=>x"9300", 1141=>x"6d00",
---- 1142=>x"9100", 1143=>x"9300", 1144=>x"9500", 1145=>x"9400", 1146=>x"9300", 1147=>x"9300", 1148=>x"9200",
---- 1149=>x"9400", 1150=>x"9100", 1151=>x"8f00", 1152=>x"9600", 1153=>x"9400", 1154=>x"9300", 1155=>x"9100",
---- 1156=>x"8f00", 1157=>x"8f00", 1158=>x"8f00", 1159=>x"8e00", 1160=>x"9300", 1161=>x"9100", 1162=>x"9300",
---- 1163=>x"9200", 1164=>x"8f00", 1165=>x"8e00", 1166=>x"8e00", 1167=>x"8c00", 1168=>x"9400", 1169=>x"9100",
---- 1170=>x"6c00", 1171=>x"9100", 1172=>x"8f00", 1173=>x"8f00", 1174=>x"8b00", 1175=>x"8900", 1176=>x"9000",
---- 1177=>x"9300", 1178=>x"9000", 1179=>x"8e00", 1180=>x"6f00", 1181=>x"9000", 1182=>x"8d00", 1183=>x"8a00",
---- 1184=>x"9000", 1185=>x"9100", 1186=>x"9300", 1187=>x"8f00", 1188=>x"8f00", 1189=>x"8e00", 1190=>x"8b00",
---- 1191=>x"8800", 1192=>x"9100", 1193=>x"9000", 1194=>x"9300", 1195=>x"9100", 1196=>x"8d00", 1197=>x"7200",
---- 1198=>x"8a00", 1199=>x"8800", 1200=>x"9000", 1201=>x"8f00", 1202=>x"8f00", 1203=>x"8f00", 1204=>x"8b00",
---- 1205=>x"8a00", 1206=>x"8500", 1207=>x"8500", 1208=>x"7000", 1209=>x"9100", 1210=>x"6f00", 1211=>x"8e00",
---- 1212=>x"8e00", 1213=>x"8800", 1214=>x"8500", 1215=>x"8300", 1216=>x"9100", 1217=>x"8d00", 1218=>x"9000",
---- 1219=>x"8d00", 1220=>x"8a00", 1221=>x"8800", 1222=>x"8500", 1223=>x"8100", 1224=>x"8f00", 1225=>x"8c00",
---- 1226=>x"8d00", 1227=>x"8a00", 1228=>x"8b00", 1229=>x"8800", 1230=>x"7d00", 1231=>x"8200", 1232=>x"8d00",
---- 1233=>x"8b00", 1234=>x"8900", 1235=>x"8a00", 1236=>x"8800", 1237=>x"8500", 1238=>x"8100", 1239=>x"8900",
---- 1240=>x"8d00", 1241=>x"8900", 1242=>x"8d00", 1243=>x"8c00", 1244=>x"8700", 1245=>x"8500", 1246=>x"8200",
---- 1247=>x"6c00", 1248=>x"8f00", 1249=>x"7500", 1250=>x"8c00", 1251=>x"8a00", 1252=>x"8600", 1253=>x"8200",
---- 1254=>x"8900", 1255=>x"a300", 1256=>x"8f00", 1257=>x"8d00", 1258=>x"8900", 1259=>x"8600", 1260=>x"8400",
---- 1261=>x"8200", 1262=>x"9600", 1263=>x"af00", 1264=>x"8d00", 1265=>x"8a00", 1266=>x"8a00", 1267=>x"8400",
---- 1268=>x"8200", 1269=>x"8800", 1270=>x"a000", 1271=>x"b800", 1272=>x"8f00", 1273=>x"8a00", 1274=>x"8800",
---- 1275=>x"8200", 1276=>x"8200", 1277=>x"9100", 1278=>x"aa00", 1279=>x"bc00", 1280=>x"8c00", 1281=>x"8b00",
---- 1282=>x"8700", 1283=>x"8300", 1284=>x"8500", 1285=>x"9e00", 1286=>x"4c00", 1287=>x"bf00", 1288=>x"8d00",
---- 1289=>x"8b00", 1290=>x"8600", 1291=>x"8100", 1292=>x"8800", 1293=>x"a400", 1294=>x"b600", 1295=>x"c000",
---- 1296=>x"7100", 1297=>x"8800", 1298=>x"8600", 1299=>x"8400", 1300=>x"9100", 1301=>x"aa00", 1302=>x"bc00",
---- 1303=>x"c100", 1304=>x"8d00", 1305=>x"7700", 1306=>x"8700", 1307=>x"8400", 1308=>x"9a00", 1309=>x"af00",
---- 1310=>x"bf00", 1311=>x"c400", 1312=>x"8c00", 1313=>x"8700", 1314=>x"8400", 1315=>x"8800", 1316=>x"a000",
---- 1317=>x"b600", 1318=>x"c100", 1319=>x"c400", 1320=>x"8900", 1321=>x"8600", 1322=>x"8300", 1323=>x"8900",
---- 1324=>x"a500", 1325=>x"b900", 1326=>x"c300", 1327=>x"c400", 1328=>x"8700", 1329=>x"8600", 1330=>x"7a00",
---- 1331=>x"9100", 1332=>x"a900", 1333=>x"bb00", 1334=>x"c300", 1335=>x"c400", 1336=>x"8800", 1337=>x"8300",
---- 1338=>x"8300", 1339=>x"9600", 1340=>x"ab00", 1341=>x"bd00", 1342=>x"c400", 1343=>x"c400", 1344=>x"7500",
---- 1345=>x"8300", 1346=>x"8600", 1347=>x"9a00", 1348=>x"b100", 1349=>x"bf00", 1350=>x"c400", 1351=>x"c400",
---- 1352=>x"8900", 1353=>x"8400", 1354=>x"8600", 1355=>x"9e00", 1356=>x"b500", 1357=>x"c200", 1358=>x"c200",
---- 1359=>x"c500", 1360=>x"8300", 1361=>x"8200", 1362=>x"8600", 1363=>x"a200", 1364=>x"b600", 1365=>x"c400",
---- 1366=>x"c500", 1367=>x"c400", 1368=>x"8300", 1369=>x"8000", 1370=>x"8800", 1371=>x"a300", 1372=>x"b700",
---- 1373=>x"c300", 1374=>x"c400", 1375=>x"c600", 1376=>x"8500", 1377=>x"7f00", 1378=>x"8900", 1379=>x"a600",
---- 1380=>x"b800", 1381=>x"c200", 1382=>x"c600", 1383=>x"ca00", 1384=>x"8400", 1385=>x"7e00", 1386=>x"8b00",
---- 1387=>x"a600", 1388=>x"b900", 1389=>x"c300", 1390=>x"c700", 1391=>x"cb00", 1392=>x"8200", 1393=>x"7d00",
---- 1394=>x"8e00", 1395=>x"5400", 1396=>x"ba00", 1397=>x"c300", 1398=>x"ca00", 1399=>x"ce00", 1400=>x"7f00",
---- 1401=>x"7e00", 1402=>x"9100", 1403=>x"ad00", 1404=>x"bc00", 1405=>x"c600", 1406=>x"cc00", 1407=>x"d100",
---- 1408=>x"8100", 1409=>x"8000", 1410=>x"9500", 1411=>x"af00", 1412=>x"c000", 1413=>x"c900", 1414=>x"cf00",
---- 1415=>x"d300", 1416=>x"7f00", 1417=>x"7f00", 1418=>x"9800", 1419=>x"b300", 1420=>x"c400", 1421=>x"cc00",
---- 1422=>x"d200", 1423=>x"2b00", 1424=>x"7e00", 1425=>x"7f00", 1426=>x"9900", 1427=>x"b500", 1428=>x"c700",
---- 1429=>x"cf00", 1430=>x"d500", 1431=>x"d400", 1432=>x"7d00", 1433=>x"7e00", 1434=>x"9d00", 1435=>x"b800",
---- 1436=>x"ca00", 1437=>x"d300", 1438=>x"d600", 1439=>x"d600", 1440=>x"7c00", 1441=>x"7e00", 1442=>x"6300",
---- 1443=>x"ba00", 1444=>x"cf00", 1445=>x"d400", 1446=>x"d700", 1447=>x"d700", 1448=>x"7a00", 1449=>x"7d00",
---- 1450=>x"9e00", 1451=>x"bf00", 1452=>x"cf00", 1453=>x"d600", 1454=>x"d800", 1455=>x"d700", 1456=>x"7700",
---- 1457=>x"7b00", 1458=>x"9e00", 1459=>x"c000", 1460=>x"d100", 1461=>x"d800", 1462=>x"d900", 1463=>x"d900",
---- 1464=>x"7500", 1465=>x"7700", 1466=>x"9b00", 1467=>x"c300", 1468=>x"d300", 1469=>x"db00", 1470=>x"dc00",
---- 1471=>x"d800", 1472=>x"7900", 1473=>x"7800", 1474=>x"6300", 1475=>x"c300", 1476=>x"d500", 1477=>x"da00",
---- 1478=>x"da00", 1479=>x"da00", 1480=>x"7700", 1481=>x"7400", 1482=>x"9d00", 1483=>x"c800", 1484=>x"d400",
---- 1485=>x"db00", 1486=>x"db00", 1487=>x"db00", 1488=>x"7600", 1489=>x"7600", 1490=>x"a300", 1491=>x"c800",
---- 1492=>x"d500", 1493=>x"db00", 1494=>x"da00", 1495=>x"da00", 1496=>x"7300", 1497=>x"7900", 1498=>x"aa00",
---- 1499=>x"cd00", 1500=>x"d800", 1501=>x"dd00", 1502=>x"da00", 1503=>x"db00", 1504=>x"7300", 1505=>x"7e00",
---- 1506=>x"b300", 1507=>x"2e00", 1508=>x"da00", 1509=>x"2100", 1510=>x"dc00", 1511=>x"db00", 1512=>x"7100",
---- 1513=>x"8200", 1514=>x"b800", 1515=>x"d400", 1516=>x"dc00", 1517=>x"de00", 1518=>x"db00", 1519=>x"d900",
---- 1520=>x"7500", 1521=>x"8c00", 1522=>x"be00", 1523=>x"d500", 1524=>x"dd00", 1525=>x"df00", 1526=>x"db00",
---- 1527=>x"d700", 1528=>x"7400", 1529=>x"9600", 1530=>x"c500", 1531=>x"d600", 1532=>x"dc00", 1533=>x"dd00",
---- 1534=>x"da00", 1535=>x"d800", 1536=>x"7600", 1537=>x"a400", 1538=>x"c900", 1539=>x"d600", 1540=>x"dd00",
---- 1541=>x"dc00", 1542=>x"d800", 1543=>x"d700", 1544=>x"7e00", 1545=>x"b100", 1546=>x"3000", 1547=>x"d900",
---- 1548=>x"db00", 1549=>x"da00", 1550=>x"d600", 1551=>x"d400", 1552=>x"8700", 1553=>x"bc00", 1554=>x"d100",
---- 1555=>x"d900", 1556=>x"db00", 1557=>x"d700", 1558=>x"d200", 1559=>x"d200", 1560=>x"9600", 1561=>x"c400",
---- 1562=>x"d500", 1563=>x"da00", 1564=>x"d900", 1565=>x"d200", 1566=>x"d000", 1567=>x"d200", 1568=>x"9c00",
---- 1569=>x"c800", 1570=>x"d400", 1571=>x"d700", 1572=>x"d600", 1573=>x"cf00", 1574=>x"cf00", 1575=>x"d000",
---- 1576=>x"9f00", 1577=>x"c900", 1578=>x"d200", 1579=>x"d600", 1580=>x"d400", 1581=>x"ce00", 1582=>x"cd00",
---- 1583=>x"ce00", 1584=>x"9f00", 1585=>x"ca00", 1586=>x"d000", 1587=>x"d400", 1588=>x"ce00", 1589=>x"cc00",
---- 1590=>x"cc00", 1591=>x"ce00", 1592=>x"9c00", 1593=>x"3d00", 1594=>x"ce00", 1595=>x"d200", 1596=>x"cf00",
---- 1597=>x"cb00", 1598=>x"cc00", 1599=>x"cf00", 1600=>x"8e00", 1601=>x"c000", 1602=>x"cf00", 1603=>x"d100",
---- 1604=>x"cd00", 1605=>x"cc00", 1606=>x"cd00", 1607=>x"d100", 1608=>x"8a00", 1609=>x"c200", 1610=>x"cf00",
---- 1611=>x"cf00", 1612=>x"cd00", 1613=>x"cc00", 1614=>x"d000", 1615=>x"d400", 1616=>x"9200", 1617=>x"c400",
---- 1618=>x"d100", 1619=>x"d100", 1620=>x"d000", 1621=>x"cf00", 1622=>x"d400", 1623=>x"d600", 1624=>x"a200",
---- 1625=>x"c800", 1626=>x"d000", 1627=>x"d200", 1628=>x"d300", 1629=>x"d200", 1630=>x"d300", 1631=>x"d700",
---- 1632=>x"b300", 1633=>x"cd00", 1634=>x"d300", 1635=>x"d400", 1636=>x"d400", 1637=>x"d400", 1638=>x"d300",
---- 1639=>x"d500", 1640=>x"be00", 1641=>x"cc00", 1642=>x"d400", 1643=>x"d400", 1644=>x"d400", 1645=>x"d400",
---- 1646=>x"d400", 1647=>x"d500", 1648=>x"c500", 1649=>x"d100", 1650=>x"d400", 1651=>x"d400", 1652=>x"d400",
---- 1653=>x"d500", 1654=>x"d500", 1655=>x"d500", 1656=>x"cb00", 1657=>x"d300", 1658=>x"d500", 1659=>x"d500",
---- 1660=>x"d500", 1661=>x"d600", 1662=>x"d600", 1663=>x"d500", 1664=>x"cd00", 1665=>x"d600", 1666=>x"d600",
---- 1667=>x"d400", 1668=>x"d600", 1669=>x"d500", 1670=>x"d400", 1671=>x"d400", 1672=>x"2d00", 1673=>x"d900",
---- 1674=>x"d600", 1675=>x"d400", 1676=>x"d500", 1677=>x"d400", 1678=>x"d500", 1679=>x"d200", 1680=>x"d300",
---- 1681=>x"d900", 1682=>x"d600", 1683=>x"d400", 1684=>x"d700", 1685=>x"d400", 1686=>x"d200", 1687=>x"d200",
---- 1688=>x"d400", 1689=>x"d700", 1690=>x"d600", 1691=>x"d600", 1692=>x"d500", 1693=>x"d300", 1694=>x"d200",
---- 1695=>x"d000", 1696=>x"d400", 1697=>x"d700", 1698=>x"d700", 1699=>x"d700", 1700=>x"d500", 1701=>x"d500",
---- 1702=>x"d000", 1703=>x"cc00", 1704=>x"d600", 1705=>x"d900", 1706=>x"d700", 1707=>x"d600", 1708=>x"d600",
---- 1709=>x"d100", 1710=>x"cf00", 1711=>x"3900", 1712=>x"2700", 1713=>x"d900", 1714=>x"d700", 1715=>x"d700",
---- 1716=>x"d500", 1717=>x"cf00", 1718=>x"cb00", 1719=>x"bd00", 1720=>x"da00", 1721=>x"d700", 1722=>x"d800",
---- 1723=>x"d600", 1724=>x"d600", 1725=>x"d000", 1726=>x"c500", 1727=>x"ab00", 1728=>x"d800", 1729=>x"d800",
---- 1730=>x"d800", 1731=>x"d600", 1732=>x"d300", 1733=>x"cb00", 1734=>x"bb00", 1735=>x"9900", 1736=>x"da00",
---- 1737=>x"d900", 1738=>x"d900", 1739=>x"d600", 1740=>x"cf00", 1741=>x"c400", 1742=>x"ac00", 1743=>x"8600",
---- 1744=>x"da00", 1745=>x"d900", 1746=>x"d800", 1747=>x"d500", 1748=>x"ce00", 1749=>x"bb00", 1750=>x"9b00",
---- 1751=>x"7700", 1752=>x"d900", 1753=>x"d800", 1754=>x"d500", 1755=>x"d100", 1756=>x"c800", 1757=>x"ad00",
---- 1758=>x"8d00", 1759=>x"7200", 1760=>x"2600", 1761=>x"d800", 1762=>x"d700", 1763=>x"ce00", 1764=>x"bc00",
---- 1765=>x"9e00", 1766=>x"8300", 1767=>x"7200", 1768=>x"da00", 1769=>x"d700", 1770=>x"d200", 1771=>x"c800",
---- 1772=>x"ad00", 1773=>x"8d00", 1774=>x"7800", 1775=>x"7800", 1776=>x"d900", 1777=>x"d600", 1778=>x"cf00",
---- 1779=>x"bd00", 1780=>x"9d00", 1781=>x"8200", 1782=>x"7600", 1783=>x"7800", 1784=>x"2700", 1785=>x"d400",
---- 1786=>x"c900", 1787=>x"b300", 1788=>x"9000", 1789=>x"7900", 1790=>x"7100", 1791=>x"8900", 1792=>x"d700",
---- 1793=>x"d000", 1794=>x"c500", 1795=>x"a800", 1796=>x"8500", 1797=>x"7800", 1798=>x"7500", 1799=>x"7300",
---- 1800=>x"d600", 1801=>x"cd00", 1802=>x"bf00", 1803=>x"9f00", 1804=>x"7c00", 1805=>x"7500", 1806=>x"7500",
---- 1807=>x"7000", 1808=>x"d200", 1809=>x"cc00", 1810=>x"ba00", 1811=>x"9600", 1812=>x"7b00", 1813=>x"7100",
---- 1814=>x"6f00", 1815=>x"7000", 1816=>x"d100", 1817=>x"c900", 1818=>x"b400", 1819=>x"8f00", 1820=>x"7900",
---- 1821=>x"6e00", 1822=>x"6c00", 1823=>x"6a00", 1824=>x"d100", 1825=>x"c600", 1826=>x"ab00", 1827=>x"8700",
---- 1828=>x"7400", 1829=>x"7000", 1830=>x"6d00", 1831=>x"6400", 1832=>x"d000", 1833=>x"be00", 1834=>x"a000",
---- 1835=>x"8000", 1836=>x"7200", 1837=>x"6f00", 1838=>x"6a00", 1839=>x"6600", 1840=>x"cc00", 1841=>x"b400",
---- 1842=>x"9300", 1843=>x"7800", 1844=>x"7000", 1845=>x"6c00", 1846=>x"6400", 1847=>x"5e00", 1848=>x"c500",
---- 1849=>x"aa00", 1850=>x"8700", 1851=>x"7600", 1852=>x"6b00", 1853=>x"6200", 1854=>x"5700", 1855=>x"4f00",
---- 1856=>x"ba00", 1857=>x"9b00", 1858=>x"8000", 1859=>x"6e00", 1860=>x"5f00", 1861=>x"5900", 1862=>x"4f00",
---- 1863=>x"4b00", 1864=>x"a700", 1865=>x"8a00", 1866=>x"7500", 1867=>x"6200", 1868=>x"5500", 1869=>x"4e00",
---- 1870=>x"4a00", 1871=>x"4e00", 1872=>x"9800", 1873=>x"7d00", 1874=>x"6300", 1875=>x"5300", 1876=>x"4700",
---- 1877=>x"3e00", 1878=>x"4400", 1879=>x"5000", 1880=>x"8a00", 1881=>x"6b00", 1882=>x"5600", 1883=>x"4700",
---- 1884=>x"3a00", 1885=>x"3900", 1886=>x"4c00", 1887=>x"5100", 1888=>x"7700", 1889=>x"5700", 1890=>x"4b00",
---- 1891=>x"3e00", 1892=>x"3800", 1893=>x"4100", 1894=>x"4d00", 1895=>x"5200", 1896=>x"6100", 1897=>x"b800",
---- 1898=>x"3d00", 1899=>x"3b00", 1900=>x"4200", 1901=>x"4d00", 1902=>x"4f00", 1903=>x"5300", 1904=>x"4500",
---- 1905=>x"3d00", 1906=>x"ca00", 1907=>x"3f00", 1908=>x"4500", 1909=>x"4c00", 1910=>x"4f00", 1911=>x"4c00",
---- 1912=>x"3700", 1913=>x"3800", 1914=>x"3d00", 1915=>x"4200", 1916=>x"4b00", 1917=>x"4a00", 1918=>x"4400",
---- 1919=>x"4500", 1920=>x"3400", 1921=>x"3400", 1922=>x"3e00", 1923=>x"4600", 1924=>x"4c00", 1925=>x"4600",
---- 1926=>x"4100", 1927=>x"4a00", 1928=>x"3600", 1929=>x"3700", 1930=>x"4300", 1931=>x"4900", 1932=>x"4100",
---- 1933=>x"4000", 1934=>x"4900", 1935=>x"5600", 1936=>x"3d00", 1937=>x"4400", 1938=>x"4900", 1939=>x"4700",
---- 1940=>x"c000", 1941=>x"4500", 1942=>x"4f00", 1943=>x"5b00", 1944=>x"4400", 1945=>x"4c00", 1946=>x"4800",
---- 1947=>x"4200", 1948=>x"4600", 1949=>x"5100", 1950=>x"5b00", 1951=>x"6700", 1952=>x"4c00", 1953=>x"4b00",
---- 1954=>x"b800", 1955=>x"4700", 1956=>x"5100", 1957=>x"6000", 1958=>x"6b00", 1959=>x"6f00", 1960=>x"4e00",
---- 1961=>x"4900", 1962=>x"4700", 1963=>x"5000", 1964=>x"5c00", 1965=>x"6800", 1966=>x"7200", 1967=>x"6c00",
---- 1968=>x"4c00", 1969=>x"4600", 1970=>x"4f00", 1971=>x"5800", 1972=>x"6300", 1973=>x"6900", 1974=>x"6e00",
---- 1975=>x"6200", 1976=>x"4800", 1977=>x"4800", 1978=>x"5400", 1979=>x"5f00", 1980=>x"6800", 1981=>x"6900",
---- 1982=>x"6300", 1983=>x"5a00", 1984=>x"5000", 1985=>x"5100", 1986=>x"5900", 1987=>x"6700", 1988=>x"6900",
---- 1989=>x"6400", 1990=>x"5700", 1991=>x"5400", 1992=>x"5400", 1993=>x"5700", 1994=>x"6000", 1995=>x"6600",
---- 1996=>x"5900", 1997=>x"5400", 1998=>x"5000", 1999=>x"4700", 2000=>x"5b00", 2001=>x"6000", 2002=>x"6300",
---- 2003=>x"5e00", 2004=>x"5400", 2005=>x"4a00", 2006=>x"4500", 2007=>x"4300", 2008=>x"6100", 2009=>x"6200",
---- 2010=>x"6400", 2011=>x"5800", 2012=>x"4f00", 2013=>x"4700", 2014=>x"4500", 2015=>x"4800", 2016=>x"6400",
---- 2017=>x"5d00", 2018=>x"5a00", 2019=>x"5700", 2020=>x"5100", 2021=>x"5200", 2022=>x"4c00", 2023=>x"5000",
---- 2024=>x"5b00", 2025=>x"5600", 2026=>x"5000", 2027=>x"5100", 2028=>x"5600", 2029=>x"5500", 2030=>x"5200",
---- 2031=>x"4f00", 2032=>x"4f00", 2033=>x"4e00", 2034=>x"4d00", 2035=>x"5500", 2036=>x"5800", 2037=>x"5700",
---- 2038=>x"5400", 2039=>x"5300", 2040=>x"4a00", 2041=>x"4a00", 2042=>x"5400", 2043=>x"5c00", 2044=>x"5b00",
---- 2045=>x"5a00", 2046=>x"5600", 2047=>x"5300"),
---- 29 => (0=>x"7b00", 1=>x"7d00", 2=>x"7a00", 3=>x"7d00", 4=>x"7e00", 5=>x"7c00", 6=>x"7c00", 7=>x"7700",
---- 8=>x"7b00", 9=>x"7c00", 10=>x"7a00", 11=>x"7d00", 12=>x"7d00", 13=>x"7c00", 14=>x"7d00",
---- 15=>x"7700", 16=>x"7c00", 17=>x"7c00", 18=>x"7b00", 19=>x"7c00", 20=>x"7e00", 21=>x"7c00",
---- 22=>x"7e00", 23=>x"7600", 24=>x"7d00", 25=>x"7d00", 26=>x"7d00", 27=>x"7b00", 28=>x"7d00",
---- 29=>x"7a00", 30=>x"7c00", 31=>x"7900", 32=>x"7e00", 33=>x"7b00", 34=>x"7c00", 35=>x"7c00",
---- 36=>x"7a00", 37=>x"7a00", 38=>x"7b00", 39=>x"7d00", 40=>x"7900", 41=>x"7b00", 42=>x"7b00",
---- 43=>x"7900", 44=>x"7b00", 45=>x"7c00", 46=>x"7b00", 47=>x"7d00", 48=>x"7b00", 49=>x"7900",
---- 50=>x"7a00", 51=>x"7900", 52=>x"7b00", 53=>x"7b00", 54=>x"7b00", 55=>x"7900", 56=>x"7a00",
---- 57=>x"7700", 58=>x"7a00", 59=>x"7b00", 60=>x"7b00", 61=>x"7e00", 62=>x"7e00", 63=>x"7b00",
---- 64=>x"7a00", 65=>x"7b00", 66=>x"7c00", 67=>x"7c00", 68=>x"7a00", 69=>x"7d00", 70=>x"8100",
---- 71=>x"7d00", 72=>x"7a00", 73=>x"7e00", 74=>x"7b00", 75=>x"7c00", 76=>x"7d00", 77=>x"7c00",
---- 78=>x"8000", 79=>x"7e00", 80=>x"7800", 81=>x"7a00", 82=>x"7a00", 83=>x"8000", 84=>x"8000",
---- 85=>x"7f00", 86=>x"8000", 87=>x"8200", 88=>x"7a00", 89=>x"7900", 90=>x"7e00", 91=>x"8000",
---- 92=>x"8100", 93=>x"8300", 94=>x"8000", 95=>x"8300", 96=>x"7800", 97=>x"7800", 98=>x"7900",
---- 99=>x"7e00", 100=>x"7d00", 101=>x"7e00", 102=>x"8100", 103=>x"8400", 104=>x"8800", 105=>x"7b00",
---- 106=>x"7b00", 107=>x"7a00", 108=>x"7b00", 109=>x"7e00", 110=>x"8300", 111=>x"8500", 112=>x"7800",
---- 113=>x"7900", 114=>x"7b00", 115=>x"7d00", 116=>x"7e00", 117=>x"8100", 118=>x"8300", 119=>x"8a00",
---- 120=>x"7900", 121=>x"7b00", 122=>x"7a00", 123=>x"7e00", 124=>x"7f00", 125=>x"8300", 126=>x"8600",
---- 127=>x"8100", 128=>x"7d00", 129=>x"7c00", 130=>x"7c00", 131=>x"7f00", 132=>x"8100", 133=>x"8300",
---- 134=>x"8500", 135=>x"7300", 136=>x"7a00", 137=>x"7f00", 138=>x"7f00", 139=>x"8200", 140=>x"8700",
---- 141=>x"8400", 142=>x"7000", 143=>x"4900", 144=>x"7b00", 145=>x"8100", 146=>x"8400", 147=>x"8600",
---- 148=>x"8200", 149=>x"6d00", 150=>x"4a00", 151=>x"2a00", 152=>x"7e00", 153=>x"8100", 154=>x"7900",
---- 155=>x"8100", 156=>x"6c00", 157=>x"4700", 158=>x"2b00", 159=>x"2c00", 160=>x"7d00", 161=>x"8200",
---- 162=>x"8200", 163=>x"6e00", 164=>x"4a00", 165=>x"3000", 166=>x"2800", 167=>x"2e00", 168=>x"8200",
---- 169=>x"8100", 170=>x"6e00", 171=>x"4e00", 172=>x"2f00", 173=>x"2b00", 174=>x"2a00", 175=>x"2b00",
---- 176=>x"8100", 177=>x"6f00", 178=>x"4c00", 179=>x"3000", 180=>x"2c00", 181=>x"2a00", 182=>x"2d00",
---- 183=>x"2b00", 184=>x"6700", 185=>x"4a00", 186=>x"3200", 187=>x"2b00", 188=>x"2f00", 189=>x"3100",
---- 190=>x"2c00", 191=>x"2d00", 192=>x"4900", 193=>x"2a00", 194=>x"2b00", 195=>x"2b00", 196=>x"2b00",
---- 197=>x"2e00", 198=>x"2b00", 199=>x"3000", 200=>x"2e00", 201=>x"2800", 202=>x"2a00", 203=>x"2c00",
---- 204=>x"d300", 205=>x"2c00", 206=>x"2c00", 207=>x"2e00", 208=>x"2800", 209=>x"2700", 210=>x"2b00",
---- 211=>x"2a00", 212=>x"2d00", 213=>x"2e00", 214=>x"2c00", 215=>x"2e00", 216=>x"2c00", 217=>x"2a00",
---- 218=>x"2e00", 219=>x"3000", 220=>x"2f00", 221=>x"3200", 222=>x"3100", 223=>x"3600", 224=>x"2900",
---- 225=>x"2a00", 226=>x"3100", 227=>x"2d00", 228=>x"3400", 229=>x"3500", 230=>x"3600", 231=>x"3500",
---- 232=>x"2e00", 233=>x"2a00", 234=>x"2e00", 235=>x"2b00", 236=>x"3300", 237=>x"3700", 238=>x"3500",
---- 239=>x"3400", 240=>x"2d00", 241=>x"3000", 242=>x"3000", 243=>x"2d00", 244=>x"3200", 245=>x"3700",
---- 246=>x"3400", 247=>x"3100", 248=>x"2c00", 249=>x"2e00", 250=>x"2f00", 251=>x"3200", 252=>x"3600",
---- 253=>x"3700", 254=>x"3500", 255=>x"3600", 256=>x"2f00", 257=>x"2e00", 258=>x"3100", 259=>x"3500",
---- 260=>x"3700", 261=>x"3200", 262=>x"3400", 263=>x"3900", 264=>x"2e00", 265=>x"3100", 266=>x"3500",
---- 267=>x"3a00", 268=>x"3600", 269=>x"3700", 270=>x"3800", 271=>x"3800", 272=>x"2e00", 273=>x"3400",
---- 274=>x"3400", 275=>x"3300", 276=>x"3300", 277=>x"3700", 278=>x"3800", 279=>x"3400", 280=>x"3100",
---- 281=>x"3200", 282=>x"3100", 283=>x"3200", 284=>x"3600", 285=>x"cb00", 286=>x"3600", 287=>x"2f00",
---- 288=>x"3200", 289=>x"3100", 290=>x"cd00", 291=>x"3600", 292=>x"3500", 293=>x"3500", 294=>x"2f00",
---- 295=>x"d700", 296=>x"3b00", 297=>x"3600", 298=>x"cc00", 299=>x"3100", 300=>x"2e00", 301=>x"2d00",
---- 302=>x"2600", 303=>x"2a00", 304=>x"3500", 305=>x"3800", 306=>x"3600", 307=>x"3200", 308=>x"2c00",
---- 309=>x"2d00", 310=>x"2e00", 311=>x"3200", 312=>x"3500", 313=>x"3200", 314=>x"2c00", 315=>x"2c00",
---- 316=>x"2c00", 317=>x"2d00", 318=>x"3300", 319=>x"3900", 320=>x"3500", 321=>x"3300", 322=>x"3100",
---- 323=>x"2e00", 324=>x"2a00", 325=>x"3000", 326=>x"3700", 327=>x"3b00", 328=>x"3500", 329=>x"3200",
---- 330=>x"2d00", 331=>x"2c00", 332=>x"2b00", 333=>x"3700", 334=>x"3b00", 335=>x"3700", 336=>x"3000",
---- 337=>x"2d00", 338=>x"2a00", 339=>x"2f00", 340=>x"2f00", 341=>x"3600", 342=>x"3500", 343=>x"2e00",
---- 344=>x"2f00", 345=>x"2700", 346=>x"2c00", 347=>x"3400", 348=>x"3800", 349=>x"3700", 350=>x"2f00",
---- 351=>x"2d00", 352=>x"2d00", 353=>x"2a00", 354=>x"3500", 355=>x"3c00", 356=>x"3700", 357=>x"3000",
---- 358=>x"2b00", 359=>x"2c00", 360=>x"2d00", 361=>x"3000", 362=>x"3800", 363=>x"3a00", 364=>x"3300",
---- 365=>x"2e00", 366=>x"2e00", 367=>x"3100", 368=>x"2e00", 369=>x"3800", 370=>x"3c00", 371=>x"3300",
---- 372=>x"2f00", 373=>x"3100", 374=>x"3300", 375=>x"3400", 376=>x"3400", 377=>x"3a00", 378=>x"3e00",
---- 379=>x"2f00", 380=>x"2d00", 381=>x"3200", 382=>x"3400", 383=>x"3100", 384=>x"3900", 385=>x"3a00",
---- 386=>x"2e00", 387=>x"2b00", 388=>x"3300", 389=>x"3400", 390=>x"3500", 391=>x"3600", 392=>x"3c00",
---- 393=>x"3200", 394=>x"2d00", 395=>x"2d00", 396=>x"3600", 397=>x"3500", 398=>x"3600", 399=>x"3700",
---- 400=>x"3500", 401=>x"2c00", 402=>x"3100", 403=>x"2f00", 404=>x"3400", 405=>x"3700", 406=>x"3600",
---- 407=>x"3600", 408=>x"3000", 409=>x"2c00", 410=>x"3700", 411=>x"3400", 412=>x"3300", 413=>x"3400",
---- 414=>x"3700", 415=>x"3400", 416=>x"d600", 417=>x"d300", 418=>x"3300", 419=>x"3500", 420=>x"3b00",
---- 421=>x"3400", 422=>x"3200", 423=>x"3300", 424=>x"2e00", 425=>x"3300", 426=>x"3600", 427=>x"3100",
---- 428=>x"3500", 429=>x"3000", 430=>x"3100", 431=>x"3700", 432=>x"3400", 433=>x"3700", 434=>x"3b00",
---- 435=>x"3500", 436=>x"3000", 437=>x"2a00", 438=>x"3000", 439=>x"4600", 440=>x"3500", 441=>x"3b00",
---- 442=>x"3500", 443=>x"3000", 444=>x"2800", 445=>x"2600", 446=>x"3600", 447=>x"5b00", 448=>x"3800",
---- 449=>x"3500", 450=>x"3200", 451=>x"2f00", 452=>x"2700", 453=>x"2c00", 454=>x"4f00", 455=>x"7a00",
---- 456=>x"3700", 457=>x"2f00", 458=>x"2900", 459=>x"2d00", 460=>x"3300", 461=>x"4a00", 462=>x"7100",
---- 463=>x"8c00", 464=>x"3500", 465=>x"2900", 466=>x"d800", 467=>x"2b00", 468=>x"c000", 469=>x"6a00",
---- 470=>x"8700", 471=>x"9500", 472=>x"3700", 473=>x"2d00", 474=>x"2900", 475=>x"3000", 476=>x"5700",
---- 477=>x"8000", 478=>x"9500", 479=>x"9700", 480=>x"3200", 481=>x"2c00", 482=>x"3200", 483=>x"4c00",
---- 484=>x"7600", 485=>x"9100", 486=>x"9900", 487=>x"9600", 488=>x"2f00", 489=>x"3100", 490=>x"4100",
---- 491=>x"6b00", 492=>x"8b00", 493=>x"9600", 494=>x"9800", 495=>x"9100", 496=>x"3100", 497=>x"3700",
---- 498=>x"5a00", 499=>x"8300", 500=>x"9500", 501=>x"9a00", 502=>x"9300", 503=>x"7100", 504=>x"2f00",
---- 505=>x"4700", 506=>x"7500", 507=>x"9300", 508=>x"9c00", 509=>x"9600", 510=>x"9100", 511=>x"8e00",
---- 512=>x"3800", 513=>x"6400", 514=>x"8d00", 515=>x"9b00", 516=>x"9a00", 517=>x"9400", 518=>x"8f00",
---- 519=>x"9100", 520=>x"4c00", 521=>x"8100", 522=>x"9a00", 523=>x"9b00", 524=>x"9400", 525=>x"9100",
---- 526=>x"8e00", 527=>x"9900", 528=>x"6e00", 529=>x"9200", 530=>x"9a00", 531=>x"9600", 532=>x"9200",
---- 533=>x"8f00", 534=>x"9300", 535=>x"9d00", 536=>x"8700", 537=>x"9900", 538=>x"9b00", 539=>x"9600",
---- 540=>x"8e00", 541=>x"9200", 542=>x"9a00", 543=>x"a000", 544=>x"9200", 545=>x"9c00", 546=>x"9900",
---- 547=>x"9400", 548=>x"9000", 549=>x"9600", 550=>x"9f00", 551=>x"a300", 552=>x"9800", 553=>x"9a00",
---- 554=>x"9600", 555=>x"9000", 556=>x"9300", 557=>x"9c00", 558=>x"9f00", 559=>x"a200", 560=>x"6400",
---- 561=>x"9500", 562=>x"9300", 563=>x"9200", 564=>x"9600", 565=>x"9e00", 566=>x"a100", 567=>x"a100",
---- 568=>x"9500", 569=>x"9200", 570=>x"9100", 571=>x"9500", 572=>x"9d00", 573=>x"a000", 574=>x"a000",
---- 575=>x"a000", 576=>x"9400", 577=>x"8f00", 578=>x"9300", 579=>x"9800", 580=>x"9f00", 581=>x"a200",
---- 582=>x"a000", 583=>x"9f00", 584=>x"9100", 585=>x"9200", 586=>x"9700", 587=>x"9c00", 588=>x"9f00",
---- 589=>x"a100", 590=>x"a100", 591=>x"a000", 592=>x"9000", 593=>x"9400", 594=>x"9b00", 595=>x"9f00",
---- 596=>x"a100", 597=>x"a200", 598=>x"a200", 599=>x"a000", 600=>x"8f00", 601=>x"9500", 602=>x"9f00",
---- 603=>x"a000", 604=>x"a100", 605=>x"a000", 606=>x"9f00", 607=>x"a100", 608=>x"9600", 609=>x"9c00",
---- 610=>x"a000", 611=>x"a000", 612=>x"a100", 613=>x"a200", 614=>x"a000", 615=>x"a100", 616=>x"9c00",
---- 617=>x"a000", 618=>x"a000", 619=>x"a000", 620=>x"a300", 621=>x"a200", 622=>x"a100", 623=>x"9f00",
---- 624=>x"9c00", 625=>x"9f00", 626=>x"a000", 627=>x"a200", 628=>x"a300", 629=>x"a000", 630=>x"a000",
---- 631=>x"a000", 632=>x"9e00", 633=>x"9f00", 634=>x"a200", 635=>x"a000", 636=>x"a100", 637=>x"9c00",
---- 638=>x"9e00", 639=>x"a100", 640=>x"a000", 641=>x"a100", 642=>x"a100", 643=>x"a100", 644=>x"a000",
---- 645=>x"9e00", 646=>x"a000", 647=>x"9f00", 648=>x"9f00", 649=>x"a200", 650=>x"a000", 651=>x"a200",
---- 652=>x"a300", 653=>x"9e00", 654=>x"9e00", 655=>x"9e00", 656=>x"a000", 657=>x"a100", 658=>x"a000",
---- 659=>x"9e00", 660=>x"9e00", 661=>x"6300", 662=>x"6400", 663=>x"9b00", 664=>x"a100", 665=>x"a000",
---- 666=>x"9e00", 667=>x"9d00", 668=>x"9c00", 669=>x"9b00", 670=>x"9e00", 671=>x"9d00", 672=>x"9f00",
---- 673=>x"9f00", 674=>x"9d00", 675=>x"9d00", 676=>x"9d00", 677=>x"9c00", 678=>x"9c00", 679=>x"9d00",
---- 680=>x"9f00", 681=>x"9e00", 682=>x"9e00", 683=>x"9e00", 684=>x"9b00", 685=>x"9c00", 686=>x"9c00",
---- 687=>x"9b00", 688=>x"a000", 689=>x"9e00", 690=>x"a000", 691=>x"9c00", 692=>x"9c00", 693=>x"9b00",
---- 694=>x"9c00", 695=>x"9c00", 696=>x"9e00", 697=>x"9f00", 698=>x"9e00", 699=>x"9c00", 700=>x"9e00",
---- 701=>x"9d00", 702=>x"9e00", 703=>x"9c00", 704=>x"9f00", 705=>x"9f00", 706=>x"9f00", 707=>x"9f00",
---- 708=>x"9c00", 709=>x"9b00", 710=>x"9d00", 711=>x"9e00", 712=>x"9f00", 713=>x"9e00", 714=>x"9f00",
---- 715=>x"9e00", 716=>x"9d00", 717=>x"9a00", 718=>x"9b00", 719=>x"9c00", 720=>x"9f00", 721=>x"9f00",
---- 722=>x"a000", 723=>x"9d00", 724=>x"a000", 725=>x"9e00", 726=>x"9d00", 727=>x"9c00", 728=>x"9f00",
---- 729=>x"a000", 730=>x"a200", 731=>x"9f00", 732=>x"9d00", 733=>x"9f00", 734=>x"9e00", 735=>x"9d00",
---- 736=>x"a200", 737=>x"9f00", 738=>x"a000", 739=>x"9f00", 740=>x"9e00", 741=>x"9e00", 742=>x"6100",
---- 743=>x"9b00", 744=>x"a000", 745=>x"a000", 746=>x"9f00", 747=>x"9f00", 748=>x"9e00", 749=>x"9e00",
---- 750=>x"9d00", 751=>x"9d00", 752=>x"a200", 753=>x"a000", 754=>x"a100", 755=>x"9e00", 756=>x"9f00",
---- 757=>x"9f00", 758=>x"9d00", 759=>x"9e00", 760=>x"a100", 761=>x"9f00", 762=>x"9f00", 763=>x"9e00",
---- 764=>x"a000", 765=>x"a000", 766=>x"9e00", 767=>x"9e00", 768=>x"a400", 769=>x"a300", 770=>x"a100",
---- 771=>x"a000", 772=>x"9f00", 773=>x"9f00", 774=>x"9c00", 775=>x"9f00", 776=>x"a200", 777=>x"a100",
---- 778=>x"a100", 779=>x"a000", 780=>x"9f00", 781=>x"9f00", 782=>x"9e00", 783=>x"a000", 784=>x"a200",
---- 785=>x"a100", 786=>x"a200", 787=>x"9f00", 788=>x"9d00", 789=>x"6100", 790=>x"9d00", 791=>x"9f00",
---- 792=>x"a200", 793=>x"a300", 794=>x"a200", 795=>x"a000", 796=>x"9f00", 797=>x"9f00", 798=>x"a000",
---- 799=>x"6000", 800=>x"a200", 801=>x"5c00", 802=>x"a200", 803=>x"a100", 804=>x"a000", 805=>x"a100",
---- 806=>x"9c00", 807=>x"9e00", 808=>x"a400", 809=>x"a300", 810=>x"a200", 811=>x"a200", 812=>x"a100",
---- 813=>x"a100", 814=>x"9d00", 815=>x"9f00", 816=>x"a200", 817=>x"a200", 818=>x"a300", 819=>x"a200",
---- 820=>x"a100", 821=>x"a000", 822=>x"a100", 823=>x"a100", 824=>x"a500", 825=>x"a400", 826=>x"a300",
---- 827=>x"5e00", 828=>x"a200", 829=>x"9f00", 830=>x"a100", 831=>x"a000", 832=>x"a400", 833=>x"a100",
---- 834=>x"a100", 835=>x"a200", 836=>x"a200", 837=>x"9f00", 838=>x"9f00", 839=>x"9f00", 840=>x"a100",
---- 841=>x"a100", 842=>x"9f00", 843=>x"a300", 844=>x"a100", 845=>x"a200", 846=>x"a200", 847=>x"9f00",
---- 848=>x"a400", 849=>x"a200", 850=>x"a100", 851=>x"a400", 852=>x"a300", 853=>x"a200", 854=>x"a100",
---- 855=>x"a100", 856=>x"a400", 857=>x"a500", 858=>x"a300", 859=>x"a000", 860=>x"a200", 861=>x"a300",
---- 862=>x"9e00", 863=>x"a000", 864=>x"a300", 865=>x"a200", 866=>x"a300", 867=>x"a400", 868=>x"a200",
---- 869=>x"a200", 870=>x"a100", 871=>x"a200", 872=>x"a400", 873=>x"a100", 874=>x"a300", 875=>x"a400",
---- 876=>x"a200", 877=>x"a300", 878=>x"a200", 879=>x"a200", 880=>x"a100", 881=>x"a200", 882=>x"a000",
---- 883=>x"a300", 884=>x"a400", 885=>x"a400", 886=>x"a100", 887=>x"a100", 888=>x"a000", 889=>x"a100",
---- 890=>x"a100", 891=>x"a200", 892=>x"a100", 893=>x"a400", 894=>x"a400", 895=>x"a100", 896=>x"a100",
---- 897=>x"a100", 898=>x"a000", 899=>x"a200", 900=>x"a300", 901=>x"a300", 902=>x"a500", 903=>x"a100",
---- 904=>x"a100", 905=>x"a000", 906=>x"a200", 907=>x"5e00", 908=>x"a000", 909=>x"a000", 910=>x"a100",
---- 911=>x"a200", 912=>x"9a00", 913=>x"9a00", 914=>x"9d00", 915=>x"9f00", 916=>x"9f00", 917=>x"a200",
---- 918=>x"a400", 919=>x"a000", 920=>x"9400", 921=>x"9200", 922=>x"9600", 923=>x"9800", 924=>x"9a00",
---- 925=>x"9e00", 926=>x"a100", 927=>x"a100", 928=>x"9200", 929=>x"9200", 930=>x"9300", 931=>x"9200",
---- 932=>x"9000", 933=>x"6900", 934=>x"9a00", 935=>x"9b00", 936=>x"9400", 937=>x"9100", 938=>x"9200",
---- 939=>x"9100", 940=>x"9100", 941=>x"9100", 942=>x"9300", 943=>x"9000", 944=>x"9900", 945=>x"9200",
---- 946=>x"9100", 947=>x"9000", 948=>x"9300", 949=>x"9500", 950=>x"9200", 951=>x"9100", 952=>x"9900",
---- 953=>x"9500", 954=>x"9300", 955=>x"9100", 956=>x"9200", 957=>x"9600", 958=>x"9200", 959=>x"9100",
---- 960=>x"9a00", 961=>x"9700", 962=>x"9400", 963=>x"9400", 964=>x"9500", 965=>x"9400", 966=>x"9200",
---- 967=>x"9000", 968=>x"9c00", 969=>x"9d00", 970=>x"9800", 971=>x"9700", 972=>x"9500", 973=>x"9300",
---- 974=>x"9400", 975=>x"9000", 976=>x"9d00", 977=>x"9e00", 978=>x"9b00", 979=>x"9d00", 980=>x"9900",
---- 981=>x"9700", 982=>x"9600", 983=>x"9300", 984=>x"9900", 985=>x"9900", 986=>x"9b00", 987=>x"9d00",
---- 988=>x"9c00", 989=>x"9a00", 990=>x"9900", 991=>x"9800", 992=>x"9800", 993=>x"9a00", 994=>x"9c00",
---- 995=>x"9b00", 996=>x"9b00", 997=>x"9a00", 998=>x"9a00", 999=>x"9b00", 1000=>x"9b00", 1001=>x"9b00",
---- 1002=>x"9a00", 1003=>x"9a00", 1004=>x"9c00", 1005=>x"9a00", 1006=>x"9a00", 1007=>x"9a00", 1008=>x"9c00",
---- 1009=>x"9a00", 1010=>x"9900", 1011=>x"9700", 1012=>x"9b00", 1013=>x"9a00", 1014=>x"9c00", 1015=>x"9d00",
---- 1016=>x"9a00", 1017=>x"9c00", 1018=>x"9a00", 1019=>x"9900", 1020=>x"9900", 1021=>x"9b00", 1022=>x"9900",
---- 1023=>x"9a00", 1024=>x"9a00", 1025=>x"9900", 1026=>x"9800", 1027=>x"9800", 1028=>x"9a00", 1029=>x"9a00",
---- 1030=>x"9900", 1031=>x"9a00", 1032=>x"9900", 1033=>x"9800", 1034=>x"9a00", 1035=>x"9800", 1036=>x"9c00",
---- 1037=>x"9a00", 1038=>x"9800", 1039=>x"9900", 1040=>x"9a00", 1041=>x"9900", 1042=>x"9900", 1043=>x"9900",
---- 1044=>x"9900", 1045=>x"9800", 1046=>x"9800", 1047=>x"9800", 1048=>x"9900", 1049=>x"9700", 1050=>x"9b00",
---- 1051=>x"9c00", 1052=>x"9900", 1053=>x"6700", 1054=>x"9800", 1055=>x"9500", 1056=>x"9900", 1057=>x"9800",
---- 1058=>x"9900", 1059=>x"9a00", 1060=>x"9a00", 1061=>x"9800", 1062=>x"9800", 1063=>x"9500", 1064=>x"9900",
---- 1065=>x"9800", 1066=>x"9700", 1067=>x"9800", 1068=>x"9700", 1069=>x"9500", 1070=>x"9200", 1071=>x"9200",
---- 1072=>x"9800", 1073=>x"9700", 1074=>x"9600", 1075=>x"9400", 1076=>x"9400", 1077=>x"9700", 1078=>x"9400",
---- 1079=>x"9000", 1080=>x"9600", 1081=>x"9700", 1082=>x"9600", 1083=>x"9100", 1084=>x"9200", 1085=>x"9500",
---- 1086=>x"9100", 1087=>x"9500", 1088=>x"9600", 1089=>x"9800", 1090=>x"9700", 1091=>x"9200", 1092=>x"9500",
---- 1093=>x"9300", 1094=>x"9000", 1095=>x"8f00", 1096=>x"9600", 1097=>x"9300", 1098=>x"9400", 1099=>x"9200",
---- 1100=>x"9100", 1101=>x"9200", 1102=>x"8f00", 1103=>x"8e00", 1104=>x"9200", 1105=>x"9300", 1106=>x"9400",
---- 1107=>x"8e00", 1108=>x"8b00", 1109=>x"8f00", 1110=>x"8e00", 1111=>x"8b00", 1112=>x"9000", 1113=>x"8e00",
---- 1114=>x"9100", 1115=>x"8d00", 1116=>x"8b00", 1117=>x"8b00", 1118=>x"8800", 1119=>x"8700", 1120=>x"9100",
---- 1121=>x"9200", 1122=>x"9000", 1123=>x"8b00", 1124=>x"8d00", 1125=>x"8a00", 1126=>x"8600", 1127=>x"8800",
---- 1128=>x"9000", 1129=>x"8e00", 1130=>x"8f00", 1131=>x"8d00", 1132=>x"8c00", 1133=>x"8900", 1134=>x"8900",
---- 1135=>x"8500", 1136=>x"8e00", 1137=>x"8e00", 1138=>x"8c00", 1139=>x"8d00", 1140=>x"8900", 1141=>x"8500",
---- 1142=>x"8300", 1143=>x"8100", 1144=>x"8f00", 1145=>x"8e00", 1146=>x"8f00", 1147=>x"8a00", 1148=>x"8600",
---- 1149=>x"8300", 1150=>x"8100", 1151=>x"9000", 1152=>x"8c00", 1153=>x"8c00", 1154=>x"8900", 1155=>x"8600",
---- 1156=>x"8500", 1157=>x"8200", 1158=>x"9000", 1159=>x"a500", 1160=>x"8b00", 1161=>x"8900", 1162=>x"8700",
---- 1163=>x"8700", 1164=>x"8300", 1165=>x"8e00", 1166=>x"a400", 1167=>x"b400", 1168=>x"8900", 1169=>x"8600",
---- 1170=>x"8600", 1171=>x"8400", 1172=>x"8b00", 1173=>x"a200", 1174=>x"4c00", 1175=>x"bd00", 1176=>x"8700",
---- 1177=>x"8400", 1178=>x"8300", 1179=>x"8600", 1180=>x"9a00", 1181=>x"b000", 1182=>x"ba00", 1183=>x"c000",
---- 1184=>x"8600", 1185=>x"8200", 1186=>x"8300", 1187=>x"9300", 1188=>x"ab00", 1189=>x"b800", 1190=>x"c000",
---- 1191=>x"c300", 1192=>x"8400", 1193=>x"7d00", 1194=>x"8a00", 1195=>x"a200", 1196=>x"b700", 1197=>x"bf00",
---- 1198=>x"c400", 1199=>x"c400", 1200=>x"8200", 1201=>x"8000", 1202=>x"9800", 1203=>x"af00", 1204=>x"bc00",
---- 1205=>x"c200", 1206=>x"c400", 1207=>x"c400", 1208=>x"8100", 1209=>x"9000", 1210=>x"a800", 1211=>x"bb00",
---- 1212=>x"c100", 1213=>x"c400", 1214=>x"c400", 1215=>x"c100", 1216=>x"8600", 1217=>x"9d00", 1218=>x"b300",
---- 1219=>x"be00", 1220=>x"c300", 1221=>x"c200", 1222=>x"c300", 1223=>x"c000", 1224=>x"9200", 1225=>x"ac00",
---- 1226=>x"bb00", 1227=>x"c200", 1228=>x"c500", 1229=>x"c300", 1230=>x"c300", 1231=>x"c000", 1232=>x"a000",
---- 1233=>x"b700", 1234=>x"bf00", 1235=>x"c300", 1236=>x"c400", 1237=>x"3c00", 1238=>x"c000", 1239=>x"c000",
---- 1240=>x"ad00", 1241=>x"bc00", 1242=>x"c300", 1243=>x"c400", 1244=>x"c300", 1245=>x"c200", 1246=>x"c100",
---- 1247=>x"c200", 1248=>x"b600", 1249=>x"c000", 1250=>x"c500", 1251=>x"c400", 1252=>x"c200", 1253=>x"c200",
---- 1254=>x"c100", 1255=>x"c300", 1256=>x"be00", 1257=>x"c500", 1258=>x"c500", 1259=>x"c300", 1260=>x"c300",
---- 1261=>x"c100", 1262=>x"c200", 1263=>x"c200", 1264=>x"c200", 1265=>x"c600", 1266=>x"c300", 1267=>x"c300",
---- 1268=>x"c200", 1269=>x"c300", 1270=>x"c200", 1271=>x"c400", 1272=>x"c400", 1273=>x"c600", 1274=>x"c400",
---- 1275=>x"c300", 1276=>x"c200", 1277=>x"c200", 1278=>x"c000", 1279=>x"c500", 1280=>x"c700", 1281=>x"c300",
---- 1282=>x"c200", 1283=>x"c200", 1284=>x"c200", 1285=>x"c200", 1286=>x"c500", 1287=>x"ca00", 1288=>x"c500",
---- 1289=>x"3a00", 1290=>x"c100", 1291=>x"c200", 1292=>x"c200", 1293=>x"c500", 1294=>x"c800", 1295=>x"cc00",
---- 1296=>x"c500", 1297=>x"c300", 1298=>x"c500", 1299=>x"c400", 1300=>x"c500", 1301=>x"c700", 1302=>x"cb00",
---- 1303=>x"ce00", 1304=>x"c400", 1305=>x"c400", 1306=>x"c400", 1307=>x"c300", 1308=>x"c700", 1309=>x"c900",
---- 1310=>x"ce00", 1311=>x"cf00", 1312=>x"c400", 1313=>x"c500", 1314=>x"c400", 1315=>x"c500", 1316=>x"ca00",
---- 1317=>x"cc00", 1318=>x"d000", 1319=>x"d100", 1320=>x"c400", 1321=>x"c400", 1322=>x"c500", 1323=>x"c800",
---- 1324=>x"cc00", 1325=>x"cc00", 1326=>x"cf00", 1327=>x"d000", 1328=>x"c300", 1329=>x"c400", 1330=>x"3a00",
---- 1331=>x"c900", 1332=>x"cd00", 1333=>x"d000", 1334=>x"d100", 1335=>x"d000", 1336=>x"c300", 1337=>x"c500",
---- 1338=>x"c700", 1339=>x"cc00", 1340=>x"cf00", 1341=>x"d100", 1342=>x"d100", 1343=>x"d000", 1344=>x"c400",
---- 1345=>x"c700", 1346=>x"ca00", 1347=>x"ce00", 1348=>x"d100", 1349=>x"d200", 1350=>x"d100", 1351=>x"cf00",
---- 1352=>x"c500", 1353=>x"c900", 1354=>x"cc00", 1355=>x"d100", 1356=>x"d100", 1357=>x"d100", 1358=>x"d100",
---- 1359=>x"ce00", 1360=>x"c600", 1361=>x"cc00", 1362=>x"ce00", 1363=>x"2e00", 1364=>x"d100", 1365=>x"d100",
---- 1366=>x"d000", 1367=>x"cf00", 1368=>x"cb00", 1369=>x"ce00", 1370=>x"d100", 1371=>x"cf00", 1372=>x"d100",
---- 1373=>x"d000", 1374=>x"d000", 1375=>x"cf00", 1376=>x"cc00", 1377=>x"cf00", 1378=>x"d300", 1379=>x"d300",
---- 1380=>x"d100", 1381=>x"cf00", 1382=>x"cf00", 1383=>x"d000", 1384=>x"cd00", 1385=>x"d100", 1386=>x"d300",
---- 1387=>x"d100", 1388=>x"d100", 1389=>x"d100", 1390=>x"d000", 1391=>x"d100", 1392=>x"cf00", 1393=>x"d400",
---- 1394=>x"d100", 1395=>x"d200", 1396=>x"d100", 1397=>x"d100", 1398=>x"d300", 1399=>x"d100", 1400=>x"d300",
---- 1401=>x"d400", 1402=>x"d400", 1403=>x"d200", 1404=>x"d200", 1405=>x"d300", 1406=>x"d100", 1407=>x"d100",
---- 1408=>x"d500", 1409=>x"d400", 1410=>x"d300", 1411=>x"d300", 1412=>x"d300", 1413=>x"d100", 1414=>x"d100",
---- 1415=>x"d100", 1416=>x"d400", 1417=>x"d400", 1418=>x"d200", 1419=>x"d200", 1420=>x"d300", 1421=>x"d200",
---- 1422=>x"d300", 1423=>x"d100", 1424=>x"d400", 1425=>x"d400", 1426=>x"d300", 1427=>x"d200", 1428=>x"d200",
---- 1429=>x"d300", 1430=>x"2c00", 1431=>x"d100", 1432=>x"2b00", 1433=>x"d300", 1434=>x"d500", 1435=>x"d200",
---- 1436=>x"d300", 1437=>x"d300", 1438=>x"d300", 1439=>x"d500", 1440=>x"d600", 1441=>x"d500", 1442=>x"d500",
---- 1443=>x"d300", 1444=>x"d200", 1445=>x"d500", 1446=>x"d600", 1447=>x"d600", 1448=>x"d500", 1449=>x"d300",
---- 1450=>x"d500", 1451=>x"d400", 1452=>x"d600", 1453=>x"d400", 1454=>x"d600", 1455=>x"d800", 1456=>x"d600",
---- 1457=>x"2a00", 1458=>x"d600", 1459=>x"d500", 1460=>x"d400", 1461=>x"d600", 1462=>x"d700", 1463=>x"d900",
---- 1464=>x"d500", 1465=>x"d700", 1466=>x"d700", 1467=>x"d500", 1468=>x"d600", 1469=>x"d700", 1470=>x"d800",
---- 1471=>x"d900", 1472=>x"d700", 1473=>x"d400", 1474=>x"d800", 1475=>x"d700", 1476=>x"d800", 1477=>x"d700",
---- 1478=>x"d700", 1479=>x"d900", 1480=>x"d700", 1481=>x"d700", 1482=>x"d700", 1483=>x"d900", 1484=>x"d800",
---- 1485=>x"d600", 1486=>x"d600", 1487=>x"d700", 1488=>x"d900", 1489=>x"d600", 1490=>x"d600", 1491=>x"d600",
---- 1492=>x"d600", 1493=>x"d500", 1494=>x"d500", 1495=>x"d400", 1496=>x"d900", 1497=>x"d500", 1498=>x"d500",
---- 1499=>x"d400", 1500=>x"d400", 1501=>x"d400", 1502=>x"2c00", 1503=>x"d500", 1504=>x"d600", 1505=>x"d400",
---- 1506=>x"d400", 1507=>x"d200", 1508=>x"d500", 1509=>x"d400", 1510=>x"d500", 1511=>x"d800", 1512=>x"d500",
---- 1513=>x"d300", 1514=>x"d300", 1515=>x"d300", 1516=>x"d500", 1517=>x"d600", 1518=>x"d600", 1519=>x"d700",
---- 1520=>x"d400", 1521=>x"d200", 1522=>x"d400", 1523=>x"d400", 1524=>x"d600", 1525=>x"d700", 1526=>x"d600",
---- 1527=>x"d800", 1528=>x"d300", 1529=>x"d200", 1530=>x"d500", 1531=>x"d500", 1532=>x"d400", 1533=>x"d600",
---- 1534=>x"d600", 1535=>x"d600", 1536=>x"d300", 1537=>x"d400", 1538=>x"d500", 1539=>x"d400", 1540=>x"d500",
---- 1541=>x"d500", 1542=>x"d500", 1543=>x"d300", 1544=>x"d300", 1545=>x"d400", 1546=>x"d200", 1547=>x"d300",
---- 1548=>x"d300", 1549=>x"d400", 1550=>x"d200", 1551=>x"d200", 1552=>x"d200", 1553=>x"d200", 1554=>x"d200",
---- 1555=>x"d200", 1556=>x"d200", 1557=>x"d200", 1558=>x"d100", 1559=>x"d000", 1560=>x"d200", 1561=>x"d000",
---- 1562=>x"2a00", 1563=>x"d100", 1564=>x"d000", 1565=>x"d000", 1566=>x"cf00", 1567=>x"ce00", 1568=>x"3000",
---- 1569=>x"d200", 1570=>x"d200", 1571=>x"d000", 1572=>x"d100", 1573=>x"d100", 1574=>x"cd00", 1575=>x"cc00",
---- 1576=>x"cf00", 1577=>x"d100", 1578=>x"d100", 1579=>x"d000", 1580=>x"d100", 1581=>x"d100", 1582=>x"cb00",
---- 1583=>x"c700", 1584=>x"d000", 1585=>x"d100", 1586=>x"d200", 1587=>x"d000", 1588=>x"d000", 1589=>x"d200",
---- 1590=>x"cc00", 1591=>x"c200", 1592=>x"cf00", 1593=>x"cf00", 1594=>x"d100", 1595=>x"d000", 1596=>x"d000",
---- 1597=>x"d100", 1598=>x"cb00", 1599=>x"bf00", 1600=>x"d100", 1601=>x"d000", 1602=>x"d000", 1603=>x"cf00",
---- 1604=>x"ce00", 1605=>x"ca00", 1606=>x"c400", 1607=>x"b600", 1608=>x"d200", 1609=>x"cf00", 1610=>x"cf00",
---- 1611=>x"ce00", 1612=>x"c800", 1613=>x"bd00", 1614=>x"b300", 1615=>x"9a00", 1616=>x"d300", 1617=>x"d100",
---- 1618=>x"d000", 1619=>x"ce00", 1620=>x"c100", 1621=>x"a800", 1622=>x"8a00", 1623=>x"5b00", 1624=>x"d300",
---- 1625=>x"d100", 1626=>x"cf00", 1627=>x"cd00", 1628=>x"b900", 1629=>x"8b00", 1630=>x"5400", 1631=>x"3300",
---- 1632=>x"d300", 1633=>x"ce00", 1634=>x"cc00", 1635=>x"c500", 1636=>x"a900", 1637=>x"7300", 1638=>x"3700",
---- 1639=>x"2a00", 1640=>x"d100", 1641=>x"cb00", 1642=>x"c500", 1643=>x"ba00", 1644=>x"9800", 1645=>x"5a00",
---- 1646=>x"2c00", 1647=>x"2b00", 1648=>x"d100", 1649=>x"c900", 1650=>x"bd00", 1651=>x"a900", 1652=>x"8500",
---- 1653=>x"4900", 1654=>x"3000", 1655=>x"3a00", 1656=>x"d000", 1657=>x"c500", 1658=>x"b400", 1659=>x"9700",
---- 1660=>x"7000", 1661=>x"4200", 1662=>x"3a00", 1663=>x"4e00", 1664=>x"ce00", 1665=>x"c100", 1666=>x"a500",
---- 1667=>x"8500", 1668=>x"5a00", 1669=>x"4200", 1670=>x"4800", 1671=>x"5900", 1672=>x"cb00", 1673=>x"bc00",
---- 1674=>x"9700", 1675=>x"6b00", 1676=>x"4c00", 1677=>x"4700", 1678=>x"5200", 1679=>x"6100", 1680=>x"c700",
---- 1681=>x"b300", 1682=>x"8300", 1683=>x"5400", 1684=>x"4b00", 1685=>x"5200", 1686=>x"5700", 1687=>x"5f00",
---- 1688=>x"c700", 1689=>x"a400", 1690=>x"6f00", 1691=>x"4c00", 1692=>x"4f00", 1693=>x"5700", 1694=>x"5d00",
---- 1695=>x"5a00", 1696=>x"ba00", 1697=>x"9100", 1698=>x"6100", 1699=>x"5100", 1700=>x"5800", 1701=>x"a200",
---- 1702=>x"5e00", 1703=>x"5800", 1704=>x"ac00", 1705=>x"7c00", 1706=>x"5700", 1707=>x"5a00", 1708=>x"5b00",
---- 1709=>x"6200", 1710=>x"5e00", 1711=>x"5b00", 1712=>x"9600", 1713=>x"6500", 1714=>x"5900", 1715=>x"5b00",
---- 1716=>x"5d00", 1717=>x"5f00", 1718=>x"5b00", 1719=>x"6200", 1720=>x"8200", 1721=>x"5e00", 1722=>x"5900",
---- 1723=>x"5d00", 1724=>x"5c00", 1725=>x"5b00", 1726=>x"5e00", 1727=>x"6800", 1728=>x"7200", 1729=>x"5b00",
---- 1730=>x"5b00", 1731=>x"5f00", 1732=>x"5c00", 1733=>x"5b00", 1734=>x"6300", 1735=>x"6600", 1736=>x"6700",
---- 1737=>x"5e00", 1738=>x"5e00", 1739=>x"5b00", 1740=>x"5a00", 1741=>x"5d00", 1742=>x"6200", 1743=>x"6800",
---- 1744=>x"6200", 1745=>x"6200", 1746=>x"5e00", 1747=>x"5900", 1748=>x"5700", 1749=>x"5e00", 1750=>x"6100",
---- 1751=>x"6b00", 1752=>x"6900", 1753=>x"6600", 1754=>x"6400", 1755=>x"5e00", 1756=>x"5e00", 1757=>x"5e00",
---- 1758=>x"6400", 1759=>x"6e00", 1760=>x"6b00", 1761=>x"6900", 1762=>x"6700", 1763=>x"6200", 1764=>x"6200",
---- 1765=>x"6100", 1766=>x"6500", 1767=>x"7100", 1768=>x"7100", 1769=>x"6700", 1770=>x"6000", 1771=>x"5f00",
---- 1772=>x"6200", 1773=>x"6500", 1774=>x"6500", 1775=>x"6c00", 1776=>x"7100", 1777=>x"6900", 1778=>x"6400",
---- 1779=>x"6200", 1780=>x"6100", 1781=>x"9b00", 1782=>x"6a00", 1783=>x"6d00", 1784=>x"7000", 1785=>x"6700",
---- 1786=>x"6900", 1787=>x"6000", 1788=>x"6000", 1789=>x"6700", 1790=>x"6a00", 1791=>x"6c00", 1792=>x"7100",
---- 1793=>x"6a00", 1794=>x"6600", 1795=>x"5d00", 1796=>x"5c00", 1797=>x"6500", 1798=>x"6600", 1799=>x"6800",
---- 1800=>x"6e00", 1801=>x"6c00", 1802=>x"6500", 1803=>x"5d00", 1804=>x"5d00", 1805=>x"6100", 1806=>x"6700",
---- 1807=>x"6200", 1808=>x"6a00", 1809=>x"6700", 1810=>x"6000", 1811=>x"5d00", 1812=>x"5c00", 1813=>x"6600",
---- 1814=>x"6600", 1815=>x"5b00", 1816=>x"6600", 1817=>x"6000", 1818=>x"5a00", 1819=>x"5e00", 1820=>x"6300",
---- 1821=>x"6400", 1822=>x"6000", 1823=>x"5600", 1824=>x"6100", 1825=>x"5c00", 1826=>x"5900", 1827=>x"6000",
---- 1828=>x"6300", 1829=>x"6000", 1830=>x"5700", 1831=>x"4a00", 1832=>x"6000", 1833=>x"5900", 1834=>x"5c00",
---- 1835=>x"6300", 1836=>x"6300", 1837=>x"5800", 1838=>x"5000", 1839=>x"4d00", 1840=>x"5700", 1841=>x"a700",
---- 1842=>x"6000", 1843=>x"6600", 1844=>x"5d00", 1845=>x"4d00", 1846=>x"4a00", 1847=>x"5100", 1848=>x"5100",
---- 1849=>x"5a00", 1850=>x"6300", 1851=>x"6100", 1852=>x"5200", 1853=>x"4700", 1854=>x"4900", 1855=>x"5200",
---- 1856=>x"5400", 1857=>x"6000", 1858=>x"6200", 1859=>x"5a00", 1860=>x"4800", 1861=>x"4700", 1862=>x"5400",
---- 1863=>x"5f00", 1864=>x"5a00", 1865=>x"6000", 1866=>x"5d00", 1867=>x"5100", 1868=>x"4700", 1869=>x"4f00",
---- 1870=>x"6000", 1871=>x"6600", 1872=>x"5a00", 1873=>x"5700", 1874=>x"5200", 1875=>x"4c00", 1876=>x"4e00",
---- 1877=>x"5a00", 1878=>x"6800", 1879=>x"6a00", 1880=>x"5400", 1881=>x"4a00", 1882=>x"4d00", 1883=>x"ad00",
---- 1884=>x"5a00", 1885=>x"6700", 1886=>x"6d00", 1887=>x"6600", 1888=>x"4f00", 1889=>x"4b00", 1890=>x"4e00",
---- 1891=>x"5d00", 1892=>x"6300", 1893=>x"6b00", 1894=>x"6c00", 1895=>x"6200", 1896=>x"4900", 1897=>x"4300",
---- 1898=>x"4f00", 1899=>x"5e00", 1900=>x"6700", 1901=>x"6b00", 1902=>x"6500", 1903=>x"5d00", 1904=>x"4600",
---- 1905=>x"4c00", 1906=>x"5a00", 1907=>x"6600", 1908=>x"7300", 1909=>x"6900", 1910=>x"5700", 1911=>x"5500",
---- 1912=>x"4a00", 1913=>x"5a00", 1914=>x"6600", 1915=>x"6d00", 1916=>x"6900", 1917=>x"5d00", 1918=>x"5500",
---- 1919=>x"5000", 1920=>x"5200", 1921=>x"6100", 1922=>x"6c00", 1923=>x"6900", 1924=>x"6100", 1925=>x"5200",
---- 1926=>x"4b00", 1927=>x"4d00", 1928=>x"6000", 1929=>x"6600", 1930=>x"6800", 1931=>x"5f00", 1932=>x"5b00",
---- 1933=>x"5100", 1934=>x"4900", 1935=>x"4d00", 1936=>x"6900", 1937=>x"6c00", 1938=>x"6600", 1939=>x"5d00",
---- 1940=>x"5000", 1941=>x"4e00", 1942=>x"4b00", 1943=>x"4c00", 1944=>x"6a00", 1945=>x"6700", 1946=>x"6200",
---- 1947=>x"5700", 1948=>x"4900", 1949=>x"4700", 1950=>x"4700", 1951=>x"4d00", 1952=>x"6a00", 1953=>x"6000",
---- 1954=>x"5700", 1955=>x"4f00", 1956=>x"4500", 1957=>x"4200", 1958=>x"4100", 1959=>x"4c00", 1960=>x"6200",
---- 1961=>x"5700", 1962=>x"4c00", 1963=>x"4f00", 1964=>x"4700", 1965=>x"3f00", 1966=>x"4200", 1967=>x"4f00",
---- 1968=>x"5700", 1969=>x"4d00", 1970=>x"4600", 1971=>x"4500", 1972=>x"4000", 1973=>x"3f00", 1974=>x"4800",
---- 1975=>x"5c00", 1976=>x"4f00", 1977=>x"4800", 1978=>x"4500", 1979=>x"4100", 1980=>x"3c00", 1981=>x"4200",
---- 1982=>x"5400", 1983=>x"6700", 1984=>x"4f00", 1985=>x"4f00", 1986=>x"4800", 1987=>x"4200", 1988=>x"4000",
---- 1989=>x"4b00", 1990=>x"5f00", 1991=>x"6c00", 1992=>x"4b00", 1993=>x"4b00", 1994=>x"4800", 1995=>x"4700",
---- 1996=>x"4800", 1997=>x"5400", 1998=>x"6300", 1999=>x"7200", 2000=>x"4900", 2001=>x"4700", 2002=>x"4b00",
---- 2003=>x"4800", 2004=>x"5000", 2005=>x"6100", 2006=>x"6f00", 2007=>x"7400", 2008=>x"4800", 2009=>x"4800",
---- 2010=>x"4b00", 2011=>x"4f00", 2012=>x"5f00", 2013=>x"6b00", 2014=>x"7600", 2015=>x"7b00", 2016=>x"4d00",
---- 2017=>x"4a00", 2018=>x"5000", 2019=>x"5900", 2020=>x"6b00", 2021=>x"7700", 2022=>x"7c00", 2023=>x"7d00",
---- 2024=>x"4b00", 2025=>x"5000", 2026=>x"5b00", 2027=>x"6900", 2028=>x"7500", 2029=>x"8000", 2030=>x"7e00",
---- 2031=>x"7e00", 2032=>x"4f00", 2033=>x"5800", 2034=>x"6600", 2035=>x"7000", 2036=>x"7d00", 2037=>x"8100",
---- 2038=>x"7f00", 2039=>x"7e00", 2040=>x"5300", 2041=>x"5e00", 2042=>x"6500", 2043=>x"7600", 2044=>x"7f00",
---- 2045=>x"8000", 2046=>x"7f00", 2047=>x"7b00"),
---- 30 => (0=>x"7c00", 1=>x"7d00", 2=>x"7f00", 3=>x"7e00", 4=>x"8300", 5=>x"7d00", 6=>x"7e00", 7=>x"7900",
---- 8=>x"7c00", 9=>x"7d00", 10=>x"7f00", 11=>x"7e00", 12=>x"7b00", 13=>x"7d00", 14=>x"7e00",
---- 15=>x"7a00", 16=>x"7c00", 17=>x"7d00", 18=>x"7f00", 19=>x"7e00", 20=>x"7d00", 21=>x"7d00",
---- 22=>x"7d00", 23=>x"7a00", 24=>x"7a00", 25=>x"7b00", 26=>x"7e00", 27=>x"7d00", 28=>x"7c00",
---- 29=>x"7f00", 30=>x"7e00", 31=>x"7d00", 32=>x"7a00", 33=>x"7d00", 34=>x"7f00", 35=>x"7e00",
---- 36=>x"7d00", 37=>x"7e00", 38=>x"7f00", 39=>x"8100", 40=>x"7b00", 41=>x"7d00", 42=>x"7d00",
---- 43=>x"7e00", 44=>x"7e00", 45=>x"7c00", 46=>x"7f00", 47=>x"8300", 48=>x"7e00", 49=>x"7e00",
---- 50=>x"7b00", 51=>x"7b00", 52=>x"7d00", 53=>x"7d00", 54=>x"8300", 55=>x"8500", 56=>x"7d00",
---- 57=>x"7d00", 58=>x"7d00", 59=>x"8000", 60=>x"8100", 61=>x"8000", 62=>x"8700", 63=>x"8400",
---- 64=>x"8000", 65=>x"8000", 66=>x"8000", 67=>x"8300", 68=>x"8500", 69=>x"8700", 70=>x"8300",
---- 71=>x"7000", 72=>x"8100", 73=>x"8300", 74=>x"8300", 75=>x"8500", 76=>x"8800", 77=>x"8300",
---- 78=>x"6e00", 79=>x"4e00", 80=>x"8400", 81=>x"8600", 82=>x"8800", 83=>x"8b00", 84=>x"8400",
---- 85=>x"7100", 86=>x"4d00", 87=>x"3400", 88=>x"8400", 89=>x"8600", 90=>x"8a00", 91=>x"8800",
---- 92=>x"7200", 93=>x"4600", 94=>x"3400", 95=>x"2f00", 96=>x"8800", 97=>x"8700", 98=>x"8700",
---- 99=>x"7100", 100=>x"4900", 101=>x"4000", 102=>x"3600", 103=>x"2f00", 104=>x"8800", 105=>x"8700",
---- 106=>x"8f00", 107=>x"4a00", 108=>x"2f00", 109=>x"3700", 110=>x"3500", 111=>x"2800", 112=>x"8600",
---- 113=>x"6c00", 114=>x"4800", 115=>x"2b00", 116=>x"2700", 117=>x"2c00", 118=>x"2f00", 119=>x"2d00",
---- 120=>x"7000", 121=>x"4600", 122=>x"2a00", 123=>x"2c00", 124=>x"2e00", 125=>x"d100", 126=>x"2e00",
---- 127=>x"2e00", 128=>x"5000", 129=>x"3000", 130=>x"2c00", 131=>x"2800", 132=>x"3300", 133=>x"2f00",
---- 134=>x"3000", 135=>x"2b00", 136=>x"3000", 137=>x"2800", 138=>x"d400", 139=>x"2b00", 140=>x"2f00",
---- 141=>x"c700", 142=>x"3700", 143=>x"3400", 144=>x"2a00", 145=>x"2900", 146=>x"2b00", 147=>x"2d00",
---- 148=>x"3000", 149=>x"3200", 150=>x"3500", 151=>x"3800", 152=>x"2d00", 153=>x"2b00", 154=>x"2a00",
---- 155=>x"2e00", 156=>x"3700", 157=>x"3800", 158=>x"3800", 159=>x"3a00", 160=>x"2b00", 161=>x"2e00",
---- 162=>x"d300", 163=>x"2d00", 164=>x"3800", 165=>x"3b00", 166=>x"3800", 167=>x"3700", 168=>x"2c00",
---- 169=>x"2d00", 170=>x"3200", 171=>x"3500", 172=>x"3700", 173=>x"3900", 174=>x"3700", 175=>x"3400",
---- 176=>x"3000", 177=>x"3100", 178=>x"3400", 179=>x"3500", 180=>x"3900", 181=>x"3c00", 182=>x"3900",
---- 183=>x"3700", 184=>x"cf00", 185=>x"3000", 186=>x"3500", 187=>x"3700", 188=>x"3800", 189=>x"3c00",
---- 190=>x"3800", 191=>x"3600", 192=>x"3300", 193=>x"3800", 194=>x"3600", 195=>x"3800", 196=>x"c300",
---- 197=>x"3c00", 198=>x"3a00", 199=>x"3800", 200=>x"3400", 201=>x"3600", 202=>x"3500", 203=>x"3700",
---- 204=>x"3900", 205=>x"3700", 206=>x"3700", 207=>x"3800", 208=>x"3500", 209=>x"3600", 210=>x"3300",
---- 211=>x"3200", 212=>x"3400", 213=>x"3200", 214=>x"3400", 215=>x"3200", 216=>x"3700", 217=>x"3700",
---- 218=>x"3500", 219=>x"3100", 220=>x"3600", 221=>x"3300", 222=>x"2e00", 223=>x"2c00", 224=>x"3700",
---- 225=>x"3600", 226=>x"3300", 227=>x"3300", 228=>x"3400", 229=>x"2e00", 230=>x"2b00", 231=>x"3200",
---- 232=>x"3800", 233=>x"3300", 234=>x"3600", 235=>x"3600", 236=>x"3300", 237=>x"3300", 238=>x"2f00",
---- 239=>x"3100", 240=>x"3400", 241=>x"3700", 242=>x"3300", 243=>x"2e00", 244=>x"2c00", 245=>x"2e00",
---- 246=>x"3000", 247=>x"3900", 248=>x"3600", 249=>x"3500", 250=>x"2d00", 251=>x"2d00", 252=>x"2b00",
---- 253=>x"2e00", 254=>x"3700", 255=>x"3400", 256=>x"3400", 257=>x"2f00", 258=>x"2c00", 259=>x"2c00",
---- 260=>x"2c00", 261=>x"3100", 262=>x"3500", 263=>x"3400", 264=>x"3400", 265=>x"2c00", 266=>x"2a00",
---- 267=>x"2d00", 268=>x"3000", 269=>x"3400", 270=>x"3200", 271=>x"2c00", 272=>x"3000", 273=>x"2d00",
---- 274=>x"2c00", 275=>x"3300", 276=>x"3500", 277=>x"3300", 278=>x"d100", 279=>x"2b00", 280=>x"2e00",
---- 281=>x"3400", 282=>x"3500", 283=>x"3600", 284=>x"3700", 285=>x"3400", 286=>x"2d00", 287=>x"2f00",
---- 288=>x"2f00", 289=>x"3a00", 290=>x"3800", 291=>x"3100", 292=>x"3100", 293=>x"2e00", 294=>x"d300",
---- 295=>x"3300", 296=>x"3300", 297=>x"3900", 298=>x"3800", 299=>x"3400", 300=>x"3200", 301=>x"3000",
---- 302=>x"3200", 303=>x"3600", 304=>x"3700", 305=>x"3900", 306=>x"3300", 307=>x"3000", 308=>x"2e00",
---- 309=>x"3100", 310=>x"3200", 311=>x"3700", 312=>x"3700", 313=>x"3600", 314=>x"3000", 315=>x"2f00",
---- 316=>x"3200", 317=>x"3100", 318=>x"3700", 319=>x"3d00", 320=>x"3100", 321=>x"2d00", 322=>x"3200",
---- 323=>x"2d00", 324=>x"2f00", 325=>x"3300", 326=>x"3e00", 327=>x"4f00", 328=>x"2e00", 329=>x"3000",
---- 330=>x"3000", 331=>x"2d00", 332=>x"3200", 333=>x"3b00", 334=>x"4200", 335=>x"4d00", 336=>x"2c00",
---- 337=>x"2f00", 338=>x"cf00", 339=>x"3100", 340=>x"3600", 341=>x"4400", 342=>x"4b00", 343=>x"4300",
---- 344=>x"2f00", 345=>x"2f00", 346=>x"3f00", 347=>x"4400", 348=>x"3e00", 349=>x"4700", 350=>x"5100",
---- 351=>x"4100", 352=>x"2e00", 353=>x"3600", 354=>x"3f00", 355=>x"4200", 356=>x"4400", 357=>x"4800",
---- 358=>x"4c00", 359=>x"4500", 360=>x"3000", 361=>x"3c00", 362=>x"3a00", 363=>x"4000", 364=>x"4900",
---- 365=>x"4a00", 366=>x"4d00", 367=>x"5800", 368=>x"3000", 369=>x"3700", 370=>x"4000", 371=>x"4500",
---- 372=>x"4d00", 373=>x"4c00", 374=>x"5800", 375=>x"6f00", 376=>x"3300", 377=>x"3600", 378=>x"3e00",
---- 379=>x"4a00", 380=>x"4e00", 381=>x"5b00", 382=>x"7000", 383=>x"8500", 384=>x"3e00", 385=>x"3f00",
---- 386=>x"3900", 387=>x"4600", 388=>x"5900", 389=>x"7100", 390=>x"8200", 391=>x"9200", 392=>x"3b00",
---- 393=>x"3e00", 394=>x"3d00", 395=>x"4900", 396=>x"6900", 397=>x"8300", 398=>x"8e00", 399=>x"9100",
---- 400=>x"3a00", 401=>x"3e00", 402=>x"4600", 403=>x"5c00", 404=>x"7e00", 405=>x"8d00", 406=>x"9200",
---- 407=>x"8f00", 408=>x"3500", 409=>x"3e00", 410=>x"5b00", 411=>x"7b00", 412=>x"8e00", 413=>x"9000",
---- 414=>x"8c00", 415=>x"8f00", 416=>x"c500", 417=>x"5600", 418=>x"7800", 419=>x"8c00", 420=>x"9400",
---- 421=>x"8f00", 422=>x"8f00", 423=>x"8d00", 424=>x"4600", 425=>x"6e00", 426=>x"7400", 427=>x"9700",
---- 428=>x"9400", 429=>x"8d00", 430=>x"8900", 431=>x"8700", 432=>x"6800", 433=>x"8700", 434=>x"9500",
---- 435=>x"9800", 436=>x"9100", 437=>x"8d00", 438=>x"8200", 439=>x"8b00", 440=>x"8300", 441=>x"9500",
---- 442=>x"9800", 443=>x"9200", 444=>x"8e00", 445=>x"8500", 446=>x"8900", 447=>x"9a00", 448=>x"9200",
---- 449=>x"9800", 450=>x"9100", 451=>x"8c00", 452=>x"8600", 453=>x"8700", 454=>x"9400", 455=>x"9e00",
---- 456=>x"9700", 457=>x"9500", 458=>x"9000", 459=>x"8900", 460=>x"8900", 461=>x"9400", 462=>x"9c00",
---- 463=>x"a200", 464=>x"9600", 465=>x"8f00", 466=>x"8e00", 467=>x"8900", 468=>x"9300", 469=>x"9c00",
---- 470=>x"a100", 471=>x"a700", 472=>x"9300", 473=>x"8f00", 474=>x"8b00", 475=>x"8f00", 476=>x"9900",
---- 477=>x"a300", 478=>x"a300", 479=>x"a600", 480=>x"9000", 481=>x"8b00", 482=>x"8e00", 483=>x"9900",
---- 484=>x"9f00", 485=>x"a200", 486=>x"a200", 487=>x"a200", 488=>x"8b00", 489=>x"8c00", 490=>x"9800",
---- 491=>x"9e00", 492=>x"a000", 493=>x"a100", 494=>x"a000", 495=>x"a100", 496=>x"8d00", 497=>x"9400",
---- 498=>x"9e00", 499=>x"9f00", 500=>x"9e00", 501=>x"a100", 502=>x"9d00", 503=>x"a000", 504=>x"9100",
---- 505=>x"9a00", 506=>x"9f00", 507=>x"5f00", 508=>x"9b00", 509=>x"9e00", 510=>x"9e00", 511=>x"9d00",
---- 512=>x"9900", 513=>x"9f00", 514=>x"a000", 515=>x"a000", 516=>x"a000", 517=>x"9e00", 518=>x"9e00",
---- 519=>x"9e00", 520=>x"9f00", 521=>x"a100", 522=>x"a300", 523=>x"9f00", 524=>x"9f00", 525=>x"9e00",
---- 526=>x"9d00", 527=>x"9f00", 528=>x"a000", 529=>x"a200", 530=>x"a300", 531=>x"9f00", 532=>x"9e00",
---- 533=>x"9d00", 534=>x"9e00", 535=>x"9d00", 536=>x"a100", 537=>x"a000", 538=>x"9f00", 539=>x"9e00",
---- 540=>x"9d00", 541=>x"9d00", 542=>x"9b00", 543=>x"9d00", 544=>x"9f00", 545=>x"a000", 546=>x"a000",
---- 547=>x"9c00", 548=>x"9f00", 549=>x"9c00", 550=>x"9c00", 551=>x"9a00", 552=>x"a100", 553=>x"9f00",
---- 554=>x"a000", 555=>x"9d00", 556=>x"9d00", 557=>x"9e00", 558=>x"9c00", 559=>x"9b00", 560=>x"a100",
---- 561=>x"a000", 562=>x"9d00", 563=>x"9e00", 564=>x"9d00", 565=>x"9f00", 566=>x"9c00", 567=>x"9e00",
---- 568=>x"a100", 569=>x"9f00", 570=>x"a100", 571=>x"9e00", 572=>x"9d00", 573=>x"9d00", 574=>x"9d00",
---- 575=>x"a000", 576=>x"9f00", 577=>x"9e00", 578=>x"9f00", 579=>x"9c00", 580=>x"9b00", 581=>x"9c00",
---- 582=>x"9c00", 583=>x"6200", 584=>x"a000", 585=>x"9f00", 586=>x"9f00", 587=>x"9d00", 588=>x"9c00",
---- 589=>x"9d00", 590=>x"9c00", 591=>x"9e00", 592=>x"9f00", 593=>x"9f00", 594=>x"9d00", 595=>x"a000",
---- 596=>x"9c00", 597=>x"9c00", 598=>x"9c00", 599=>x"9e00", 600=>x"9e00", 601=>x"a000", 602=>x"a000",
---- 603=>x"9d00", 604=>x"9c00", 605=>x"9f00", 606=>x"9f00", 607=>x"9e00", 608=>x"a000", 609=>x"a000",
---- 610=>x"a100", 611=>x"9f00", 612=>x"9d00", 613=>x"9d00", 614=>x"9e00", 615=>x"a000", 616=>x"a000",
---- 617=>x"a100", 618=>x"a000", 619=>x"9f00", 620=>x"9d00", 621=>x"9d00", 622=>x"9c00", 623=>x"9f00",
---- 624=>x"9e00", 625=>x"a200", 626=>x"a000", 627=>x"9b00", 628=>x"9e00", 629=>x"9d00", 630=>x"9f00",
---- 631=>x"9d00", 632=>x"9f00", 633=>x"9f00", 634=>x"9f00", 635=>x"9e00", 636=>x"9d00", 637=>x"9d00",
---- 638=>x"9e00", 639=>x"6200", 640=>x"9f00", 641=>x"9e00", 642=>x"9d00", 643=>x"9f00", 644=>x"a000",
---- 645=>x"9c00", 646=>x"9b00", 647=>x"9c00", 648=>x"9f00", 649=>x"9d00", 650=>x"9f00", 651=>x"9e00",
---- 652=>x"a000", 653=>x"9c00", 654=>x"9d00", 655=>x"9d00", 656=>x"9d00", 657=>x"9d00", 658=>x"9d00",
---- 659=>x"9f00", 660=>x"9b00", 661=>x"9d00", 662=>x"9d00", 663=>x"9b00", 664=>x"9d00", 665=>x"5f00",
---- 666=>x"9f00", 667=>x"9d00", 668=>x"9b00", 669=>x"9d00", 670=>x"9d00", 671=>x"9c00", 672=>x"9b00",
---- 673=>x"9e00", 674=>x"a000", 675=>x"9e00", 676=>x"9d00", 677=>x"9c00", 678=>x"9d00", 679=>x"6400",
---- 680=>x"9c00", 681=>x"9d00", 682=>x"9c00", 683=>x"9c00", 684=>x"9c00", 685=>x"9b00", 686=>x"9c00",
---- 687=>x"9c00", 688=>x"9b00", 689=>x"9e00", 690=>x"9c00", 691=>x"9b00", 692=>x"9c00", 693=>x"9c00",
---- 694=>x"9b00", 695=>x"9c00", 696=>x"9c00", 697=>x"9d00", 698=>x"9d00", 699=>x"9b00", 700=>x"9b00",
---- 701=>x"9b00", 702=>x"9b00", 703=>x"9c00", 704=>x"9c00", 705=>x"9b00", 706=>x"9b00", 707=>x"9b00",
---- 708=>x"9b00", 709=>x"9900", 710=>x"9900", 711=>x"9900", 712=>x"9d00", 713=>x"9b00", 714=>x"9b00",
---- 715=>x"9c00", 716=>x"9c00", 717=>x"9b00", 718=>x"9a00", 719=>x"9b00", 720=>x"9e00", 721=>x"9a00",
---- 722=>x"9800", 723=>x"9a00", 724=>x"9a00", 725=>x"9c00", 726=>x"9c00", 727=>x"9a00", 728=>x"9d00",
---- 729=>x"9a00", 730=>x"6600", 731=>x"9900", 732=>x"9900", 733=>x"9a00", 734=>x"9d00", 735=>x"9b00",
---- 736=>x"9b00", 737=>x"9b00", 738=>x"9c00", 739=>x"9b00", 740=>x"9c00", 741=>x"9a00", 742=>x"9800",
---- 743=>x"9c00", 744=>x"9c00", 745=>x"9d00", 746=>x"9c00", 747=>x"9c00", 748=>x"9b00", 749=>x"9a00",
---- 750=>x"9900", 751=>x"9a00", 752=>x"9e00", 753=>x"9f00", 754=>x"9b00", 755=>x"9d00", 756=>x"9c00",
---- 757=>x"9c00", 758=>x"9c00", 759=>x"9b00", 760=>x"9f00", 761=>x"9e00", 762=>x"9c00", 763=>x"9c00",
---- 764=>x"9c00", 765=>x"9c00", 766=>x"9b00", 767=>x"9b00", 768=>x"9f00", 769=>x"9c00", 770=>x"9a00",
---- 771=>x"9b00", 772=>x"9c00", 773=>x"9c00", 774=>x"9a00", 775=>x"9d00", 776=>x"9d00", 777=>x"9d00",
---- 778=>x"9b00", 779=>x"9a00", 780=>x"9b00", 781=>x"9a00", 782=>x"9900", 783=>x"9b00", 784=>x"9e00",
---- 785=>x"9e00", 786=>x"9e00", 787=>x"9c00", 788=>x"9d00", 789=>x"9c00", 790=>x"9b00", 791=>x"9d00",
---- 792=>x"a000", 793=>x"9c00", 794=>x"9b00", 795=>x"9c00", 796=>x"9d00", 797=>x"9c00", 798=>x"9b00",
---- 799=>x"9c00", 800=>x"9e00", 801=>x"9c00", 802=>x"9c00", 803=>x"9e00", 804=>x"9e00", 805=>x"9d00",
---- 806=>x"9e00", 807=>x"9e00", 808=>x"9e00", 809=>x"9d00", 810=>x"9e00", 811=>x"9d00", 812=>x"9d00",
---- 813=>x"9e00", 814=>x"9c00", 815=>x"9c00", 816=>x"9f00", 817=>x"9f00", 818=>x"a000", 819=>x"9e00",
---- 820=>x"9e00", 821=>x"9f00", 822=>x"9d00", 823=>x"9d00", 824=>x"9e00", 825=>x"9e00", 826=>x"9f00",
---- 827=>x"9f00", 828=>x"a000", 829=>x"9f00", 830=>x"6200", 831=>x"9d00", 832=>x"9d00", 833=>x"9f00",
---- 834=>x"a000", 835=>x"a000", 836=>x"9f00", 837=>x"9e00", 838=>x"9e00", 839=>x"9c00", 840=>x"a100",
---- 841=>x"5f00", 842=>x"a100", 843=>x"6000", 844=>x"9e00", 845=>x"9d00", 846=>x"9e00", 847=>x"9e00",
---- 848=>x"a300", 849=>x"a300", 850=>x"a200", 851=>x"9f00", 852=>x"9d00", 853=>x"9b00", 854=>x"9e00",
---- 855=>x"9e00", 856=>x"a100", 857=>x"a100", 858=>x"a200", 859=>x"9f00", 860=>x"a000", 861=>x"9d00",
---- 862=>x"9d00", 863=>x"9d00", 864=>x"a200", 865=>x"a100", 866=>x"9f00", 867=>x"a000", 868=>x"a000",
---- 869=>x"9e00", 870=>x"a000", 871=>x"a000", 872=>x"a000", 873=>x"a000", 874=>x"a100", 875=>x"a000",
---- 876=>x"9d00", 877=>x"9d00", 878=>x"9d00", 879=>x"9e00", 880=>x"a100", 881=>x"9e00", 882=>x"a000",
---- 883=>x"9e00", 884=>x"9e00", 885=>x"9e00", 886=>x"9f00", 887=>x"9e00", 888=>x"a000", 889=>x"9e00",
---- 890=>x"9f00", 891=>x"9e00", 892=>x"9d00", 893=>x"9d00", 894=>x"9f00", 895=>x"9e00", 896=>x"9f00",
---- 897=>x"9f00", 898=>x"a100", 899=>x"a100", 900=>x"9c00", 901=>x"9e00", 902=>x"9d00", 903=>x"9c00",
---- 904=>x"a200", 905=>x"9f00", 906=>x"9f00", 907=>x"9e00", 908=>x"9f00", 909=>x"9d00", 910=>x"9d00",
---- 911=>x"9c00", 912=>x"a100", 913=>x"a100", 914=>x"a100", 915=>x"9d00", 916=>x"9f00", 917=>x"9d00",
---- 918=>x"9b00", 919=>x"9d00", 920=>x"a000", 921=>x"9f00", 922=>x"9e00", 923=>x"9c00", 924=>x"9c00",
---- 925=>x"9d00", 926=>x"9c00", 927=>x"9a00", 928=>x"9b00", 929=>x"6300", 930=>x"9d00", 931=>x"9d00",
---- 932=>x"9a00", 933=>x"9c00", 934=>x"9900", 935=>x"9900", 936=>x"9200", 937=>x"9600", 938=>x"6700",
---- 939=>x"9900", 940=>x"9900", 941=>x"9900", 942=>x"9900", 943=>x"9700", 944=>x"9100", 945=>x"8f00",
---- 946=>x"9200", 947=>x"8e00", 948=>x"9300", 949=>x"9500", 950=>x"9700", 951=>x"6600", 952=>x"9000",
---- 953=>x"9000", 954=>x"9000", 955=>x"8e00", 956=>x"8e00", 957=>x"8f00", 958=>x"9000", 959=>x"9300",
---- 960=>x"9100", 961=>x"8e00", 962=>x"8f00", 963=>x"8e00", 964=>x"8e00", 965=>x"9100", 966=>x"8d00",
---- 967=>x"8d00", 968=>x"9000", 969=>x"8f00", 970=>x"9000", 971=>x"9000", 972=>x"8e00", 973=>x"9000",
---- 974=>x"8e00", 975=>x"9000", 976=>x"9300", 977=>x"9200", 978=>x"9300", 979=>x"9200", 980=>x"6e00",
---- 981=>x"9000", 982=>x"9000", 983=>x"8d00", 984=>x"9500", 985=>x"9500", 986=>x"9600", 987=>x"9400",
---- 988=>x"9600", 989=>x"9100", 990=>x"8e00", 991=>x"8e00", 992=>x"9800", 993=>x"9b00", 994=>x"9900",
---- 995=>x"9800", 996=>x"9500", 997=>x"9600", 998=>x"9100", 999=>x"8f00", 1000=>x"9b00", 1001=>x"9c00",
---- 1002=>x"9c00", 1003=>x"9d00", 1004=>x"9900", 1005=>x"9900", 1006=>x"9200", 1007=>x"9200", 1008=>x"9900",
---- 1009=>x"9b00", 1010=>x"9c00", 1011=>x"9b00", 1012=>x"9a00", 1013=>x"9900", 1014=>x"6700", 1015=>x"9700",
---- 1016=>x"9a00", 1017=>x"9d00", 1018=>x"9d00", 1019=>x"9c00", 1020=>x"9e00", 1021=>x"9a00", 1022=>x"9600",
---- 1023=>x"9600", 1024=>x"9c00", 1025=>x"9b00", 1026=>x"6200", 1027=>x"9c00", 1028=>x"9a00", 1029=>x"9600",
---- 1030=>x"9400", 1031=>x"9100", 1032=>x"9a00", 1033=>x"9a00", 1034=>x"9b00", 1035=>x"9a00", 1036=>x"9a00",
---- 1037=>x"9800", 1038=>x"9200", 1039=>x"9300", 1040=>x"9900", 1041=>x"9900", 1042=>x"9800", 1043=>x"9900",
---- 1044=>x"9600", 1045=>x"9300", 1046=>x"9300", 1047=>x"9100", 1048=>x"6800", 1049=>x"9700", 1050=>x"9800",
---- 1051=>x"9700", 1052=>x"9300", 1053=>x"9100", 1054=>x"9000", 1055=>x"8f00", 1056=>x"9500", 1057=>x"9700",
---- 1058=>x"9800", 1059=>x"9200", 1060=>x"8f00", 1061=>x"8e00", 1062=>x"8e00", 1063=>x"8c00", 1064=>x"9500",
---- 1065=>x"9300", 1066=>x"9300", 1067=>x"8f00", 1068=>x"8f00", 1069=>x"8e00", 1070=>x"8d00", 1071=>x"8b00",
---- 1072=>x"9200", 1073=>x"9100", 1074=>x"8f00", 1075=>x"9000", 1076=>x"8c00", 1077=>x"8c00", 1078=>x"8b00",
---- 1079=>x"8700", 1080=>x"9100", 1081=>x"9100", 1082=>x"8e00", 1083=>x"8a00", 1084=>x"8900", 1085=>x"7600",
---- 1086=>x"8800", 1087=>x"8400", 1088=>x"8d00", 1089=>x"8d00", 1090=>x"8e00", 1091=>x"8b00", 1092=>x"8800",
---- 1093=>x"8600", 1094=>x"8500", 1095=>x"8100", 1096=>x"8900", 1097=>x"8a00", 1098=>x"8d00", 1099=>x"8a00",
---- 1100=>x"8600", 1101=>x"8400", 1102=>x"8300", 1103=>x"8600", 1104=>x"8800", 1105=>x"8800", 1106=>x"8a00",
---- 1107=>x"7700", 1108=>x"8500", 1109=>x"7900", 1110=>x"8f00", 1111=>x"9d00", 1112=>x"8800", 1113=>x"8600",
---- 1114=>x"8700", 1115=>x"8800", 1116=>x"9000", 1117=>x"9b00", 1118=>x"a500", 1119=>x"ad00", 1120=>x"8800",
---- 1121=>x"8300", 1122=>x"8900", 1123=>x"9700", 1124=>x"a300", 1125=>x"ab00", 1126=>x"b400", 1127=>x"b900",
---- 1128=>x"8400", 1129=>x"8a00", 1130=>x"9d00", 1131=>x"a900", 1132=>x"b400", 1133=>x"b900", 1134=>x"be00",
---- 1135=>x"c000", 1136=>x"8e00", 1137=>x"a600", 1138=>x"b200", 1139=>x"bd00", 1140=>x"bf00", 1141=>x"c100",
---- 1142=>x"c100", 1143=>x"c100", 1144=>x"a700", 1145=>x"b200", 1146=>x"bc00", 1147=>x"c300", 1148=>x"c500",
---- 1149=>x"c600", 1150=>x"c300", 1151=>x"c000", 1152=>x"b500", 1153=>x"bd00", 1154=>x"c200", 1155=>x"c400",
---- 1156=>x"c600", 1157=>x"c500", 1158=>x"c300", 1159=>x"c000", 1160=>x"bd00", 1161=>x"c300", 1162=>x"c600",
---- 1163=>x"c500", 1164=>x"c600", 1165=>x"c400", 1166=>x"c200", 1167=>x"c000", 1168=>x"c100", 1169=>x"c600",
---- 1170=>x"c600", 1171=>x"c400", 1172=>x"c500", 1173=>x"c300", 1174=>x"c200", 1175=>x"c100", 1176=>x"c300",
---- 1177=>x"c400", 1178=>x"c400", 1179=>x"c300", 1180=>x"c500", 1181=>x"c300", 1182=>x"c300", 1183=>x"c200",
---- 1184=>x"c200", 1185=>x"c200", 1186=>x"c200", 1187=>x"c300", 1188=>x"c400", 1189=>x"c200", 1190=>x"c100",
---- 1191=>x"c100", 1192=>x"c200", 1193=>x"c100", 1194=>x"c100", 1195=>x"c100", 1196=>x"c400", 1197=>x"c300",
---- 1198=>x"c200", 1199=>x"c300", 1200=>x"c200", 1201=>x"c200", 1202=>x"c200", 1203=>x"c300", 1204=>x"c300",
---- 1205=>x"c300", 1206=>x"c200", 1207=>x"c300", 1208=>x"c300", 1209=>x"c100", 1210=>x"c000", 1211=>x"c200",
---- 1212=>x"c200", 1213=>x"c200", 1214=>x"c400", 1215=>x"c700", 1216=>x"c100", 1217=>x"c000", 1218=>x"c100",
---- 1219=>x"c200", 1220=>x"c300", 1221=>x"c300", 1222=>x"c600", 1223=>x"ca00", 1224=>x"c000", 1225=>x"c100",
---- 1226=>x"c100", 1227=>x"c100", 1228=>x"c500", 1229=>x"c700", 1230=>x"cc00", 1231=>x"cd00", 1232=>x"c000",
---- 1233=>x"c100", 1234=>x"c200", 1235=>x"c500", 1236=>x"c900", 1237=>x"cc00", 1238=>x"ce00", 1239=>x"d000",
---- 1240=>x"c100", 1241=>x"c200", 1242=>x"c300", 1243=>x"ca00", 1244=>x"cd00", 1245=>x"3000", 1246=>x"ce00",
---- 1247=>x"cf00", 1248=>x"c100", 1249=>x"c400", 1250=>x"c800", 1251=>x"cc00", 1252=>x"2f00", 1253=>x"d200",
---- 1254=>x"d000", 1255=>x"ce00", 1256=>x"c300", 1257=>x"c900", 1258=>x"cd00", 1259=>x"d100", 1260=>x"d100",
---- 1261=>x"d100", 1262=>x"d000", 1263=>x"ce00", 1264=>x"c700", 1265=>x"cb00", 1266=>x"ce00", 1267=>x"d100",
---- 1268=>x"d000", 1269=>x"cf00", 1270=>x"ce00", 1271=>x"cd00", 1272=>x"c800", 1273=>x"cd00", 1274=>x"d000",
---- 1275=>x"cf00", 1276=>x"cf00", 1277=>x"ce00", 1278=>x"cd00", 1279=>x"cc00", 1280=>x"ca00", 1281=>x"cd00",
---- 1282=>x"ce00", 1283=>x"cd00", 1284=>x"cf00", 1285=>x"cd00", 1286=>x"ce00", 1287=>x"ce00", 1288=>x"cd00",
---- 1289=>x"ce00", 1290=>x"cd00", 1291=>x"cd00", 1292=>x"ce00", 1293=>x"ce00", 1294=>x"d000", 1295=>x"d000",
---- 1296=>x"cd00", 1297=>x"ce00", 1298=>x"cc00", 1299=>x"cc00", 1300=>x"cf00", 1301=>x"d000", 1302=>x"d000",
---- 1303=>x"d300", 1304=>x"cf00", 1305=>x"d000", 1306=>x"d000", 1307=>x"cf00", 1308=>x"cf00", 1309=>x"cf00",
---- 1310=>x"cf00", 1311=>x"d400", 1312=>x"cf00", 1313=>x"cf00", 1314=>x"2f00", 1315=>x"cf00", 1316=>x"ce00",
---- 1317=>x"cf00", 1318=>x"2d00", 1319=>x"d400", 1320=>x"ce00", 1321=>x"ce00", 1322=>x"d000", 1323=>x"cc00",
---- 1324=>x"cf00", 1325=>x"ce00", 1326=>x"d200", 1327=>x"d100", 1328=>x"cf00", 1329=>x"d000", 1330=>x"ce00",
---- 1331=>x"ce00", 1332=>x"2e00", 1333=>x"d100", 1334=>x"d100", 1335=>x"d300", 1336=>x"cf00", 1337=>x"ce00",
---- 1338=>x"cd00", 1339=>x"ce00", 1340=>x"d000", 1341=>x"cf00", 1342=>x"d000", 1343=>x"d200", 1344=>x"ce00",
---- 1345=>x"ce00", 1346=>x"cd00", 1347=>x"ce00", 1348=>x"cf00", 1349=>x"d000", 1350=>x"d100", 1351=>x"d200",
---- 1352=>x"cf00", 1353=>x"d000", 1354=>x"d000", 1355=>x"ce00", 1356=>x"d000", 1357=>x"cf00", 1358=>x"cf00",
---- 1359=>x"d100", 1360=>x"cf00", 1361=>x"d300", 1362=>x"d000", 1363=>x"d000", 1364=>x"d100", 1365=>x"cf00",
---- 1366=>x"cf00", 1367=>x"d200", 1368=>x"d100", 1369=>x"d200", 1370=>x"d000", 1371=>x"cf00", 1372=>x"cf00",
---- 1373=>x"cf00", 1374=>x"d100", 1375=>x"d300", 1376=>x"d100", 1377=>x"d100", 1378=>x"d200", 1379=>x"d000",
---- 1380=>x"d000", 1381=>x"2f00", 1382=>x"d200", 1383=>x"d200", 1384=>x"d100", 1385=>x"d200", 1386=>x"d200",
---- 1387=>x"d000", 1388=>x"d100", 1389=>x"d100", 1390=>x"d200", 1391=>x"d300", 1392=>x"ce00", 1393=>x"d100",
---- 1394=>x"d200", 1395=>x"d000", 1396=>x"d300", 1397=>x"d300", 1398=>x"2a00", 1399=>x"d500", 1400=>x"cf00",
---- 1401=>x"d100", 1402=>x"d100", 1403=>x"2e00", 1404=>x"d300", 1405=>x"d300", 1406=>x"d300", 1407=>x"d300",
---- 1408=>x"d000", 1409=>x"d300", 1410=>x"d300", 1411=>x"d100", 1412=>x"d300", 1413=>x"d200", 1414=>x"d300",
---- 1415=>x"d500", 1416=>x"d300", 1417=>x"d400", 1418=>x"d300", 1419=>x"d400", 1420=>x"d400", 1421=>x"d500",
---- 1422=>x"d600", 1423=>x"d500", 1424=>x"d300", 1425=>x"d500", 1426=>x"2b00", 1427=>x"d500", 1428=>x"d500",
---- 1429=>x"d500", 1430=>x"d400", 1431=>x"d600", 1432=>x"d400", 1433=>x"d500", 1434=>x"d400", 1435=>x"d500",
---- 1436=>x"d600", 1437=>x"d600", 1438=>x"d500", 1439=>x"d500", 1440=>x"d600", 1441=>x"d600", 1442=>x"d600",
---- 1443=>x"2800", 1444=>x"d800", 1445=>x"d700", 1446=>x"d500", 1447=>x"d200", 1448=>x"d900", 1449=>x"d700",
---- 1450=>x"d700", 1451=>x"d600", 1452=>x"d700", 1453=>x"d500", 1454=>x"d100", 1455=>x"cf00", 1456=>x"d900",
---- 1457=>x"d800", 1458=>x"d600", 1459=>x"d400", 1460=>x"d300", 1461=>x"d000", 1462=>x"ce00", 1463=>x"cd00",
---- 1464=>x"d900", 1465=>x"d800", 1466=>x"d500", 1467=>x"2d00", 1468=>x"d100", 1469=>x"ce00", 1470=>x"cd00",
---- 1471=>x"cf00", 1472=>x"d500", 1473=>x"d500", 1474=>x"d300", 1475=>x"d100", 1476=>x"d000", 1477=>x"d000",
---- 1478=>x"d100", 1479=>x"d200", 1480=>x"d500", 1481=>x"d400", 1482=>x"d200", 1483=>x"d200", 1484=>x"d200",
---- 1485=>x"d300", 1486=>x"d400", 1487=>x"d400", 1488=>x"d500", 1489=>x"d400", 1490=>x"d400", 1491=>x"d400",
---- 1492=>x"d600", 1493=>x"d500", 1494=>x"d500", 1495=>x"d400", 1496=>x"d600", 1497=>x"d600", 1498=>x"d600",
---- 1499=>x"d500", 1500=>x"d400", 1501=>x"d400", 1502=>x"d200", 1503=>x"d200", 1504=>x"d700", 1505=>x"d700",
---- 1506=>x"d700", 1507=>x"d400", 1508=>x"d200", 1509=>x"d200", 1510=>x"d000", 1511=>x"cf00", 1512=>x"d700",
---- 1513=>x"d700", 1514=>x"d500", 1515=>x"d300", 1516=>x"d200", 1517=>x"cf00", 1518=>x"cd00", 1519=>x"cf00",
---- 1520=>x"d600", 1521=>x"d500", 1522=>x"d400", 1523=>x"d100", 1524=>x"cf00", 1525=>x"cd00", 1526=>x"ce00",
---- 1527=>x"cc00", 1528=>x"d500", 1529=>x"d400", 1530=>x"d200", 1531=>x"d000", 1532=>x"cd00", 1533=>x"ce00",
---- 1534=>x"cd00", 1535=>x"cc00", 1536=>x"d300", 1537=>x"d200", 1538=>x"d000", 1539=>x"cf00", 1540=>x"cd00",
---- 1541=>x"ca00", 1542=>x"c500", 1543=>x"c100", 1544=>x"d200", 1545=>x"d100", 1546=>x"ce00", 1547=>x"ca00",
---- 1548=>x"3800", 1549=>x"bf00", 1550=>x"b100", 1551=>x"a200", 1552=>x"d200", 1553=>x"cd00", 1554=>x"c700",
---- 1555=>x"bf00", 1556=>x"b700", 1557=>x"a700", 1558=>x"8b00", 1559=>x"6400", 1560=>x"cd00", 1561=>x"c800",
---- 1562=>x"be00", 1563=>x"b200", 1564=>x"a500", 1565=>x"8b00", 1566=>x"6200", 1567=>x"3a00", 1568=>x"c900",
---- 1569=>x"3a00", 1570=>x"ba00", 1571=>x"ab00", 1572=>x"9600", 1573=>x"7400", 1574=>x"4700", 1575=>x"3100",
---- 1576=>x"be00", 1577=>x"bb00", 1578=>x"b200", 1579=>x"a100", 1580=>x"7e00", 1581=>x"4d00", 1582=>x"2f00",
---- 1583=>x"2a00", 1584=>x"b900", 1585=>x"af00", 1586=>x"9600", 1587=>x"7200", 1588=>x"4a00", 1589=>x"2c00",
---- 1590=>x"2700", 1591=>x"2d00", 1592=>x"b100", 1593=>x"9700", 1594=>x"5f00", 1595=>x"3600", 1596=>x"d200",
---- 1597=>x"2e00", 1598=>x"3200", 1599=>x"3c00", 1600=>x"9e00", 1601=>x"6b00", 1602=>x"3100", 1603=>x"2900",
---- 1604=>x"3300", 1605=>x"3f00", 1606=>x"4300", 1607=>x"4600", 1608=>x"6f00", 1609=>x"3f00", 1610=>x"d300",
---- 1611=>x"3500", 1612=>x"4400", 1613=>x"5000", 1614=>x"4f00", 1615=>x"4b00", 1616=>x"3200", 1617=>x"2a00",
---- 1618=>x"3600", 1619=>x"4600", 1620=>x"5000", 1621=>x"4f00", 1622=>x"4f00", 1623=>x"5000", 1624=>x"2800",
---- 1625=>x"3100", 1626=>x"4d00", 1627=>x"5700", 1628=>x"5500", 1629=>x"4f00", 1630=>x"4d00", 1631=>x"4d00",
---- 1632=>x"3500", 1633=>x"4b00", 1634=>x"5c00", 1635=>x"5b00", 1636=>x"5600", 1637=>x"5400", 1638=>x"5000",
---- 1639=>x"5200", 1640=>x"4300", 1641=>x"5600", 1642=>x"5b00", 1643=>x"5a00", 1644=>x"5600", 1645=>x"5600",
---- 1646=>x"5500", 1647=>x"5a00", 1648=>x"5400", 1649=>x"5c00", 1650=>x"5900", 1651=>x"5d00", 1652=>x"6000",
---- 1653=>x"5800", 1654=>x"5500", 1655=>x"6300", 1656=>x"6100", 1657=>x"5f00", 1658=>x"5800", 1659=>x"5b00",
---- 1660=>x"5c00", 1661=>x"5b00", 1662=>x"6100", 1663=>x"6e00", 1664=>x"6200", 1665=>x"5800", 1666=>x"5a00",
---- 1667=>x"5c00", 1668=>x"5c00", 1669=>x"6000", 1670=>x"6900", 1671=>x"6e00", 1672=>x"5e00", 1673=>x"5900",
---- 1674=>x"6100", 1675=>x"5f00", 1676=>x"6200", 1677=>x"6800", 1678=>x"6f00", 1679=>x"7400", 1680=>x"5800",
---- 1681=>x"5e00", 1682=>x"6400", 1683=>x"6100", 1684=>x"6500", 1685=>x"6f00", 1686=>x"7500", 1687=>x"6f00",
---- 1688=>x"5800", 1689=>x"6200", 1690=>x"6800", 1691=>x"6900", 1692=>x"6b00", 1693=>x"7200", 1694=>x"6b00",
---- 1695=>x"6200", 1696=>x"5e00", 1697=>x"6700", 1698=>x"6800", 1699=>x"6e00", 1700=>x"7100", 1701=>x"7100",
---- 1702=>x"6600", 1703=>x"5d00", 1704=>x"6400", 1705=>x"6600", 1706=>x"6a00", 1707=>x"7000", 1708=>x"7000",
---- 1709=>x"6b00", 1710=>x"6100", 1711=>x"5a00", 1712=>x"6800", 1713=>x"6900", 1714=>x"6e00", 1715=>x"7200",
---- 1716=>x"6f00", 1717=>x"6500", 1718=>x"5b00", 1719=>x"5800", 1720=>x"6b00", 1721=>x"6f00", 1722=>x"7100",
---- 1723=>x"8c00", 1724=>x"6c00", 1725=>x"5f00", 1726=>x"5d00", 1727=>x"5b00", 1728=>x"9100", 1729=>x"7300",
---- 1730=>x"7200", 1731=>x"7400", 1732=>x"6800", 1733=>x"5c00", 1734=>x"5900", 1735=>x"5b00", 1736=>x"7000",
---- 1737=>x"7200", 1738=>x"7300", 1739=>x"6f00", 1740=>x"6300", 1741=>x"5c00", 1742=>x"5700", 1743=>x"5b00",
---- 1744=>x"6f00", 1745=>x"7300", 1746=>x"6f00", 1747=>x"6400", 1748=>x"5f00", 1749=>x"5c00", 1750=>x"5a00",
---- 1751=>x"6000", 1752=>x"7500", 1753=>x"7000", 1754=>x"6900", 1755=>x"6300", 1756=>x"5c00", 1757=>x"5b00",
---- 1758=>x"5e00", 1759=>x"6400", 1760=>x"7400", 1761=>x"7000", 1762=>x"6a00", 1763=>x"6500", 1764=>x"5c00",
---- 1765=>x"5b00", 1766=>x"a100", 1767=>x"6400", 1768=>x"7000", 1769=>x"6f00", 1770=>x"6800", 1771=>x"5c00",
---- 1772=>x"5a00", 1773=>x"5c00", 1774=>x"6000", 1775=>x"6a00", 1776=>x"6f00", 1777=>x"6800", 1778=>x"5f00",
---- 1779=>x"5c00", 1780=>x"5a00", 1781=>x"5a00", 1782=>x"6200", 1783=>x"6b00", 1784=>x"6800", 1785=>x"6300",
---- 1786=>x"5a00", 1787=>x"5600", 1788=>x"5500", 1789=>x"6000", 1790=>x"6700", 1791=>x"6900", 1792=>x"6400",
---- 1793=>x"5a00", 1794=>x"5700", 1795=>x"5500", 1796=>x"5c00", 1797=>x"6400", 1798=>x"6a00", 1799=>x"6800",
---- 1800=>x"5900", 1801=>x"4d00", 1802=>x"5600", 1803=>x"6000", 1804=>x"6600", 1805=>x"6900", 1806=>x"6500",
---- 1807=>x"9a00", 1808=>x"b700", 1809=>x"4900", 1810=>x"5900", 1811=>x"6600", 1812=>x"6900", 1813=>x"6600",
---- 1814=>x"6500", 1815=>x"6100", 1816=>x"4b00", 1817=>x"5000", 1818=>x"6000", 1819=>x"6c00", 1820=>x"6c00",
---- 1821=>x"6300", 1822=>x"6600", 1823=>x"5c00", 1824=>x"4d00", 1825=>x"5900", 1826=>x"6600", 1827=>x"6c00",
---- 1828=>x"6900", 1829=>x"6100", 1830=>x"5d00", 1831=>x"5a00", 1832=>x"5300", 1833=>x"5d00", 1834=>x"6800",
---- 1835=>x"6900", 1836=>x"6500", 1837=>x"6000", 1838=>x"5d00", 1839=>x"5600", 1840=>x"5e00", 1841=>x"6500",
---- 1842=>x"6700", 1843=>x"6300", 1844=>x"6100", 1845=>x"6100", 1846=>x"5800", 1847=>x"5900", 1848=>x"6400",
---- 1849=>x"6a00", 1850=>x"6300", 1851=>x"5f00", 1852=>x"6000", 1853=>x"5f00", 1854=>x"5900", 1855=>x"5a00",
---- 1856=>x"6b00", 1857=>x"6300", 1858=>x"5e00", 1859=>x"5f00", 1860=>x"5e00", 1861=>x"5d00", 1862=>x"5d00",
---- 1863=>x"5c00", 1864=>x"6a00", 1865=>x"6000", 1866=>x"5c00", 1867=>x"5f00", 1868=>x"5d00", 1869=>x"5b00",
---- 1870=>x"5d00", 1871=>x"6300", 1872=>x"5b00", 1873=>x"5c00", 1874=>x"5d00", 1875=>x"6000", 1876=>x"5c00",
---- 1877=>x"5900", 1878=>x"5e00", 1879=>x"6500", 1880=>x"5a00", 1881=>x"5900", 1882=>x"5a00", 1883=>x"5a00",
---- 1884=>x"5d00", 1885=>x"5a00", 1886=>x"5e00", 1887=>x"6600", 1888=>x"5b00", 1889=>x"5900", 1890=>x"5600",
---- 1891=>x"5500", 1892=>x"5a00", 1893=>x"5d00", 1894=>x"6200", 1895=>x"6700", 1896=>x"5600", 1897=>x"5500",
---- 1898=>x"5500", 1899=>x"5400", 1900=>x"5700", 1901=>x"5e00", 1902=>x"6800", 1903=>x"6a00", 1904=>x"5200",
---- 1905=>x"5400", 1906=>x"5400", 1907=>x"5200", 1908=>x"5600", 1909=>x"6300", 1910=>x"6c00", 1911=>x"7100",
---- 1912=>x"4e00", 1913=>x"5100", 1914=>x"5100", 1915=>x"5600", 1916=>x"5b00", 1917=>x"6900", 1918=>x"7300",
---- 1919=>x"6d00", 1920=>x"4d00", 1921=>x"4c00", 1922=>x"5100", 1923=>x"5c00", 1924=>x"6300", 1925=>x"6c00",
---- 1926=>x"7400", 1927=>x"6900", 1928=>x"4e00", 1929=>x"5000", 1930=>x"5300", 1931=>x"5f00", 1932=>x"6a00",
---- 1933=>x"7200", 1934=>x"6d00", 1935=>x"6300", 1936=>x"4e00", 1937=>x"5300", 1938=>x"6100", 1939=>x"6b00",
---- 1940=>x"7200", 1941=>x"7000", 1942=>x"6700", 1943=>x"5c00", 1944=>x"5100", 1945=>x"5a00", 1946=>x"6300",
---- 1947=>x"7000", 1948=>x"7300", 1949=>x"6a00", 1950=>x"6700", 1951=>x"6000", 1952=>x"5800", 1953=>x"5e00",
---- 1954=>x"6900", 1955=>x"7100", 1956=>x"6f00", 1957=>x"9400", 1958=>x"6500", 1959=>x"6100", 1960=>x"6000",
---- 1961=>x"6700", 1962=>x"7000", 1963=>x"7200", 1964=>x"7000", 1965=>x"6a00", 1966=>x"6600", 1967=>x"6200",
---- 1968=>x"6a00", 1969=>x"6f00", 1970=>x"7400", 1971=>x"7500", 1972=>x"7400", 1973=>x"6800", 1974=>x"6500",
---- 1975=>x"5d00", 1976=>x"6c00", 1977=>x"6d00", 1978=>x"7300", 1979=>x"7600", 1980=>x"7100", 1981=>x"6b00",
---- 1982=>x"6500", 1983=>x"5700", 1984=>x"6f00", 1985=>x"7400", 1986=>x"7900", 1987=>x"7300", 1988=>x"6a00",
---- 1989=>x"6800", 1990=>x"5f00", 1991=>x"4e00", 1992=>x"7300", 1993=>x"7900", 1994=>x"7900", 1995=>x"6d00",
---- 1996=>x"6b00", 1997=>x"6200", 1998=>x"5500", 1999=>x"4700", 2000=>x"7e00", 2001=>x"7d00", 2002=>x"7100",
---- 2003=>x"6b00", 2004=>x"6100", 2005=>x"5a00", 2006=>x"5000", 2007=>x"4300", 2008=>x"7a00", 2009=>x"7500",
---- 2010=>x"6d00", 2011=>x"6700", 2012=>x"5b00", 2013=>x"5300", 2014=>x"4700", 2015=>x"3f00", 2016=>x"8400",
---- 2017=>x"6f00", 2018=>x"6b00", 2019=>x"6200", 2020=>x"5600", 2021=>x"4a00", 2022=>x"3d00", 2023=>x"3600",
---- 2024=>x"7500", 2025=>x"6d00", 2026=>x"6300", 2027=>x"5800", 2028=>x"4b00", 2029=>x"3d00", 2030=>x"3a00",
---- 2031=>x"2f00", 2032=>x"7800", 2033=>x"6600", 2034=>x"5600", 2035=>x"4d00", 2036=>x"3d00", 2037=>x"3300",
---- 2038=>x"3200", 2039=>x"3100", 2040=>x"7100", 2041=>x"5e00", 2042=>x"4a00", 2043=>x"3d00", 2044=>x"3a00",
---- 2045=>x"3400", 2046=>x"2c00", 2047=>x"2b00"),
---- 31 => (0=>x"7600", 1=>x"7700", 2=>x"7500", 3=>x"7500", 4=>x"8c00", 5=>x"a900", 6=>x"ac00", 7=>x"9500",
---- 8=>x"7500", 9=>x"7600", 10=>x"7500", 11=>x"7500", 12=>x"8d00", 13=>x"a900", 14=>x"ae00",
---- 15=>x"9900", 16=>x"7600", 17=>x"7500", 18=>x"7700", 19=>x"7700", 20=>x"8c00", 21=>x"a700",
---- 22=>x"a800", 23=>x"8c00", 24=>x"7800", 25=>x"7700", 26=>x"7e00", 27=>x"7f00", 28=>x"7f00",
---- 29=>x"7700", 30=>x"6000", 31=>x"4300", 32=>x"7e00", 33=>x"7e00", 34=>x"8000", 35=>x"7a00",
---- 36=>x"5f00", 37=>x"3c00", 38=>x"2f00", 39=>x"2d00", 40=>x"8400", 41=>x"8100", 42=>x"7400",
---- 43=>x"5a00", 44=>x"3c00", 45=>x"2f00", 46=>x"2f00", 47=>x"3000", 48=>x"8500", 49=>x"7a00",
---- 50=>x"5c00", 51=>x"3c00", 52=>x"3100", 53=>x"2900", 54=>x"2e00", 55=>x"3000", 56=>x"7100",
---- 57=>x"5700", 58=>x"3600", 59=>x"3600", 60=>x"3600", 61=>x"2c00", 62=>x"3300", 63=>x"3200",
---- 64=>x"4f00", 65=>x"3200", 66=>x"2d00", 67=>x"2a00", 68=>x"2e00", 69=>x"3000", 70=>x"2d00",
---- 71=>x"2f00", 72=>x"3000", 73=>x"2c00", 74=>x"3000", 75=>x"2e00", 76=>x"3200", 77=>x"3100",
---- 78=>x"2c00", 79=>x"2f00", 80=>x"2a00", 81=>x"3200", 82=>x"3400", 83=>x"2f00", 84=>x"3300",
---- 85=>x"3000", 86=>x"2e00", 87=>x"3100", 88=>x"2f00", 89=>x"d200", 90=>x"3600", 91=>x"3300",
---- 92=>x"2e00", 93=>x"2e00", 94=>x"3100", 95=>x"3400", 96=>x"3200", 97=>x"2e00", 98=>x"2c00",
---- 99=>x"d100", 100=>x"2e00", 101=>x"3200", 102=>x"3300", 103=>x"3500", 104=>x"2800", 105=>x"2d00",
---- 106=>x"2a00", 107=>x"2e00", 108=>x"2d00", 109=>x"3200", 110=>x"3800", 111=>x"3300", 112=>x"2b00",
---- 113=>x"2e00", 114=>x"2f00", 115=>x"3000", 116=>x"2f00", 117=>x"3400", 118=>x"3200", 119=>x"3900",
---- 120=>x"3100", 121=>x"2e00", 122=>x"3200", 123=>x"3300", 124=>x"3300", 125=>x"3100", 126=>x"3200",
---- 127=>x"3800", 128=>x"3100", 129=>x"3300", 130=>x"3500", 131=>x"3200", 132=>x"3200", 133=>x"2f00",
---- 134=>x"3500", 135=>x"3900", 136=>x"3600", 137=>x"3200", 138=>x"3500", 139=>x"3300", 140=>x"3100",
---- 141=>x"3300", 142=>x"3600", 143=>x"3600", 144=>x"3200", 145=>x"3200", 146=>x"3500", 147=>x"3100",
---- 148=>x"cf00", 149=>x"3600", 150=>x"3400", 151=>x"2d00", 152=>x"3900", 153=>x"3600", 154=>x"3500",
---- 155=>x"3400", 156=>x"3200", 157=>x"2f00", 158=>x"2f00", 159=>x"3000", 160=>x"3400", 161=>x"3400",
---- 162=>x"3200", 163=>x"2f00", 164=>x"3000", 165=>x"2d00", 166=>x"2c00", 167=>x"2f00", 168=>x"3300",
---- 169=>x"3500", 170=>x"3200", 171=>x"3000", 172=>x"2f00", 173=>x"2d00", 174=>x"2e00", 175=>x"2b00",
---- 176=>x"3500", 177=>x"3300", 178=>x"3600", 179=>x"2e00", 180=>x"2b00", 181=>x"2f00", 182=>x"3100",
---- 183=>x"2c00", 184=>x"ca00", 185=>x"3200", 186=>x"3400", 187=>x"2f00", 188=>x"2c00", 189=>x"2f00",
---- 190=>x"2e00", 191=>x"2e00", 192=>x"3400", 193=>x"2d00", 194=>x"2a00", 195=>x"2b00", 196=>x"3000",
---- 197=>x"2e00", 198=>x"2f00", 199=>x"3100", 200=>x"cd00", 201=>x"2b00", 202=>x"2a00", 203=>x"2b00",
---- 204=>x"d200", 205=>x"2e00", 206=>x"2f00", 207=>x"2d00", 208=>x"2f00", 209=>x"2c00", 210=>x"2f00",
---- 211=>x"3000", 212=>x"3000", 213=>x"2a00", 214=>x"2b00", 215=>x"2c00", 216=>x"3100", 217=>x"3500",
---- 218=>x"3500", 219=>x"3100", 220=>x"3000", 221=>x"2f00", 222=>x"2c00", 223=>x"2e00", 224=>x"c900",
---- 225=>x"3700", 226=>x"3000", 227=>x"2d00", 228=>x"2d00", 229=>x"2a00", 230=>x"3000", 231=>x"3000",
---- 232=>x"3600", 233=>x"3100", 234=>x"2e00", 235=>x"3200", 236=>x"2d00", 237=>x"2d00", 238=>x"2d00",
---- 239=>x"3000", 240=>x"3300", 241=>x"3100", 242=>x"2d00", 243=>x"3300", 244=>x"3600", 245=>x"2d00",
---- 246=>x"3000", 247=>x"3300", 248=>x"3000", 249=>x"2f00", 250=>x"2a00", 251=>x"2e00", 252=>x"2f00",
---- 253=>x"2c00", 254=>x"3600", 255=>x"3700", 256=>x"3000", 257=>x"2b00", 258=>x"2c00", 259=>x"2c00",
---- 260=>x"2f00", 261=>x"3600", 262=>x"3600", 263=>x"3200", 264=>x"2e00", 265=>x"2d00", 266=>x"2f00",
---- 267=>x"3100", 268=>x"3600", 269=>x"3700", 270=>x"2d00", 271=>x"2200", 272=>x"2c00", 273=>x"2d00",
---- 274=>x"3300", 275=>x"3900", 276=>x"3b00", 277=>x"3400", 278=>x"2200", 279=>x"1d00", 280=>x"3000",
---- 281=>x"3000", 282=>x"3a00", 283=>x"4300", 284=>x"3c00", 285=>x"2600", 286=>x"1a00", 287=>x"2000",
---- 288=>x"3300", 289=>x"3b00", 290=>x"4800", 291=>x"4300", 292=>x"3100", 293=>x"2300", 294=>x"1a00",
---- 295=>x"3e00", 296=>x"3800", 297=>x"4300", 298=>x"4200", 299=>x"3100", 300=>x"2100", 301=>x"1d00",
---- 302=>x"3500", 303=>x"7a00", 304=>x"4500", 305=>x"4300", 306=>x"3200", 307=>x"2700", 308=>x"2200",
---- 309=>x"3100", 310=>x"6a00", 311=>x"9a00", 312=>x"4f00", 313=>x"4100", 314=>x"2900", 315=>x"2500",
---- 316=>x"2f00", 317=>x"5900", 318=>x"8c00", 319=>x"a300", 320=>x"5300", 321=>x"3e00", 322=>x"2900",
---- 323=>x"3000", 324=>x"5800", 325=>x"8300", 326=>x"9800", 327=>x"a600", 328=>x"4b00", 329=>x"3600",
---- 330=>x"2f00", 331=>x"5400", 332=>x"8000", 333=>x"9400", 334=>x"9b00", 335=>x"a300", 336=>x"3e00",
---- 337=>x"3c00", 338=>x"5400", 339=>x"7900", 340=>x"9000", 341=>x"9600", 342=>x"6700", 343=>x"9c00",
---- 344=>x"3e00", 345=>x"5600", 346=>x"7800", 347=>x"8b00", 348=>x"9700", 349=>x"9300", 350=>x"9200",
---- 351=>x"9700", 352=>x"5b00", 353=>x"7600", 354=>x"8b00", 355=>x"9600", 356=>x"9800", 357=>x"9100",
---- 358=>x"8e00", 359=>x"8e00", 360=>x"7100", 361=>x"8800", 362=>x"9300", 363=>x"9600", 364=>x"9c00",
---- 365=>x"8f00", 366=>x"8300", 367=>x"9100", 368=>x"8300", 369=>x"8f00", 370=>x"9300", 371=>x"9600",
---- 372=>x"9900", 373=>x"8900", 374=>x"8a00", 375=>x"9c00", 376=>x"6e00", 377=>x"9400", 378=>x"9300",
---- 379=>x"9700", 380=>x"8f00", 381=>x"8900", 382=>x"9b00", 383=>x"a400", 384=>x"9500", 385=>x"9700",
---- 386=>x"9100", 387=>x"8b00", 388=>x"8d00", 389=>x"9800", 390=>x"a000", 391=>x"a300", 392=>x"9500",
---- 393=>x"9700", 394=>x"8f00", 395=>x"8a00", 396=>x"9b00", 397=>x"a200", 398=>x"a100", 399=>x"a500",
---- 400=>x"9600", 401=>x"9700", 402=>x"8b00", 403=>x"9600", 404=>x"a300", 405=>x"a500", 406=>x"a400",
---- 407=>x"a400", 408=>x"9300", 409=>x"8d00", 410=>x"9400", 411=>x"9f00", 412=>x"a600", 413=>x"a500",
---- 414=>x"a500", 415=>x"a200", 416=>x"8800", 417=>x"8d00", 418=>x"9c00", 419=>x"a400", 420=>x"a700",
---- 421=>x"a500", 422=>x"a400", 423=>x"a300", 424=>x"8e00", 425=>x"9b00", 426=>x"a000", 427=>x"a500",
---- 428=>x"a500", 429=>x"a500", 430=>x"a400", 431=>x"a300", 432=>x"9900", 433=>x"9e00", 434=>x"a200",
---- 435=>x"a100", 436=>x"a300", 437=>x"a000", 438=>x"a400", 439=>x"a600", 440=>x"9e00", 441=>x"9e00",
---- 442=>x"a300", 443=>x"a300", 444=>x"a100", 445=>x"a200", 446=>x"a200", 447=>x"5e00", 448=>x"a000",
---- 449=>x"a200", 450=>x"a300", 451=>x"a100", 452=>x"a000", 453=>x"9e00", 454=>x"9f00", 455=>x"9f00",
---- 456=>x"a200", 457=>x"a200", 458=>x"a000", 459=>x"a000", 460=>x"a000", 461=>x"9f00", 462=>x"9e00",
---- 463=>x"9f00", 464=>x"a100", 465=>x"a100", 466=>x"a000", 467=>x"a000", 468=>x"a000", 469=>x"9e00",
---- 470=>x"9e00", 471=>x"9e00", 472=>x"a100", 473=>x"a000", 474=>x"9e00", 475=>x"9f00", 476=>x"9e00",
---- 477=>x"9d00", 478=>x"9e00", 479=>x"9e00", 480=>x"9f00", 481=>x"a000", 482=>x"a000", 483=>x"a000",
---- 484=>x"9f00", 485=>x"9e00", 486=>x"9d00", 487=>x"9d00", 488=>x"a100", 489=>x"a000", 490=>x"9e00",
---- 491=>x"9f00", 492=>x"9e00", 493=>x"9d00", 494=>x"9d00", 495=>x"9d00", 496=>x"a000", 497=>x"a000",
---- 498=>x"9e00", 499=>x"9f00", 500=>x"9e00", 501=>x"9e00", 502=>x"9e00", 503=>x"9d00", 504=>x"9f00",
---- 505=>x"9f00", 506=>x"9f00", 507=>x"9b00", 508=>x"9d00", 509=>x"9d00", 510=>x"9d00", 511=>x"9f00",
---- 512=>x"9e00", 513=>x"6300", 514=>x"9d00", 515=>x"9d00", 516=>x"9c00", 517=>x"9e00", 518=>x"9d00",
---- 519=>x"a000", 520=>x"9e00", 521=>x"9f00", 522=>x"9e00", 523=>x"9b00", 524=>x"9c00", 525=>x"9900",
---- 526=>x"6100", 527=>x"9f00", 528=>x"9e00", 529=>x"9d00", 530=>x"9c00", 531=>x"9d00", 532=>x"9c00",
---- 533=>x"9900", 534=>x"9b00", 535=>x"9c00", 536=>x"9c00", 537=>x"9b00", 538=>x"9c00", 539=>x"9a00",
---- 540=>x"9c00", 541=>x"9c00", 542=>x"9a00", 543=>x"9a00", 544=>x"9d00", 545=>x"9d00", 546=>x"9b00",
---- 547=>x"9c00", 548=>x"9b00", 549=>x"9a00", 550=>x"9a00", 551=>x"9900", 552=>x"9e00", 553=>x"9d00",
---- 554=>x"9c00", 555=>x"9b00", 556=>x"9c00", 557=>x"9900", 558=>x"9a00", 559=>x"9a00", 560=>x"9c00",
---- 561=>x"9a00", 562=>x"9c00", 563=>x"9b00", 564=>x"9c00", 565=>x"9a00", 566=>x"9a00", 567=>x"9900",
---- 568=>x"9e00", 569=>x"9a00", 570=>x"9a00", 571=>x"9800", 572=>x"9b00", 573=>x"9800", 574=>x"9800",
---- 575=>x"9a00", 576=>x"9b00", 577=>x"9900", 578=>x"9c00", 579=>x"9b00", 580=>x"6300", 581=>x"9a00",
---- 582=>x"9a00", 583=>x"9a00", 584=>x"9c00", 585=>x"6500", 586=>x"9c00", 587=>x"9c00", 588=>x"9b00",
---- 589=>x"9900", 590=>x"9b00", 591=>x"9c00", 592=>x"9c00", 593=>x"9b00", 594=>x"9b00", 595=>x"9b00",
---- 596=>x"9d00", 597=>x"9b00", 598=>x"9c00", 599=>x"9b00", 600=>x"9d00", 601=>x"9d00", 602=>x"9f00",
---- 603=>x"9a00", 604=>x"9b00", 605=>x"9c00", 606=>x"9d00", 607=>x"9c00", 608=>x"9e00", 609=>x"9e00",
---- 610=>x"9e00", 611=>x"9f00", 612=>x"9c00", 613=>x"9d00", 614=>x"a000", 615=>x"9e00", 616=>x"9d00",
---- 617=>x"9d00", 618=>x"9c00", 619=>x"a000", 620=>x"9e00", 621=>x"9d00", 622=>x"9d00", 623=>x"9d00",
---- 624=>x"9c00", 625=>x"9e00", 626=>x"9f00", 627=>x"9f00", 628=>x"9d00", 629=>x"9b00", 630=>x"9c00",
---- 631=>x"9d00", 632=>x"9e00", 633=>x"9d00", 634=>x"9f00", 635=>x"9f00", 636=>x"9e00", 637=>x"9c00",
---- 638=>x"9e00", 639=>x"9d00", 640=>x"9e00", 641=>x"9c00", 642=>x"9e00", 643=>x"9d00", 644=>x"9f00",
---- 645=>x"9b00", 646=>x"9900", 647=>x"9e00", 648=>x"9c00", 649=>x"9a00", 650=>x"9d00", 651=>x"9e00",
---- 652=>x"9c00", 653=>x"9c00", 654=>x"9f00", 655=>x"9e00", 656=>x"9e00", 657=>x"9c00", 658=>x"9f00",
---- 659=>x"9c00", 660=>x"9c00", 661=>x"9b00", 662=>x"9c00", 663=>x"9c00", 664=>x"9d00", 665=>x"9d00",
---- 666=>x"9c00", 667=>x"9c00", 668=>x"9d00", 669=>x"9c00", 670=>x"9d00", 671=>x"9d00", 672=>x"9c00",
---- 673=>x"9c00", 674=>x"9e00", 675=>x"9d00", 676=>x"9e00", 677=>x"9b00", 678=>x"9c00", 679=>x"9b00",
---- 680=>x"9c00", 681=>x"6100", 682=>x"9b00", 683=>x"9c00", 684=>x"9b00", 685=>x"9b00", 686=>x"9b00",
---- 687=>x"9a00", 688=>x"9a00", 689=>x"9d00", 690=>x"9d00", 691=>x"9c00", 692=>x"9a00", 693=>x"9a00",
---- 694=>x"9a00", 695=>x"9a00", 696=>x"9b00", 697=>x"9c00", 698=>x"9b00", 699=>x"9c00", 700=>x"6400",
---- 701=>x"9800", 702=>x"9b00", 703=>x"9a00", 704=>x"9a00", 705=>x"9b00", 706=>x"9900", 707=>x"9a00",
---- 708=>x"9a00", 709=>x"9700", 710=>x"9a00", 711=>x"9900", 712=>x"9a00", 713=>x"9a00", 714=>x"9b00",
---- 715=>x"9a00", 716=>x"9b00", 717=>x"9800", 718=>x"9c00", 719=>x"9a00", 720=>x"9b00", 721=>x"9800",
---- 722=>x"9a00", 723=>x"9900", 724=>x"9b00", 725=>x"9c00", 726=>x"9b00", 727=>x"9900", 728=>x"9a00",
---- 729=>x"9b00", 730=>x"9b00", 731=>x"9a00", 732=>x"9700", 733=>x"9900", 734=>x"9a00", 735=>x"9a00",
---- 736=>x"9c00", 737=>x"9b00", 738=>x"9a00", 739=>x"9a00", 740=>x"9a00", 741=>x"9700", 742=>x"9700",
---- 743=>x"9900", 744=>x"9900", 745=>x"9800", 746=>x"9900", 747=>x"9900", 748=>x"9900", 749=>x"9b00",
---- 750=>x"9a00", 751=>x"9900", 752=>x"9a00", 753=>x"9900", 754=>x"9c00", 755=>x"9b00", 756=>x"9c00",
---- 757=>x"9900", 758=>x"6500", 759=>x"9800", 760=>x"9a00", 761=>x"9a00", 762=>x"9b00", 763=>x"9a00",
---- 764=>x"9b00", 765=>x"9800", 766=>x"9800", 767=>x"9600", 768=>x"9b00", 769=>x"9c00", 770=>x"9b00",
---- 771=>x"9b00", 772=>x"9c00", 773=>x"9700", 774=>x"9800", 775=>x"9600", 776=>x"9d00", 777=>x"9c00",
---- 778=>x"9c00", 779=>x"9a00", 780=>x"9a00", 781=>x"9800", 782=>x"9800", 783=>x"9700", 784=>x"9b00",
---- 785=>x"9900", 786=>x"9b00", 787=>x"9900", 788=>x"9b00", 789=>x"9900", 790=>x"9800", 791=>x"9800",
---- 792=>x"9b00", 793=>x"9a00", 794=>x"9a00", 795=>x"9800", 796=>x"9a00", 797=>x"9a00", 798=>x"9a00",
---- 799=>x"9700", 800=>x"9c00", 801=>x"9b00", 802=>x"9c00", 803=>x"9900", 804=>x"9b00", 805=>x"9900",
---- 806=>x"9800", 807=>x"9700", 808=>x"9c00", 809=>x"9c00", 810=>x"9a00", 811=>x"9800", 812=>x"9900",
---- 813=>x"9800", 814=>x"9600", 815=>x"9a00", 816=>x"9d00", 817=>x"9a00", 818=>x"9b00", 819=>x"9a00",
---- 820=>x"9a00", 821=>x"9800", 822=>x"9600", 823=>x"9600", 824=>x"9d00", 825=>x"9d00", 826=>x"9b00",
---- 827=>x"9a00", 828=>x"9c00", 829=>x"9800", 830=>x"9900", 831=>x"9900", 832=>x"9b00", 833=>x"9c00",
---- 834=>x"9c00", 835=>x"9900", 836=>x"9b00", 837=>x"9900", 838=>x"9900", 839=>x"9800", 840=>x"9d00",
---- 841=>x"9c00", 842=>x"9d00", 843=>x"9900", 844=>x"9800", 845=>x"9800", 846=>x"9600", 847=>x"9700",
---- 848=>x"9c00", 849=>x"9c00", 850=>x"9d00", 851=>x"9a00", 852=>x"9b00", 853=>x"9900", 854=>x"9700",
---- 855=>x"9900", 856=>x"9e00", 857=>x"9d00", 858=>x"9c00", 859=>x"9a00", 860=>x"9b00", 861=>x"9900",
---- 862=>x"9a00", 863=>x"9800", 864=>x"9e00", 865=>x"9e00", 866=>x"9d00", 867=>x"9e00", 868=>x"9b00",
---- 869=>x"9900", 870=>x"9600", 871=>x"9700", 872=>x"9c00", 873=>x"9f00", 874=>x"9e00", 875=>x"9b00",
---- 876=>x"9c00", 877=>x"9a00", 878=>x"9900", 879=>x"9600", 880=>x"9d00", 881=>x"9e00", 882=>x"9b00",
---- 883=>x"9a00", 884=>x"9c00", 885=>x"9a00", 886=>x"9900", 887=>x"9700", 888=>x"9d00", 889=>x"6000",
---- 890=>x"9d00", 891=>x"9b00", 892=>x"9b00", 893=>x"9800", 894=>x"9900", 895=>x"9700", 896=>x"9d00",
---- 897=>x"9d00", 898=>x"9c00", 899=>x"9c00", 900=>x"9b00", 901=>x"9900", 902=>x"9600", 903=>x"9700",
---- 904=>x"9c00", 905=>x"9c00", 906=>x"9c00", 907=>x"9a00", 908=>x"9d00", 909=>x"6400", 910=>x"9900",
---- 911=>x"9700", 912=>x"9d00", 913=>x"9b00", 914=>x"9b00", 915=>x"9b00", 916=>x"9b00", 917=>x"9900",
---- 918=>x"9900", 919=>x"9600", 920=>x"9b00", 921=>x"9a00", 922=>x"9c00", 923=>x"9a00", 924=>x"9700",
---- 925=>x"9400", 926=>x"9700", 927=>x"9400", 928=>x"9a00", 929=>x"9900", 930=>x"9a00", 931=>x"9b00",
---- 932=>x"9900", 933=>x"9900", 934=>x"9800", 935=>x"9600", 936=>x"9700", 937=>x"9800", 938=>x"9800",
---- 939=>x"9b00", 940=>x"9a00", 941=>x"9800", 942=>x"9700", 943=>x"9600", 944=>x"9800", 945=>x"9500",
---- 946=>x"9a00", 947=>x"9b00", 948=>x"9a00", 949=>x"9800", 950=>x"9700", 951=>x"9700", 952=>x"9400",
---- 953=>x"9900", 954=>x"9a00", 955=>x"9800", 956=>x"9700", 957=>x"6700", 958=>x"9600", 959=>x"9500",
---- 960=>x"9000", 961=>x"9300", 962=>x"9600", 963=>x"9600", 964=>x"9600", 965=>x"9800", 966=>x"9800",
---- 967=>x"9800", 968=>x"8c00", 969=>x"8d00", 970=>x"8f00", 971=>x"9000", 972=>x"9000", 973=>x"9300",
---- 974=>x"9500", 975=>x"9600", 976=>x"8c00", 977=>x"8f00", 978=>x"8f00", 979=>x"8c00", 980=>x"8c00",
---- 981=>x"8d00", 982=>x"8c00", 983=>x"8e00", 984=>x"8d00", 985=>x"8e00", 986=>x"8d00", 987=>x"8c00",
---- 988=>x"8b00", 989=>x"8c00", 990=>x"8800", 991=>x"8800", 992=>x"8e00", 993=>x"8e00", 994=>x"8f00",
---- 995=>x"7300", 996=>x"8c00", 997=>x"8a00", 998=>x"8500", 999=>x"8600", 1000=>x"9000", 1001=>x"8f00",
---- 1002=>x"9000", 1003=>x"8b00", 1004=>x"8d00", 1005=>x"8600", 1006=>x"8600", 1007=>x"8500", 1008=>x"9400",
---- 1009=>x"9100", 1010=>x"8f00", 1011=>x"8d00", 1012=>x"8b00", 1013=>x"8700", 1014=>x"8500", 1015=>x"8400",
---- 1016=>x"9900", 1017=>x"9800", 1018=>x"9300", 1019=>x"8e00", 1020=>x"8900", 1021=>x"8700", 1022=>x"8700",
---- 1023=>x"8400", 1024=>x"9400", 1025=>x"9500", 1026=>x"9300", 1027=>x"9100", 1028=>x"9000", 1029=>x"8b00",
---- 1030=>x"8b00", 1031=>x"8800", 1032=>x"9100", 1033=>x"9100", 1034=>x"9200", 1035=>x"8e00", 1036=>x"8e00",
---- 1037=>x"8e00", 1038=>x"8a00", 1039=>x"8700", 1040=>x"9100", 1041=>x"9000", 1042=>x"9000", 1043=>x"8f00",
---- 1044=>x"8b00", 1045=>x"8b00", 1046=>x"8900", 1047=>x"8700", 1048=>x"8f00", 1049=>x"8a00", 1050=>x"8900",
---- 1051=>x"8a00", 1052=>x"8900", 1053=>x"8900", 1054=>x"8800", 1055=>x"8600", 1056=>x"8a00", 1057=>x"8900",
---- 1058=>x"8600", 1059=>x"8700", 1060=>x"8700", 1061=>x"8500", 1062=>x"8700", 1063=>x"8400", 1064=>x"8800",
---- 1065=>x"8400", 1066=>x"8700", 1067=>x"8400", 1068=>x"8300", 1069=>x"7e00", 1070=>x"7f00", 1071=>x"8300",
---- 1072=>x"7b00", 1073=>x"8400", 1074=>x"8100", 1075=>x"8000", 1076=>x"8000", 1077=>x"8500", 1078=>x"8b00",
---- 1079=>x"9700", 1080=>x"8200", 1081=>x"8000", 1082=>x"8100", 1083=>x"7c00", 1084=>x"8d00", 1085=>x"9600",
---- 1086=>x"9f00", 1087=>x"5700", 1088=>x"8200", 1089=>x"8700", 1090=>x"9100", 1091=>x"9900", 1092=>x"a100",
---- 1093=>x"a600", 1094=>x"ac00", 1095=>x"b400", 1096=>x"9300", 1097=>x"9e00", 1098=>x"a300", 1099=>x"ac00",
---- 1100=>x"b100", 1101=>x"b300", 1102=>x"b700", 1103=>x"bb00", 1104=>x"a500", 1105=>x"ae00", 1106=>x"b200",
---- 1107=>x"b500", 1108=>x"b900", 1109=>x"ba00", 1110=>x"bb00", 1111=>x"be00", 1112=>x"b300", 1113=>x"b700",
---- 1114=>x"bd00", 1115=>x"bc00", 1116=>x"bd00", 1117=>x"bc00", 1118=>x"bb00", 1119=>x"bd00", 1120=>x"bd00",
---- 1121=>x"bd00", 1122=>x"be00", 1123=>x"be00", 1124=>x"bf00", 1125=>x"be00", 1126=>x"bc00", 1127=>x"bc00",
---- 1128=>x"c000", 1129=>x"c000", 1130=>x"be00", 1131=>x"bd00", 1132=>x"be00", 1133=>x"be00", 1134=>x"bc00",
---- 1135=>x"bd00", 1136=>x"c100", 1137=>x"c000", 1138=>x"c000", 1139=>x"bd00", 1140=>x"bc00", 1141=>x"bd00",
---- 1142=>x"bd00", 1143=>x"be00", 1144=>x"bf00", 1145=>x"bf00", 1146=>x"bf00", 1147=>x"bd00", 1148=>x"bd00",
---- 1149=>x"be00", 1150=>x"bd00", 1151=>x"be00", 1152=>x"c000", 1153=>x"bf00", 1154=>x"bc00", 1155=>x"bc00",
---- 1156=>x"be00", 1157=>x"be00", 1158=>x"be00", 1159=>x"bf00", 1160=>x"c000", 1161=>x"be00", 1162=>x"bd00",
---- 1163=>x"bc00", 1164=>x"bf00", 1165=>x"c000", 1166=>x"bf00", 1167=>x"3d00", 1168=>x"be00", 1169=>x"bf00",
---- 1170=>x"be00", 1171=>x"be00", 1172=>x"c100", 1173=>x"c100", 1174=>x"c100", 1175=>x"c300", 1176=>x"c000",
---- 1177=>x"bf00", 1178=>x"bd00", 1179=>x"c000", 1180=>x"c200", 1181=>x"c500", 1182=>x"c700", 1183=>x"c700",
---- 1184=>x"c300", 1185=>x"c000", 1186=>x"c100", 1187=>x"c300", 1188=>x"c500", 1189=>x"c800", 1190=>x"c900",
---- 1191=>x"ca00", 1192=>x"c300", 1193=>x"c100", 1194=>x"c500", 1195=>x"c600", 1196=>x"cb00", 1197=>x"cb00",
---- 1198=>x"cc00", 1199=>x"cb00", 1200=>x"c500", 1201=>x"c800", 1202=>x"ca00", 1203=>x"ca00", 1204=>x"cc00",
---- 1205=>x"ce00", 1206=>x"cc00", 1207=>x"cc00", 1208=>x"ca00", 1209=>x"cb00", 1210=>x"cd00", 1211=>x"ce00",
---- 1212=>x"cc00", 1213=>x"cd00", 1214=>x"cc00", 1215=>x"cb00", 1216=>x"cc00", 1217=>x"d000", 1218=>x"d000",
---- 1219=>x"ce00", 1220=>x"cc00", 1221=>x"cb00", 1222=>x"cb00", 1223=>x"ca00", 1224=>x"d000", 1225=>x"d300",
---- 1226=>x"d100", 1227=>x"cf00", 1228=>x"cd00", 1229=>x"ca00", 1230=>x"c900", 1231=>x"c900", 1232=>x"d100",
---- 1233=>x"d100", 1234=>x"d100", 1235=>x"cf00", 1236=>x"cd00", 1237=>x"cc00", 1238=>x"ca00", 1239=>x"cb00",
---- 1240=>x"d100", 1241=>x"cf00", 1242=>x"d000", 1243=>x"d000", 1244=>x"cd00", 1245=>x"cd00", 1246=>x"cc00",
---- 1247=>x"cd00", 1248=>x"cf00", 1249=>x"ce00", 1250=>x"d100", 1251=>x"cf00", 1252=>x"cf00", 1253=>x"d000",
---- 1254=>x"ce00", 1255=>x"ce00", 1256=>x"cc00", 1257=>x"ce00", 1258=>x"ce00", 1259=>x"cf00", 1260=>x"d000",
---- 1261=>x"d000", 1262=>x"ce00", 1263=>x"cf00", 1264=>x"cc00", 1265=>x"ce00", 1266=>x"ce00", 1267=>x"ce00",
---- 1268=>x"d100", 1269=>x"d000", 1270=>x"ce00", 1271=>x"cf00", 1272=>x"cd00", 1273=>x"cd00", 1274=>x"cf00",
---- 1275=>x"cf00", 1276=>x"d000", 1277=>x"2d00", 1278=>x"d100", 1279=>x"ce00", 1280=>x"cd00", 1281=>x"ce00",
---- 1282=>x"cf00", 1283=>x"d100", 1284=>x"d000", 1285=>x"d000", 1286=>x"d000", 1287=>x"cf00", 1288=>x"cf00",
---- 1289=>x"d200", 1290=>x"d100", 1291=>x"d100", 1292=>x"d200", 1293=>x"d000", 1294=>x"d000", 1295=>x"cf00",
---- 1296=>x"d200", 1297=>x"d100", 1298=>x"d200", 1299=>x"d100", 1300=>x"d200", 1301=>x"d200", 1302=>x"cf00",
---- 1303=>x"cf00", 1304=>x"d200", 1305=>x"d100", 1306=>x"d200", 1307=>x"2c00", 1308=>x"2d00", 1309=>x"cf00",
---- 1310=>x"ce00", 1311=>x"cf00", 1312=>x"d300", 1313=>x"d100", 1314=>x"d200", 1315=>x"d200", 1316=>x"d000",
---- 1317=>x"3000", 1318=>x"cf00", 1319=>x"d000", 1320=>x"d200", 1321=>x"d200", 1322=>x"d300", 1323=>x"d100",
---- 1324=>x"d000", 1325=>x"cf00", 1326=>x"cf00", 1327=>x"d200", 1328=>x"d100", 1329=>x"d100", 1330=>x"d400",
---- 1331=>x"d100", 1332=>x"d100", 1333=>x"d200", 1334=>x"d200", 1335=>x"d300", 1336=>x"d200", 1337=>x"d200",
---- 1338=>x"d300", 1339=>x"d200", 1340=>x"d200", 1341=>x"d300", 1342=>x"d300", 1343=>x"d300", 1344=>x"d000",
---- 1345=>x"d300", 1346=>x"d300", 1347=>x"d300", 1348=>x"d200", 1349=>x"d500", 1350=>x"d400", 1351=>x"d400",
---- 1352=>x"d200", 1353=>x"d500", 1354=>x"d300", 1355=>x"d000", 1356=>x"d200", 1357=>x"d300", 1358=>x"d200",
---- 1359=>x"d400", 1360=>x"d200", 1361=>x"d500", 1362=>x"d400", 1363=>x"d100", 1364=>x"d200", 1365=>x"d300",
---- 1366=>x"d200", 1367=>x"2c00", 1368=>x"d400", 1369=>x"d300", 1370=>x"d400", 1371=>x"d400", 1372=>x"d200",
---- 1373=>x"d400", 1374=>x"d400", 1375=>x"d400", 1376=>x"d500", 1377=>x"d500", 1378=>x"d500", 1379=>x"d300",
---- 1380=>x"d400", 1381=>x"d500", 1382=>x"d500", 1383=>x"d300", 1384=>x"d500", 1385=>x"d500", 1386=>x"d700",
---- 1387=>x"d400", 1388=>x"d400", 1389=>x"d600", 1390=>x"d300", 1391=>x"d300", 1392=>x"d500", 1393=>x"d500",
---- 1394=>x"d500", 1395=>x"d500", 1396=>x"d500", 1397=>x"d400", 1398=>x"d400", 1399=>x"d600", 1400=>x"2b00",
---- 1401=>x"d600", 1402=>x"d700", 1403=>x"d500", 1404=>x"d400", 1405=>x"d600", 1406=>x"d500", 1407=>x"d500",
---- 1408=>x"d500", 1409=>x"d600", 1410=>x"d700", 1411=>x"d600", 1412=>x"d600", 1413=>x"d600", 1414=>x"d500",
---- 1415=>x"d400", 1416=>x"d600", 1417=>x"d400", 1418=>x"d500", 1419=>x"d500", 1420=>x"d300", 1421=>x"d400",
---- 1422=>x"d500", 1423=>x"d500", 1424=>x"d600", 1425=>x"d600", 1426=>x"d400", 1427=>x"d300", 1428=>x"d300",
---- 1429=>x"d300", 1430=>x"d400", 1431=>x"d200", 1432=>x"d600", 1433=>x"d300", 1434=>x"d200", 1435=>x"d200",
---- 1436=>x"d100", 1437=>x"d000", 1438=>x"cf00", 1439=>x"cf00", 1440=>x"d200", 1441=>x"d000", 1442=>x"cf00",
---- 1443=>x"cf00", 1444=>x"cf00", 1445=>x"cd00", 1446=>x"cd00", 1447=>x"cd00", 1448=>x"cf00", 1449=>x"cd00",
---- 1450=>x"cd00", 1451=>x"cc00", 1452=>x"cc00", 1453=>x"cd00", 1454=>x"cc00", 1455=>x"cb00", 1456=>x"3100",
---- 1457=>x"cd00", 1458=>x"cd00", 1459=>x"cd00", 1460=>x"ce00", 1461=>x"d100", 1462=>x"d000", 1463=>x"cf00",
---- 1464=>x"d000", 1465=>x"d000", 1466=>x"d100", 1467=>x"d100", 1468=>x"d100", 1469=>x"d100", 1470=>x"d300",
---- 1471=>x"d100", 1472=>x"2e00", 1473=>x"d000", 1474=>x"d300", 1475=>x"d200", 1476=>x"d200", 1477=>x"d400",
---- 1478=>x"2c00", 1479=>x"d500", 1480=>x"d300", 1481=>x"d300", 1482=>x"d200", 1483=>x"d200", 1484=>x"d200",
---- 1485=>x"d200", 1486=>x"d200", 1487=>x"d100", 1488=>x"d200", 1489=>x"d100", 1490=>x"d100", 1491=>x"cf00",
---- 1492=>x"d000", 1493=>x"d000", 1494=>x"ce00", 1495=>x"cf00", 1496=>x"d100", 1497=>x"d000", 1498=>x"cf00",
---- 1499=>x"cf00", 1500=>x"cf00", 1501=>x"cf00", 1502=>x"cf00", 1503=>x"cd00", 1504=>x"cf00", 1505=>x"cf00",
---- 1506=>x"cf00", 1507=>x"cf00", 1508=>x"d000", 1509=>x"cf00", 1510=>x"cd00", 1511=>x"cb00", 1512=>x"cd00",
---- 1513=>x"cb00", 1514=>x"cc00", 1515=>x"cc00", 1516=>x"cc00", 1517=>x"c900", 1518=>x"c800", 1519=>x"c300",
---- 1520=>x"cb00", 1521=>x"c900", 1522=>x"c700", 1523=>x"3900", 1524=>x"c300", 1525=>x"bc00", 1526=>x"b200",
---- 1527=>x"9900", 1528=>x"c800", 1529=>x"c400", 1530=>x"b800", 1531=>x"af00", 1532=>x"9a00", 1533=>x"7f00",
---- 1534=>x"6200", 1535=>x"4400", 1536=>x"ba00", 1537=>x"aa00", 1538=>x"8e00", 1539=>x"6700", 1540=>x"4600",
---- 1541=>x"3300", 1542=>x"2d00", 1543=>x"2a00", 1544=>x"8700", 1545=>x"6100", 1546=>x"4000", 1547=>x"2d00",
---- 1548=>x"2600", 1549=>x"2800", 1550=>x"2b00", 1551=>x"2d00", 1552=>x"3f00", 1553=>x"2e00", 1554=>x"2900",
---- 1555=>x"2a00", 1556=>x"2700", 1557=>x"2b00", 1558=>x"3300", 1559=>x"3500", 1560=>x"2a00", 1561=>x"2b00",
---- 1562=>x"2a00", 1563=>x"2c00", 1564=>x"2b00", 1565=>x"3500", 1566=>x"4400", 1567=>x"4500", 1568=>x"2a00",
---- 1569=>x"2700", 1570=>x"2a00", 1571=>x"3400", 1572=>x"3d00", 1573=>x"4900", 1574=>x"5000", 1575=>x"4d00",
---- 1576=>x"2e00", 1577=>x"3300", 1578=>x"3800", 1579=>x"4000", 1580=>x"4b00", 1581=>x"5500", 1582=>x"5200",
---- 1583=>x"4c00", 1584=>x"3600", 1585=>x"3c00", 1586=>x"4100", 1587=>x"4b00", 1588=>x"5300", 1589=>x"5700",
---- 1590=>x"5300", 1591=>x"5600", 1592=>x"3f00", 1593=>x"4000", 1594=>x"4600", 1595=>x"5100", 1596=>x"5400",
---- 1597=>x"5100", 1598=>x"5300", 1599=>x"5700", 1600=>x"4600", 1601=>x"4a00", 1602=>x"4f00", 1603=>x"5300",
---- 1604=>x"5100", 1605=>x"5400", 1606=>x"5700", 1607=>x"5500", 1608=>x"4c00", 1609=>x"4d00", 1610=>x"5400",
---- 1611=>x"5600", 1612=>x"a900", 1613=>x"5800", 1614=>x"5a00", 1615=>x"5700", 1616=>x"5200", 1617=>x"5600",
---- 1618=>x"5900", 1619=>x"5b00", 1620=>x"5e00", 1621=>x"5400", 1622=>x"5300", 1623=>x"5500", 1624=>x"5500",
---- 1625=>x"5c00", 1626=>x"5d00", 1627=>x"6100", 1628=>x"5b00", 1629=>x"5600", 1630=>x"5000", 1631=>x"5500",
---- 1632=>x"5e00", 1633=>x"6000", 1634=>x"6500", 1635=>x"6200", 1636=>x"5e00", 1637=>x"5700", 1638=>x"5100",
---- 1639=>x"5900", 1640=>x"6400", 1641=>x"6600", 1642=>x"6800", 1643=>x"5f00", 1644=>x"5a00", 1645=>x"5b00",
---- 1646=>x"5600", 1647=>x"6200", 1648=>x"6a00", 1649=>x"7100", 1650=>x"6800", 1651=>x"6200", 1652=>x"5c00",
---- 1653=>x"5500", 1654=>x"5800", 1655=>x"6000", 1656=>x"8d00", 1657=>x"7100", 1658=>x"6700", 1659=>x"6000",
---- 1660=>x"5c00", 1661=>x"5700", 1662=>x"6100", 1663=>x"6500", 1664=>x"6f00", 1665=>x"6b00", 1666=>x"6500",
---- 1667=>x"5e00", 1668=>x"5b00", 1669=>x"5d00", 1670=>x"6400", 1671=>x"6800", 1672=>x"6f00", 1673=>x"6200",
---- 1674=>x"5e00", 1675=>x"5d00", 1676=>x"5d00", 1677=>x"6500", 1678=>x"6600", 1679=>x"6600", 1680=>x"6300",
---- 1681=>x"5900", 1682=>x"5c00", 1683=>x"5d00", 1684=>x"6200", 1685=>x"6600", 1686=>x"6b00", 1687=>x"6700",
---- 1688=>x"5a00", 1689=>x"5800", 1690=>x"5b00", 1691=>x"6300", 1692=>x"6700", 1693=>x"6800", 1694=>x"6700",
---- 1695=>x"6600", 1696=>x"5700", 1697=>x"5800", 1698=>x"5b00", 1699=>x"6500", 1700=>x"6800", 1701=>x"6800",
---- 1702=>x"6400", 1703=>x"6500", 1704=>x"5800", 1705=>x"5b00", 1706=>x"6000", 1707=>x"6800", 1708=>x"6700",
---- 1709=>x"6500", 1710=>x"6400", 1711=>x"6900", 1712=>x"5b00", 1713=>x"5e00", 1714=>x"6500", 1715=>x"6a00",
---- 1716=>x"6500", 1717=>x"5e00", 1718=>x"6500", 1719=>x"6700", 1720=>x"5b00", 1721=>x"6300", 1722=>x"6600",
---- 1723=>x"6800", 1724=>x"6300", 1725=>x"6200", 1726=>x"9500", 1727=>x"6a00", 1728=>x"5e00", 1729=>x"6800",
---- 1730=>x"6800", 1731=>x"6900", 1732=>x"6500", 1733=>x"6200", 1734=>x"6700", 1735=>x"6500", 1736=>x"6500",
---- 1737=>x"6800", 1738=>x"6a00", 1739=>x"6600", 1740=>x"6600", 1741=>x"6500", 1742=>x"6800", 1743=>x"5f00",
---- 1744=>x"6800", 1745=>x"6900", 1746=>x"6800", 1747=>x"6700", 1748=>x"6700", 1749=>x"6600", 1750=>x"6800",
---- 1751=>x"5a00", 1752=>x"6a00", 1753=>x"6a00", 1754=>x"6800", 1755=>x"6500", 1756=>x"5f00", 1757=>x"6200",
---- 1758=>x"5800", 1759=>x"5600", 1760=>x"6800", 1761=>x"6800", 1762=>x"6700", 1763=>x"6100", 1764=>x"5f00",
---- 1765=>x"5b00", 1766=>x"5400", 1767=>x"5100", 1768=>x"6500", 1769=>x"6a00", 1770=>x"6400", 1771=>x"5e00",
---- 1772=>x"9f00", 1773=>x"5700", 1774=>x"5700", 1775=>x"5100", 1776=>x"6600", 1777=>x"6500", 1778=>x"6200",
---- 1779=>x"6200", 1780=>x"5d00", 1781=>x"5200", 1782=>x"5c00", 1783=>x"5800", 1784=>x"6900", 1785=>x"5d00",
---- 1786=>x"5c00", 1787=>x"6000", 1788=>x"5800", 1789=>x"5900", 1790=>x"5d00", 1791=>x"5b00", 1792=>x"6700",
---- 1793=>x"5f00", 1794=>x"5e00", 1795=>x"6000", 1796=>x"5a00", 1797=>x"5900", 1798=>x"5e00", 1799=>x"5f00",
---- 1800=>x"6200", 1801=>x"5c00", 1802=>x"6200", 1803=>x"5e00", 1804=>x"5e00", 1805=>x"5c00", 1806=>x"5c00",
---- 1807=>x"6100", 1808=>x"5a00", 1809=>x"5a00", 1810=>x"5f00", 1811=>x"a300", 1812=>x"5f00", 1813=>x"5f00",
---- 1814=>x"5f00", 1815=>x"6100", 1816=>x"5800", 1817=>x"5b00", 1818=>x"5d00", 1819=>x"6000", 1820=>x"5f00",
---- 1821=>x"5f00", 1822=>x"6100", 1823=>x"5800", 1824=>x"5800", 1825=>x"5800", 1826=>x"5d00", 1827=>x"6200",
---- 1828=>x"5f00", 1829=>x"6300", 1830=>x"5e00", 1831=>x"4d00", 1832=>x"5900", 1833=>x"5a00", 1834=>x"6000",
---- 1835=>x"5e00", 1836=>x"5c00", 1837=>x"6000", 1838=>x"5900", 1839=>x"4700", 1840=>x"5e00", 1841=>x"6300",
---- 1842=>x"6500", 1843=>x"5d00", 1844=>x"5d00", 1845=>x"5900", 1846=>x"4a00", 1847=>x"3d00", 1848=>x"6300",
---- 1849=>x"6a00", 1850=>x"6300", 1851=>x"5c00", 1852=>x"5900", 1853=>x"5300", 1854=>x"4400", 1855=>x"3b00",
---- 1856=>x"6500", 1857=>x"6b00", 1858=>x"6100", 1859=>x"5e00", 1860=>x"5600", 1861=>x"4c00", 1862=>x"3c00",
---- 1863=>x"3800", 1864=>x"6800", 1865=>x"6500", 1866=>x"6100", 1867=>x"5e00", 1868=>x"4f00", 1869=>x"4500",
---- 1870=>x"3500", 1871=>x"3400", 1872=>x"6900", 1873=>x"5e00", 1874=>x"6000", 1875=>x"5a00", 1876=>x"4f00",
---- 1877=>x"4200", 1878=>x"3800", 1879=>x"3400", 1880=>x"6500", 1881=>x"6200", 1882=>x"5e00", 1883=>x"a700",
---- 1884=>x"4500", 1885=>x"3a00", 1886=>x"3800", 1887=>x"3600", 1888=>x"6400", 1889=>x"6200", 1890=>x"5a00",
---- 1891=>x"b100", 1892=>x"3d00", 1893=>x"3b00", 1894=>x"3300", 1895=>x"3200", 1896=>x"6700", 1897=>x"5f00",
---- 1898=>x"5500", 1899=>x"4600", 1900=>x"3d00", 1901=>x"3c00", 1902=>x"3400", 1903=>x"3500", 1904=>x"6600",
---- 1905=>x"5a00", 1906=>x"5400", 1907=>x"4800", 1908=>x"4700", 1909=>x"3f00", 1910=>x"3600", 1911=>x"3a00",
---- 1912=>x"6300", 1913=>x"5d00", 1914=>x"5200", 1915=>x"4d00", 1916=>x"4a00", 1917=>x"3f00", 1918=>x"3b00",
---- 1919=>x"3d00", 1920=>x"6000", 1921=>x"5700", 1922=>x"5200", 1923=>x"5500", 1924=>x"4800", 1925=>x"3c00",
---- 1926=>x"3a00", 1927=>x"4100", 1928=>x"5f00", 1929=>x"a800", 1930=>x"5000", 1931=>x"4b00", 1932=>x"4100",
---- 1933=>x"3900", 1934=>x"4400", 1935=>x"4600", 1936=>x"5e00", 1937=>x"5900", 1938=>x"4f00", 1939=>x"4700",
---- 1940=>x"3e00", 1941=>x"4100", 1942=>x"4400", 1943=>x"3d00", 1944=>x"5d00", 1945=>x"5600", 1946=>x"4c00",
---- 1947=>x"3e00", 1948=>x"3d00", 1949=>x"4700", 1950=>x"4900", 1951=>x"3e00", 1952=>x"5c00", 1953=>x"4b00",
---- 1954=>x"3f00", 1955=>x"3b00", 1956=>x"4500", 1957=>x"4500", 1958=>x"4900", 1959=>x"3e00", 1960=>x"5500",
---- 1961=>x"4400", 1962=>x"3d00", 1963=>x"4400", 1964=>x"4900", 1965=>x"4200", 1966=>x"4100", 1967=>x"3900",
---- 1968=>x"4b00", 1969=>x"4300", 1970=>x"4100", 1971=>x"3e00", 1972=>x"3f00", 1973=>x"4000", 1974=>x"3a00",
---- 1975=>x"cf00", 1976=>x"4b00", 1977=>x"4400", 1978=>x"3f00", 1979=>x"3d00", 1980=>x"3c00", 1981=>x"3c00",
---- 1982=>x"3500", 1983=>x"3400", 1984=>x"b700", 1985=>x"4100", 1986=>x"3a00", 1987=>x"3b00", 1988=>x"3e00",
---- 1989=>x"3900", 1990=>x"3600", 1991=>x"3700", 1992=>x"3e00", 1993=>x"3a00", 1994=>x"3b00", 1995=>x"3900",
---- 1996=>x"3500", 1997=>x"3400", 1998=>x"3300", 1999=>x"3000", 2000=>x"3d00", 2001=>x"3900", 2002=>x"3800",
---- 2003=>x"3b00", 2004=>x"3500", 2005=>x"3700", 2006=>x"3200", 2007=>x"3500", 2008=>x"3800", 2009=>x"3700",
---- 2010=>x"3d00", 2011=>x"3700", 2012=>x"3400", 2013=>x"3700", 2014=>x"3800", 2015=>x"4600", 2016=>x"3200",
---- 2017=>x"3300", 2018=>x"3a00", 2019=>x"c200", 2020=>x"3900", 2021=>x"3a00", 2022=>x"4700", 2023=>x"5100",
---- 2024=>x"2f00", 2025=>x"3600", 2026=>x"3400", 2027=>x"3d00", 2028=>x"4100", 2029=>x"4b00", 2030=>x"5900",
---- 2031=>x"5b00", 2032=>x"3300", 2033=>x"3200", 2034=>x"3700", 2035=>x"3c00", 2036=>x"4900", 2037=>x"5700",
---- 2038=>x"6100", 2039=>x"6100", 2040=>x"3000", 2041=>x"3300", 2042=>x"3f00", 2043=>x"4b00", 2044=>x"5700",
---- 2045=>x"6000", 2046=>x"6500", 2047=>x"6800")
---- );
--
--
---- -- 256x256 - 64 FDAs
---- constant c_PIXEL  : matrix := (
---- 0 => (0=>x"a200", 1=>x"a200", 2=>x"a000", 3=>x"a000", 4=>x"a200",
---- 5=>x"a200", 6=>x"a000", 7=>x"a000", 8=>x"a300",
---- 9=>x"a100", 10=>x"a000", 11=>x"a100", 12=>x"a200",
---- 13=>x"9f00", 14=>x"9e00", 15=>x"9e00", 16=>x"9c00",
---- 17=>x"9d00", 18=>x"9e00", 19=>x"9d00", 20=>x"9b00",
---- 21=>x"9d00", 22=>x"9d00", 23=>x"9700", 24=>x"9d00",
---- 25=>x"9d00", 26=>x"9d00", 27=>x"9a00", 28=>x"9e00",
---- 29=>x"9e00", 30=>x"9d00", 31=>x"9c00", 32=>x"9d00",
---- 33=>x"6100", 34=>x"9c00", 35=>x"9a00", 36=>x"9c00",
---- 37=>x"9c00", 38=>x"9f00", 39=>x"9a00", 40=>x"9b00",
---- 41=>x"9c00", 42=>x"9d00", 43=>x"9c00", 44=>x"9e00",
---- 45=>x"9d00", 46=>x"9900", 47=>x"9c00", 48=>x"9c00",
---- 49=>x"9a00", 50=>x"9900", 51=>x"9d00", 52=>x"9a00",
---- 53=>x"9a00", 54=>x"9900", 55=>x"9c00", 56=>x"9e00",
---- 57=>x"9e00", 58=>x"9d00", 59=>x"9d00", 60=>x"9d00",
---- 61=>x"6000", 62=>x"6000", 63=>x"9e00", 64=>x"9d00",
---- 65=>x"9f00", 66=>x"9f00", 67=>x"9c00", 68=>x"9f00",
---- 69=>x"9f00", 70=>x"9d00", 71=>x"9c00", 72=>x"a000",
---- 73=>x"9d00", 74=>x"9e00", 75=>x"6000", 76=>x"a100",
---- 77=>x"a000", 78=>x"a100", 79=>x"6100", 80=>x"a500",
---- 81=>x"a200", 82=>x"a200", 83=>x"a000", 84=>x"a000",
---- 85=>x"a000", 86=>x"a200", 87=>x"a100", 88=>x"a100",
---- 89=>x"9f00", 90=>x"a100", 91=>x"a200", 92=>x"a300",
---- 93=>x"a000", 94=>x"a200", 95=>x"a000", 96=>x"a300",
---- 97=>x"a200", 98=>x"a200", 99=>x"a100", 100=>x"a200",
---- 101=>x"a300", 102=>x"a000", 103=>x"a000", 104=>x"a100",
---- 105=>x"9f00", 106=>x"9d00", 107=>x"a100", 108=>x"a100",
---- 109=>x"a200", 110=>x"a000", 111=>x"a300", 112=>x"9e00",
---- 113=>x"a000", 114=>x"a000", 115=>x"a400", 116=>x"5f00",
---- 117=>x"5f00", 118=>x"a200", 119=>x"a600", 120=>x"a100",
---- 121=>x"a200", 122=>x"a700", 123=>x"aa00", 124=>x"a200",
---- 125=>x"a300", 126=>x"a800", 127=>x"ab00", 128=>x"a500",
---- 129=>x"a700", 130=>x"ac00", 131=>x"ae00", 132=>x"a700",
---- 133=>x"ab00", 134=>x"b000", 135=>x"ad00", 136=>x"a900",
---- 137=>x"ad00", 138=>x"ae00", 139=>x"aa00", 140=>x"ad00",
---- 141=>x"ac00", 142=>x"ab00", 143=>x"a600", 144=>x"ad00",
---- 145=>x"ab00", 146=>x"a900", 147=>x"a400", 148=>x"ad00",
---- 149=>x"ad00", 150=>x"a700", 151=>x"9f00", 152=>x"aa00",
---- 153=>x"a700", 154=>x"a300", 155=>x"9e00", 156=>x"a700",
---- 157=>x"a400", 158=>x"9f00", 159=>x"9900", 160=>x"a200",
---- 161=>x"a200", 162=>x"6600", 163=>x"9300", 164=>x"a200",
---- 165=>x"9f00", 166=>x"9700", 167=>x"8c00", 168=>x"9b00",
---- 169=>x"9900", 170=>x"9200", 171=>x"8400", 172=>x"9700",
---- 173=>x"9400", 174=>x"8900", 175=>x"7700", 176=>x"9400",
---- 177=>x"8d00", 178=>x"7e00", 179=>x"6a00", 180=>x"8b00",
---- 181=>x"7900", 182=>x"7300", 183=>x"5d00", 184=>x"8300",
---- 185=>x"7c00", 186=>x"6700", 187=>x"5500", 188=>x"7b00",
---- 189=>x"6f00", 190=>x"5800", 191=>x"5300", 192=>x"6d00",
---- 193=>x"6100", 194=>x"5100", 195=>x"5500", 196=>x"6100",
---- 197=>x"5700", 198=>x"5400", 199=>x"5600", 200=>x"5800",
---- 201=>x"5400", 202=>x"5500", 203=>x"5b00", 204=>x"5b00",
---- 205=>x"5800", 206=>x"5600", 207=>x"5c00", 208=>x"5500",
---- 209=>x"5700", 210=>x"5900", 211=>x"5d00", 212=>x"5600",
---- 213=>x"5400", 214=>x"5500", 215=>x"5d00", 216=>x"5b00",
---- 217=>x"5900", 218=>x"5a00", 219=>x"5e00", 220=>x"5b00",
---- 221=>x"5b00", 222=>x"5a00", 223=>x"5d00", 224=>x"5c00",
---- 225=>x"5f00", 226=>x"5a00", 227=>x"5b00", 228=>x"5c00",
---- 229=>x"5f00", 230=>x"5b00", 231=>x"5900", 232=>x"5700",
---- 233=>x"5900", 234=>x"5a00", 235=>x"5a00", 236=>x"5d00",
---- 237=>x"5a00", 238=>x"a700", 239=>x"5a00", 240=>x"5900",
---- 241=>x"5900", 242=>x"5900", 243=>x"5900", 244=>x"5700",
---- 245=>x"5700", 246=>x"5900", 247=>x"5900", 248=>x"5c00",
---- 249=>x"5b00", 250=>x"5a00", 251=>x"5d00", 252=>x"5d00",
---- 253=>x"5b00", 254=>x"5b00", 255=>x"5c00", 256=>x"5d00",
---- 257=>x"a300", 258=>x"5d00", 259=>x"5e00", 260=>x"5e00",
---- 261=>x"5f00", 262=>x"5f00", 263=>x"6000", 264=>x"5e00",
---- 265=>x"6300", 266=>x"6100", 267=>x"6000", 268=>x"6300",
---- 269=>x"6400", 270=>x"6300", 271=>x"6200", 272=>x"6400",
---- 273=>x"6400", 274=>x"6100", 275=>x"6300", 276=>x"6300",
---- 277=>x"6500", 278=>x"6400", 279=>x"6500", 280=>x"6300",
---- 281=>x"6300", 282=>x"6400", 283=>x"6400", 284=>x"6500",
---- 285=>x"6400", 286=>x"6300", 287=>x"6100", 288=>x"6500",
---- 289=>x"6500", 290=>x"6300", 291=>x"6300", 292=>x"6200",
---- 293=>x"6300", 294=>x"6400", 295=>x"6500", 296=>x"6500",
---- 297=>x"6300", 298=>x"6300", 299=>x"6400", 300=>x"6a00",
---- 301=>x"6500", 302=>x"6000", 303=>x"6400", 304=>x"6200",
---- 305=>x"6000", 306=>x"5f00", 307=>x"6300", 308=>x"6000",
---- 309=>x"6200", 310=>x"6500", 311=>x"6200", 312=>x"6100",
---- 313=>x"6100", 314=>x"6200", 315=>x"6100", 316=>x"6100",
---- 317=>x"6100", 318=>x"5e00", 319=>x"6400", 320=>x"6300",
---- 321=>x"6100", 322=>x"5f00", 323=>x"5e00", 324=>x"5d00",
---- 325=>x"6500", 326=>x"5f00", 327=>x"5e00", 328=>x"5f00",
---- 329=>x"6300", 330=>x"6200", 331=>x"5e00", 332=>x"5f00",
---- 333=>x"6000", 334=>x"6300", 335=>x"5e00", 336=>x"6000",
---- 337=>x"6000", 338=>x"6400", 339=>x"6200", 340=>x"5e00",
---- 341=>x"6000", 342=>x"6000", 343=>x"6000", 344=>x"6400",
---- 345=>x"6100", 346=>x"6200", 347=>x"6200", 348=>x"6300",
---- 349=>x"6300", 350=>x"6200", 351=>x"6300", 352=>x"6200",
---- 353=>x"6300", 354=>x"9f00", 355=>x"6200", 356=>x"6200",
---- 357=>x"6400", 358=>x"6200", 359=>x"6200", 360=>x"6300",
---- 361=>x"6400", 362=>x"6400", 363=>x"6600", 364=>x"6000",
---- 365=>x"6200", 366=>x"6500", 367=>x"6800", 368=>x"6100",
---- 369=>x"6400", 370=>x"6500", 371=>x"6800", 372=>x"6400",
---- 373=>x"6500", 374=>x"6600", 375=>x"6600", 376=>x"6700",
---- 377=>x"6800", 378=>x"6700", 379=>x"6800", 380=>x"6a00",
---- 381=>x"6800", 382=>x"6b00", 383=>x"9700", 384=>x"6a00",
---- 385=>x"6900", 386=>x"6900", 387=>x"6a00", 388=>x"7000",
---- 389=>x"6900", 390=>x"6600", 391=>x"6800", 392=>x"6d00",
---- 393=>x"6b00", 394=>x"6900", 395=>x"6800", 396=>x"6a00",
---- 397=>x"6b00", 398=>x"6b00", 399=>x"6800", 400=>x"6800",
---- 401=>x"6800", 402=>x"6900", 403=>x"6900", 404=>x"6f00",
---- 405=>x"6b00", 406=>x"6a00", 407=>x"6c00", 408=>x"6c00",
---- 409=>x"6d00", 410=>x"6c00", 411=>x"6d00", 412=>x"6d00",
---- 413=>x"6c00", 414=>x"6a00", 415=>x"6b00", 416=>x"6b00",
---- 417=>x"6b00", 418=>x"6c00", 419=>x"6b00", 420=>x"6b00",
---- 421=>x"6c00", 422=>x"6d00", 423=>x"6b00", 424=>x"6b00",
---- 425=>x"6c00", 426=>x"6d00", 427=>x"6900", 428=>x"6900",
---- 429=>x"6d00", 430=>x"6b00", 431=>x"6800", 432=>x"9200",
---- 433=>x"6900", 434=>x"6900", 435=>x"6900", 436=>x"6a00",
---- 437=>x"6a00", 438=>x"6600", 439=>x"6a00", 440=>x"6800",
---- 441=>x"6b00", 442=>x"6900", 443=>x"6a00", 444=>x"6600",
---- 445=>x"6800", 446=>x"6a00", 447=>x"6900", 448=>x"6500",
---- 449=>x"6600", 450=>x"6700", 451=>x"6600", 452=>x"6300",
---- 453=>x"6700", 454=>x"6a00", 455=>x"6600", 456=>x"6900",
---- 457=>x"6a00", 458=>x"6900", 459=>x"6800", 460=>x"6700",
---- 461=>x"6a00", 462=>x"6b00", 463=>x"6700", 464=>x"6900",
---- 465=>x"6900", 466=>x"6a00", 467=>x"6900", 468=>x"6700",
---- 469=>x"6a00", 470=>x"6900", 471=>x"9800", 472=>x"6500",
---- 473=>x"6700", 474=>x"6700", 475=>x"6500", 476=>x"6400",
---- 477=>x"6700", 478=>x"6600", 479=>x"6700", 480=>x"6600",
---- 481=>x"6700", 482=>x"6700", 483=>x"6600", 484=>x"6100",
---- 485=>x"6700", 486=>x"6600", 487=>x"6300", 488=>x"6600",
---- 489=>x"6700", 490=>x"6600", 491=>x"6500", 492=>x"6300",
---- 493=>x"6400", 494=>x"6300", 495=>x"6400", 496=>x"6300",
---- 497=>x"6400", 498=>x"6500", 499=>x"6400", 500=>x"9700",
---- 501=>x"6800", 502=>x"6800", 503=>x"6600", 504=>x"6500",
---- 505=>x"9b00", 506=>x"6500", 507=>x"6500", 508=>x"6200",
---- 509=>x"6500", 510=>x"6600", 511=>x"6700", 512=>x"6300",
---- 513=>x"6500", 514=>x"6400", 515=>x"6800", 516=>x"6300",
---- 517=>x"6600", 518=>x"6500", 519=>x"6500", 520=>x"6000",
---- 521=>x"6500", 522=>x"6500", 523=>x"6000", 524=>x"5e00",
---- 525=>x"5d00", 526=>x"6000", 527=>x"5f00", 528=>x"6000",
---- 529=>x"6100", 530=>x"6200", 531=>x"5f00", 532=>x"6100",
---- 533=>x"6400", 534=>x"6300", 535=>x"5f00", 536=>x"6600",
---- 537=>x"6200", 538=>x"6300", 539=>x"6100", 540=>x"6600",
---- 541=>x"6300", 542=>x"6300", 543=>x"6100", 544=>x"6200",
---- 545=>x"6500", 546=>x"6200", 547=>x"6300", 548=>x"6400",
---- 549=>x"6300", 550=>x"6600", 551=>x"6300", 552=>x"6a00",
---- 553=>x"6800", 554=>x"6400", 555=>x"6400", 556=>x"6700",
---- 557=>x"6500", 558=>x"6800", 559=>x"6a00", 560=>x"6800",
---- 561=>x"6600", 562=>x"6700", 563=>x"6700", 564=>x"6500",
---- 565=>x"6600", 566=>x"6400", 567=>x"6200", 568=>x"6600",
---- 569=>x"6400", 570=>x"6200", 571=>x"6000", 572=>x"6500",
---- 573=>x"6100", 574=>x"5d00", 575=>x"a600", 576=>x"5f00",
---- 577=>x"5d00", 578=>x"5b00", 579=>x"5900", 580=>x"5a00",
---- 581=>x"5c00", 582=>x"5e00", 583=>x"5b00", 584=>x"5a00",
---- 585=>x"5b00", 586=>x"6300", 587=>x"5a00", 588=>x"5600",
---- 589=>x"5300", 590=>x"5800", 591=>x"5800", 592=>x"5200",
---- 593=>x"5400", 594=>x"5200", 595=>x"5000", 596=>x"5400",
---- 597=>x"5100", 598=>x"4e00", 599=>x"4f00", 600=>x"5100",
---- 601=>x"5100", 602=>x"4c00", 603=>x"4b00", 604=>x"4b00",
---- 605=>x"4c00", 606=>x"4a00", 607=>x"4a00", 608=>x"4c00",
---- 609=>x"4b00", 610=>x"4d00", 611=>x"4b00", 612=>x"5300",
---- 613=>x"4d00", 614=>x"4a00", 615=>x"4c00", 616=>x"4f00",
---- 617=>x"4d00", 618=>x"4c00", 619=>x"4c00", 620=>x"4e00",
---- 621=>x"4f00", 622=>x"4d00", 623=>x"4b00", 624=>x"5000",
---- 625=>x"5200", 626=>x"5200", 627=>x"4a00", 628=>x"5100",
---- 629=>x"4f00", 630=>x"4f00", 631=>x"4c00", 632=>x"5300",
---- 633=>x"5000", 634=>x"4e00", 635=>x"4f00", 636=>x"5500",
---- 637=>x"5600", 638=>x"5300", 639=>x"5100", 640=>x"5900",
---- 641=>x"5600", 642=>x"5100", 643=>x"5000", 644=>x"5600",
---- 645=>x"5400", 646=>x"4f00", 647=>x"5100", 648=>x"4f00",
---- 649=>x"5100", 650=>x"5000", 651=>x"4f00", 652=>x"4f00",
---- 653=>x"5200", 654=>x"4e00", 655=>x"4d00", 656=>x"4c00",
---- 657=>x"5200", 658=>x"4d00", 659=>x"4f00", 660=>x"4d00",
---- 661=>x"4f00", 662=>x"4f00", 663=>x"4d00", 664=>x"4e00",
---- 665=>x"5000", 666=>x"4e00", 667=>x"4900", 668=>x"5100",
---- 669=>x"5100", 670=>x"4b00", 671=>x"4b00", 672=>x"4b00",
---- 673=>x"4c00", 674=>x"b800", 675=>x"4800", 676=>x"4800",
---- 677=>x"4a00", 678=>x"4600", 679=>x"4a00", 680=>x"4900",
---- 681=>x"4b00", 682=>x"4700", 683=>x"4800", 684=>x"4b00",
---- 685=>x"4700", 686=>x"4600", 687=>x"4500", 688=>x"4700",
---- 689=>x"4200", 690=>x"3d00", 691=>x"4100", 692=>x"4800",
---- 693=>x"4000", 694=>x"3c00", 695=>x"3d00", 696=>x"3d00",
---- 697=>x"3c00", 698=>x"3900", 699=>x"3b00", 700=>x"3800",
---- 701=>x"3700", 702=>x"c600", 703=>x"3b00", 704=>x"3800",
---- 705=>x"3800", 706=>x"3600", 707=>x"3900", 708=>x"3500",
---- 709=>x"3700", 710=>x"3a00", 711=>x"3a00", 712=>x"3800",
---- 713=>x"3800", 714=>x"3b00", 715=>x"3900", 716=>x"3600",
---- 717=>x"3800", 718=>x"3600", 719=>x"3800", 720=>x"3c00",
---- 721=>x"3700", 722=>x"3500", 723=>x"3700", 724=>x"3600",
---- 725=>x"3100", 726=>x"3400", 727=>x"3700", 728=>x"3b00",
---- 729=>x"3400", 730=>x"3000", 731=>x"3200", 732=>x"3400",
---- 733=>x"3200", 734=>x"3200", 735=>x"3700", 736=>x"3400",
---- 737=>x"3100", 738=>x"3300", 739=>x"3600", 740=>x"3800",
---- 741=>x"3300", 742=>x"3200", 743=>x"3300", 744=>x"3200",
---- 745=>x"3100", 746=>x"3000", 747=>x"3300", 748=>x"2d00",
---- 749=>x"3000", 750=>x"2f00", 751=>x"2f00", 752=>x"d100",
---- 753=>x"2f00", 754=>x"2d00", 755=>x"3100", 756=>x"2e00",
---- 757=>x"2e00", 758=>x"3200", 759=>x"3600", 760=>x"3100",
---- 761=>x"2e00", 762=>x"3200", 763=>x"3700", 764=>x"3400",
---- 765=>x"3100", 766=>x"2f00", 767=>x"2f00", 768=>x"2b00",
---- 769=>x"2b00", 770=>x"2d00", 771=>x"2f00", 772=>x"2e00",
---- 773=>x"2c00", 774=>x"2f00", 775=>x"3200", 776=>x"2f00",
---- 777=>x"2e00", 778=>x"3000", 779=>x"3200", 780=>x"3300",
---- 781=>x"3700", 782=>x"3600", 783=>x"3500", 784=>x"3800",
---- 785=>x"c800", 786=>x"3b00", 787=>x"3d00", 788=>x"3e00",
---- 789=>x"4000", 790=>x"4200", 791=>x"3e00", 792=>x"5f00",
---- 793=>x"5500", 794=>x"4a00", 795=>x"4500", 796=>x"7b00",
---- 797=>x"7500", 798=>x"6800", 799=>x"5900", 800=>x"8100",
---- 801=>x"8100", 802=>x"7e00", 803=>x"7200", 804=>x"8900",
---- 805=>x"8600", 806=>x"8400", 807=>x"8300", 808=>x"8b00",
---- 809=>x"8700", 810=>x"8b00", 811=>x"8800", 812=>x"8700",
---- 813=>x"8500", 814=>x"8b00", 815=>x"8e00", 816=>x"8000",
---- 817=>x"8300", 818=>x"8b00", 819=>x"9200", 820=>x"7c00",
---- 821=>x"8300", 822=>x"8b00", 823=>x"9100", 824=>x"8200",
---- 825=>x"7d00", 826=>x"8200", 827=>x"8e00", 828=>x"6700",
---- 829=>x"6c00", 830=>x"7a00", 831=>x"8800", 832=>x"4700",
---- 833=>x"5000", 834=>x"6e00", 835=>x"7f00", 836=>x"2e00",
---- 837=>x"3c00", 838=>x"5f00", 839=>x"7700", 840=>x"2300",
---- 841=>x"2e00", 842=>x"4c00", 843=>x"6c00", 844=>x"2300",
---- 845=>x"2800", 846=>x"3600", 847=>x"5300", 848=>x"2000",
---- 849=>x"2200", 850=>x"2a00", 851=>x"4100", 852=>x"2400",
---- 853=>x"2300", 854=>x"2a00", 855=>x"3f00", 856=>x"2000",
---- 857=>x"2700", 858=>x"2c00", 859=>x"3900", 860=>x"1f00",
---- 861=>x"2400", 862=>x"2c00", 863=>x"3c00", 864=>x"1f00",
---- 865=>x"2000", 866=>x"2200", 867=>x"cd00", 868=>x"1e00",
---- 869=>x"2100", 870=>x"2100", 871=>x"d500", 872=>x"1f00",
---- 873=>x"2000", 874=>x"1e00", 875=>x"2800", 876=>x"1e00",
---- 877=>x"2000", 878=>x"2200", 879=>x"2b00", 880=>x"1d00",
---- 881=>x"2000", 882=>x"1f00", 883=>x"2800", 884=>x"2000",
---- 885=>x"1f00", 886=>x"2000", 887=>x"2600", 888=>x"1e00",
---- 889=>x"1d00", 890=>x"2000", 891=>x"2500", 892=>x"2000",
---- 893=>x"1e00", 894=>x"2000", 895=>x"2600", 896=>x"2000",
---- 897=>x"2000", 898=>x"2100", 899=>x"2500", 900=>x"2500",
---- 901=>x"2400", 902=>x"2400", 903=>x"2800", 904=>x"2200",
---- 905=>x"2300", 906=>x"2200", 907=>x"2300", 908=>x"2800",
---- 909=>x"2700", 910=>x"2600", 911=>x"2300", 912=>x"2a00",
---- 913=>x"2900", 914=>x"2500", 915=>x"2100", 916=>x"2600",
---- 917=>x"2500", 918=>x"2400", 919=>x"2700", 920=>x"2600",
---- 921=>x"2600", 922=>x"2200", 923=>x"2400", 924=>x"2400",
---- 925=>x"2400", 926=>x"1f00", 927=>x"2400", 928=>x"2300",
---- 929=>x"2500", 930=>x"2200", 931=>x"2300", 932=>x"2100",
---- 933=>x"2100", 934=>x"2000", 935=>x"2400", 936=>x"2500",
---- 937=>x"2300", 938=>x"2200", 939=>x"1e00", 940=>x"2900",
---- 941=>x"2700", 942=>x"2200", 943=>x"2200", 944=>x"2f00",
---- 945=>x"2d00", 946=>x"2d00", 947=>x"3300", 948=>x"2f00",
---- 949=>x"3b00", 950=>x"4500", 951=>x"4400", 952=>x"4900",
---- 953=>x"5400", 954=>x"5400", 955=>x"5100", 956=>x"5d00",
---- 957=>x"5d00", 958=>x"5a00", 959=>x"5700", 960=>x"5400",
---- 961=>x"5a00", 962=>x"5a00", 963=>x"5a00", 964=>x"5500",
---- 965=>x"5a00", 966=>x"5a00", 967=>x"6000", 968=>x"4900",
---- 969=>x"5300", 970=>x"6000", 971=>x"6800", 972=>x"3b00",
---- 973=>x"4f00", 974=>x"6100", 975=>x"7000", 976=>x"3100",
---- 977=>x"4800", 978=>x"5e00", 979=>x"6c00", 980=>x"2900",
---- 981=>x"3b00", 982=>x"5000", 983=>x"5d00", 984=>x"2a00",
---- 985=>x"3500", 986=>x"4200", 987=>x"5200", 988=>x"2e00",
---- 989=>x"3300", 990=>x"3900", 991=>x"4600", 992=>x"3300",
---- 993=>x"3800", 994=>x"3500", 995=>x"3c00", 996=>x"3500",
---- 997=>x"3c00", 998=>x"3f00", 999=>x"c100", 1000=>x"3200",
---- 1001=>x"3700", 1002=>x"3b00", 1003=>x"3800", 1004=>x"3000",
---- 1005=>x"3700", 1006=>x"3900", 1007=>x"3100", 1008=>x"2f00",
---- 1009=>x"3300", 1010=>x"3500", 1011=>x"3300", 1012=>x"3200",
---- 1013=>x"3400", 1014=>x"3500", 1015=>x"3500", 1016=>x"2f00",
---- 1017=>x"3000", 1018=>x"3300", 1019=>x"3200", 1020=>x"2a00",
---- 1021=>x"3200", 1022=>x"3200", 1023=>x"3200"),
----
---- 1=> (0=>x"a300", 1=>x"a100", 2=>x"9f00", 3=>x"9f00", 4=>x"a300",
---- 5=>x"a100", 6=>x"9f00", 7=>x"9f00", 8=>x"a200",
---- 9=>x"9e00", 10=>x"9e00", 11=>x"9d00", 12=>x"9f00",
---- 13=>x"a000", 14=>x"9b00", 15=>x"9900", 16=>x"9f00",
---- 17=>x"9e00", 18=>x"9d00", 19=>x"9a00", 20=>x"9d00",
---- 21=>x"9d00", 22=>x"9d00", 23=>x"9c00", 24=>x"9d00",
---- 25=>x"9d00", 26=>x"9b00", 27=>x"9c00", 28=>x"6300",
---- 29=>x"9b00", 30=>x"9c00", 31=>x"9b00", 32=>x"9c00",
---- 33=>x"9d00", 34=>x"9c00", 35=>x"9c00", 36=>x"9c00",
---- 37=>x"9c00", 38=>x"9c00", 39=>x"9e00", 40=>x"9b00",
---- 41=>x"9d00", 42=>x"9e00", 43=>x"9e00", 44=>x"9d00",
---- 45=>x"9b00", 46=>x"9e00", 47=>x"9d00", 48=>x"9f00",
---- 49=>x"9f00", 50=>x"9d00", 51=>x"9e00", 52=>x"9e00",
---- 53=>x"9f00", 54=>x"9f00", 55=>x"9d00", 56=>x"9d00",
---- 57=>x"9f00", 58=>x"9f00", 59=>x"9d00", 60=>x"9f00",
---- 61=>x"6100", 62=>x"a100", 63=>x"9f00", 64=>x"9d00",
---- 65=>x"9e00", 66=>x"a000", 67=>x"a000", 68=>x"9d00",
---- 69=>x"9e00", 70=>x"9f00", 71=>x"a100", 72=>x"a100",
---- 73=>x"a400", 74=>x"a300", 75=>x"a100", 76=>x"a100",
---- 77=>x"a300", 78=>x"a000", 79=>x"a100", 80=>x"9f00",
---- 81=>x"a200", 82=>x"a200", 83=>x"a100", 84=>x"9f00",
---- 85=>x"a100", 86=>x"a100", 87=>x"a400", 88=>x"a000",
---- 89=>x"a000", 90=>x"a200", 91=>x"a700", 92=>x"9e00",
---- 93=>x"a100", 94=>x"a300", 95=>x"5700", 96=>x"9f00",
---- 97=>x"a200", 98=>x"a600", 99=>x"a900", 100=>x"9f00",
---- 101=>x"a300", 102=>x"aa00", 103=>x"ac00", 104=>x"a100",
---- 105=>x"a600", 106=>x"aa00", 107=>x"aa00", 108=>x"a600",
---- 109=>x"a800", 110=>x"a900", 111=>x"a700", 112=>x"a800",
---- 113=>x"ab00", 114=>x"a900", 115=>x"a500", 116=>x"aa00",
---- 117=>x"ad00", 118=>x"a700", 119=>x"a100", 120=>x"ac00",
---- 121=>x"a800", 122=>x"a400", 123=>x"9d00", 124=>x"ab00",
---- 125=>x"a700", 126=>x"a000", 127=>x"9800", 128=>x"a900",
---- 129=>x"a300", 130=>x"9d00", 131=>x"9600", 132=>x"a700",
---- 133=>x"9f00", 134=>x"9900", 135=>x"9300", 136=>x"a300",
---- 137=>x"9c00", 138=>x"9600", 139=>x"8b00", 140=>x"a000",
---- 141=>x"9a00", 142=>x"9200", 143=>x"8300", 144=>x"9e00",
---- 145=>x"9400", 146=>x"8b00", 147=>x"7e00", 148=>x"9a00",
---- 149=>x"8f00", 150=>x"8000", 151=>x"7000", 152=>x"9500",
---- 153=>x"8a00", 154=>x"7700", 155=>x"6000", 156=>x"8f00",
---- 157=>x"8100", 158=>x"6d00", 159=>x"5200", 160=>x"8600",
---- 161=>x"7600", 162=>x"6100", 163=>x"5100", 164=>x"7b00",
---- 165=>x"6a00", 166=>x"5500", 167=>x"5000", 168=>x"8e00",
---- 169=>x"5e00", 170=>x"4f00", 171=>x"5200", 172=>x"6200",
---- 173=>x"5100", 174=>x"5300", 175=>x"5600", 176=>x"5700",
---- 177=>x"5100", 178=>x"5600", 179=>x"5900", 180=>x"5300",
---- 181=>x"5400", 182=>x"5800", 183=>x"5800", 184=>x"5400",
---- 185=>x"5700", 186=>x"5d00", 187=>x"5900", 188=>x"5500",
---- 189=>x"5b00", 190=>x"6000", 191=>x"5c00", 192=>x"5700",
---- 193=>x"a500", 194=>x"5b00", 195=>x"5b00", 196=>x"5700",
---- 197=>x"5b00", 198=>x"6000", 199=>x"5d00", 200=>x"5800",
---- 201=>x"5900", 202=>x"5c00", 203=>x"5800", 204=>x"5d00",
---- 205=>x"5b00", 206=>x"5b00", 207=>x"5d00", 208=>x"5d00",
---- 209=>x"5b00", 210=>x"5d00", 211=>x"5d00", 212=>x"5d00",
---- 213=>x"5c00", 214=>x"5d00", 215=>x"5f00", 216=>x"5c00",
---- 217=>x"5c00", 218=>x"5b00", 219=>x"5a00", 220=>x"5e00",
---- 221=>x"5a00", 222=>x"5b00", 223=>x"5d00", 224=>x"5c00",
---- 225=>x"5c00", 226=>x"5d00", 227=>x"5d00", 228=>x"5b00",
---- 229=>x"5900", 230=>x"5700", 231=>x"5900", 232=>x"5a00",
---- 233=>x"5900", 234=>x"5600", 235=>x"5900", 236=>x"5800",
---- 237=>x"5700", 238=>x"5800", 239=>x"5a00", 240=>x"5a00",
---- 241=>x"5c00", 242=>x"5b00", 243=>x"5b00", 244=>x"5c00",
---- 245=>x"5a00", 246=>x"5c00", 247=>x"5e00", 248=>x"5e00",
---- 249=>x"5c00", 250=>x"a100", 251=>x"6000", 252=>x"5d00",
---- 253=>x"5c00", 254=>x"5f00", 255=>x"6000", 256=>x"5e00",
---- 257=>x"6200", 258=>x"5f00", 259=>x"5e00", 260=>x"6100",
---- 261=>x"6100", 262=>x"6400", 263=>x"6300", 264=>x"6100",
---- 265=>x"6300", 266=>x"6400", 267=>x"6100", 268=>x"6300",
---- 269=>x"6400", 270=>x"6500", 271=>x"9b00", 272=>x"6600",
---- 273=>x"6200", 274=>x"6300", 275=>x"6500", 276=>x"6700",
---- 277=>x"6300", 278=>x"6300", 279=>x"6300", 280=>x"6300",
---- 281=>x"6400", 282=>x"6500", 283=>x"6300", 284=>x"6200",
---- 285=>x"6200", 286=>x"6400", 287=>x"6200", 288=>x"6400",
---- 289=>x"6300", 290=>x"6200", 291=>x"6500", 292=>x"6700",
---- 293=>x"6500", 294=>x"6100", 295=>x"6200", 296=>x"6500",
---- 297=>x"5f00", 298=>x"6200", 299=>x"6300", 300=>x"6300",
---- 301=>x"6000", 302=>x"6100", 303=>x"6000", 304=>x"6500",
---- 305=>x"6500", 306=>x"6000", 307=>x"6000", 308=>x"9f00",
---- 309=>x"6300", 310=>x"6100", 311=>x"6000", 312=>x"6100",
---- 313=>x"6200", 314=>x"6100", 315=>x"6200", 316=>x"6000",
---- 317=>x"5d00", 318=>x"6000", 319=>x"6000", 320=>x"5d00",
---- 321=>x"5e00", 322=>x"5d00", 323=>x"6000", 324=>x"5e00",
---- 325=>x"a000", 326=>x"6000", 327=>x"5e00", 328=>x"5e00",
---- 329=>x"6100", 330=>x"6000", 331=>x"5d00", 332=>x"5b00",
---- 333=>x"5d00", 334=>x"5f00", 335=>x"5f00", 336=>x"9f00",
---- 337=>x"5f00", 338=>x"6000", 339=>x"6000", 340=>x"6500",
---- 341=>x"6100", 342=>x"5e00", 343=>x"5e00", 344=>x"5f00",
---- 345=>x"6100", 346=>x"6100", 347=>x"6100", 348=>x"6000",
---- 349=>x"6100", 350=>x"6300", 351=>x"6200", 352=>x"6300",
---- 353=>x"6100", 354=>x"6000", 355=>x"6200", 356=>x"6100",
---- 357=>x"6500", 358=>x"6100", 359=>x"6300", 360=>x"9c00",
---- 361=>x"6300", 362=>x"6200", 363=>x"6200", 364=>x"6600",
---- 365=>x"6200", 366=>x"6300", 367=>x"6300", 368=>x"6900",
---- 369=>x"6500", 370=>x"6200", 371=>x"6000", 372=>x"6600",
---- 373=>x"6500", 374=>x"6300", 375=>x"5e00", 376=>x"6700",
---- 377=>x"6400", 378=>x"6100", 379=>x"6100", 380=>x"6700",
---- 381=>x"6300", 382=>x"9f00", 383=>x"6300", 384=>x"6600",
---- 385=>x"6600", 386=>x"6700", 387=>x"6600", 388=>x"6600",
---- 389=>x"6600", 390=>x"6900", 391=>x"6300", 392=>x"6700",
---- 393=>x"6700", 394=>x"6800", 395=>x"6400", 396=>x"6800",
---- 397=>x"9600", 398=>x"6700", 399=>x"6300", 400=>x"6800",
---- 401=>x"6600", 402=>x"6400", 403=>x"6400", 404=>x"6a00",
---- 405=>x"6800", 406=>x"6700", 407=>x"6300", 408=>x"6c00",
---- 409=>x"6b00", 410=>x"6a00", 411=>x"6400", 412=>x"6900",
---- 413=>x"6600", 414=>x"6800", 415=>x"6700", 416=>x"6800",
---- 417=>x"6700", 418=>x"6800", 419=>x"9b00", 420=>x"6700",
---- 421=>x"9a00", 422=>x"6700", 423=>x"6700", 424=>x"6600",
---- 425=>x"6900", 426=>x"6600", 427=>x"6500", 428=>x"6900",
---- 429=>x"6800", 430=>x"6700", 431=>x"6400", 432=>x"6900",
---- 433=>x"6800", 434=>x"6800", 435=>x"6100", 436=>x"6a00",
---- 437=>x"6b00", 438=>x"6900", 439=>x"6500", 440=>x"6a00",
---- 441=>x"6800", 442=>x"6800", 443=>x"6600", 444=>x"6800",
---- 445=>x"6400", 446=>x"6400", 447=>x"6400", 448=>x"6900",
---- 449=>x"6800", 450=>x"6700", 451=>x"6800", 452=>x"6700",
---- 453=>x"6800", 454=>x"6700", 455=>x"6500", 456=>x"6700",
---- 457=>x"6600", 458=>x"6600", 459=>x"6600", 460=>x"6700",
---- 461=>x"6300", 462=>x"6300", 463=>x"6500", 464=>x"6600",
---- 465=>x"6000", 466=>x"6200", 467=>x"6400", 468=>x"6500",
---- 469=>x"6400", 470=>x"6400", 471=>x"6300", 472=>x"6300",
---- 473=>x"6600", 474=>x"6300", 475=>x"6300", 476=>x"6700",
---- 477=>x"6300", 478=>x"6300", 479=>x"6000", 480=>x"6600",
---- 481=>x"6300", 482=>x"6300", 483=>x"5f00", 484=>x"6500",
---- 485=>x"6200", 486=>x"6200", 487=>x"6000", 488=>x"6300",
---- 489=>x"5f00", 490=>x"6400", 491=>x"6300", 492=>x"6400",
---- 493=>x"6300", 494=>x"6300", 495=>x"6300", 496=>x"6500",
---- 497=>x"9900", 498=>x"6600", 499=>x"6400", 500=>x"6600",
---- 501=>x"6400", 502=>x"6300", 503=>x"6400", 504=>x"6700",
---- 505=>x"6a00", 506=>x"6600", 507=>x"6400", 508=>x"6800",
---- 509=>x"6800", 510=>x"6800", 511=>x"6600", 512=>x"6a00",
---- 513=>x"6600", 514=>x"6500", 515=>x"6300", 516=>x"6400",
---- 517=>x"6400", 518=>x"6200", 519=>x"6300", 520=>x"6200",
---- 521=>x"6300", 522=>x"6100", 523=>x"5f00", 524=>x"5d00",
---- 525=>x"5f00", 526=>x"5d00", 527=>x"5b00", 528=>x"5e00",
---- 529=>x"5e00", 530=>x"5d00", 531=>x"5b00", 532=>x"5f00",
---- 533=>x"5d00", 534=>x"5f00", 535=>x"5f00", 536=>x"6100",
---- 537=>x"6000", 538=>x"5f00", 539=>x"5b00", 540=>x"6100",
---- 541=>x"6100", 542=>x"9e00", 543=>x"5c00", 544=>x"6200",
---- 545=>x"6200", 546=>x"6100", 547=>x"5b00", 548=>x"6000",
---- 549=>x"6300", 550=>x"6100", 551=>x"5c00", 552=>x"6500",
---- 553=>x"6700", 554=>x"6000", 555=>x"5900", 556=>x"6400",
---- 557=>x"6500", 558=>x"5e00", 559=>x"5a00", 560=>x"6200",
---- 561=>x"6300", 562=>x"5d00", 563=>x"5900", 564=>x"5e00",
---- 565=>x"6000", 566=>x"5c00", 567=>x"5700", 568=>x"5e00",
---- 569=>x"5a00", 570=>x"5800", 571=>x"5300", 572=>x"5c00",
---- 573=>x"5800", 574=>x"5200", 575=>x"5000", 576=>x"5800",
---- 577=>x"5500", 578=>x"5300", 579=>x"5000", 580=>x"ab00",
---- 581=>x"5500", 582=>x"5400", 583=>x"5100", 584=>x"5500",
---- 585=>x"ac00", 586=>x"5200", 587=>x"5200", 588=>x"5100",
---- 589=>x"4e00", 590=>x"5100", 591=>x"5000", 592=>x"4f00",
---- 593=>x"4c00", 594=>x"4e00", 595=>x"5100", 596=>x"4e00",
---- 597=>x"4c00", 598=>x"4b00", 599=>x"4d00", 600=>x"4900",
---- 601=>x"4b00", 602=>x"4800", 603=>x"4600", 604=>x"4a00",
---- 605=>x"4c00", 606=>x"4a00", 607=>x"b600", 608=>x"4a00",
---- 609=>x"4b00", 610=>x"4e00", 611=>x"4900", 612=>x"4b00",
---- 613=>x"4c00", 614=>x"4900", 615=>x"4800", 616=>x"5000",
---- 617=>x"4d00", 618=>x"4c00", 619=>x"4900", 620=>x"4a00",
---- 621=>x"4a00", 622=>x"4b00", 623=>x"4700", 624=>x"4a00",
---- 625=>x"4700", 626=>x"4700", 627=>x"4800", 628=>x"4d00",
---- 629=>x"4b00", 630=>x"4c00", 631=>x"4a00", 632=>x"4f00",
---- 633=>x"4e00", 634=>x"4a00", 635=>x"4800", 636=>x"4f00",
---- 637=>x"4c00", 638=>x"4900", 639=>x"4500", 640=>x"5000",
---- 641=>x"4c00", 642=>x"4c00", 643=>x"4900", 644=>x"5100",
---- 645=>x"4d00", 646=>x"4b00", 647=>x"4b00", 648=>x"4c00",
---- 649=>x"4e00", 650=>x"4f00", 651=>x"4c00", 652=>x"4d00",
---- 653=>x"4e00", 654=>x"4d00", 655=>x"4900", 656=>x"4e00",
---- 657=>x"4a00", 658=>x"4a00", 659=>x"4900", 660=>x"4800",
---- 661=>x"4c00", 662=>x"5000", 663=>x"4b00", 664=>x"4e00",
---- 665=>x"4f00", 666=>x"5200", 667=>x"4c00", 668=>x"5000",
---- 669=>x"5000", 670=>x"4c00", 671=>x"4900", 672=>x"4a00",
---- 673=>x"4900", 674=>x"4c00", 675=>x"4a00", 676=>x"4800",
---- 677=>x"4700", 678=>x"4c00", 679=>x"4700", 680=>x"4600",
---- 681=>x"4300", 682=>x"4500", 683=>x"4500", 684=>x"ba00",
---- 685=>x"4400", 686=>x"4400", 687=>x"4500", 688=>x"4300",
---- 689=>x"4500", 690=>x"4600", 691=>x"4300", 692=>x"4100",
---- 693=>x"4500", 694=>x"4600", 695=>x"4400", 696=>x"3d00",
---- 697=>x"3c00", 698=>x"4200", 699=>x"4500", 700=>x"3c00",
---- 701=>x"3e00", 702=>x"4300", 703=>x"4000", 704=>x"3c00",
---- 705=>x"3e00", 706=>x"4300", 707=>x"4000", 708=>x"3b00",
---- 709=>x"3b00", 710=>x"4000", 711=>x"4000", 712=>x"3b00",
---- 713=>x"3d00", 714=>x"4200", 715=>x"4000", 716=>x"3b00",
---- 717=>x"3d00", 718=>x"3e00", 719=>x"3f00", 720=>x"3900",
---- 721=>x"3600", 722=>x"3c00", 723=>x"3b00", 724=>x"3700",
---- 725=>x"3700", 726=>x"3900", 727=>x"3700", 728=>x"3300",
---- 729=>x"3a00", 730=>x"3900", 731=>x"3900", 732=>x"3300",
---- 733=>x"3400", 734=>x"3300", 735=>x"3100", 736=>x"3300",
---- 737=>x"3200", 738=>x"3200", 739=>x"3100", 740=>x"3000",
---- 741=>x"3100", 742=>x"2f00", 743=>x"3000", 744=>x"3200",
---- 745=>x"3100", 746=>x"3000", 747=>x"2f00", 748=>x"3400",
---- 749=>x"3100", 750=>x"3200", 751=>x"3400", 752=>x"3000",
---- 753=>x"2f00", 754=>x"3200", 755=>x"3000", 756=>x"2e00",
---- 757=>x"2a00", 758=>x"3000", 759=>x"3100", 760=>x"3100",
---- 761=>x"2e00", 762=>x"3000", 763=>x"3000", 764=>x"2e00",
---- 765=>x"2c00", 766=>x"2e00", 767=>x"3000", 768=>x"3000",
---- 769=>x"2c00", 770=>x"2900", 771=>x"3000", 772=>x"2d00",
---- 773=>x"2b00", 774=>x"2c00", 775=>x"2c00", 776=>x"2c00",
---- 777=>x"2900", 778=>x"2c00", 779=>x"2900", 780=>x"3100",
---- 781=>x"d600", 782=>x"2700", 783=>x"2800", 784=>x"3200",
---- 785=>x"3000", 786=>x"2a00", 787=>x"2800", 788=>x"3700",
---- 789=>x"3300", 790=>x"3400", 791=>x"3000", 792=>x"3d00",
---- 793=>x"3700", 794=>x"3400", 795=>x"3400", 796=>x"4c00",
---- 797=>x"b900", 798=>x"3d00", 799=>x"3600", 800=>x"6000",
---- 801=>x"5500", 802=>x"4f00", 803=>x"4000", 804=>x"7600",
---- 805=>x"6800", 806=>x"5b00", 807=>x"5000", 808=>x"8200",
---- 809=>x"7b00", 810=>x"6d00", 811=>x"6100", 812=>x"8d00",
---- 813=>x"8900", 814=>x"7e00", 815=>x"7200", 816=>x"9700",
---- 817=>x"9200", 818=>x"8c00", 819=>x"8100", 820=>x"9700",
---- 821=>x"9500", 822=>x"9300", 823=>x"8e00", 824=>x"9600",
---- 825=>x"9800", 826=>x"9800", 827=>x"9100", 828=>x"8f00",
---- 829=>x"9500", 830=>x"9b00", 831=>x"9700", 832=>x"8a00",
---- 833=>x"9400", 834=>x"9f00", 835=>x"9f00", 836=>x"8400",
---- 837=>x"9200", 838=>x"a400", 839=>x"a400", 840=>x"7e00",
---- 841=>x"9800", 842=>x"a400", 843=>x"a400", 844=>x"8d00",
---- 845=>x"9600", 846=>x"a500", 847=>x"a800", 848=>x"7200",
---- 849=>x"9300", 850=>x"a400", 851=>x"a900", 852=>x"6e00",
---- 853=>x"9400", 854=>x"a500", 855=>x"ab00", 856=>x"6200",
---- 857=>x"8c00", 858=>x"a300", 859=>x"ad00", 860=>x"5e00",
---- 861=>x"8b00", 862=>x"9e00", 863=>x"aa00", 864=>x"5900",
---- 865=>x"8900", 866=>x"9a00", 867=>x"a400", 868=>x"5300",
---- 869=>x"8500", 870=>x"9a00", 871=>x"a600", 872=>x"4a00",
---- 873=>x"7c00", 874=>x"9c00", 875=>x"a800", 876=>x"4c00",
---- 877=>x"7a00", 878=>x"9a00", 879=>x"aa00", 880=>x"4b00",
---- 881=>x"7b00", 882=>x"9700", 883=>x"a600", 884=>x"4600",
---- 885=>x"7d00", 886=>x"9500", 887=>x"a400", 888=>x"4400",
---- 889=>x"7200", 890=>x"9600", 891=>x"a500", 892=>x"4000",
---- 893=>x"6c00", 894=>x"9400", 895=>x"a400", 896=>x"ca00",
---- 897=>x"6500", 898=>x"8f00", 899=>x"a000", 900=>x"3100",
---- 901=>x"6300", 902=>x"8b00", 903=>x"9d00", 904=>x"3100",
---- 905=>x"5b00", 906=>x"8900", 907=>x"9b00", 908=>x"2c00",
---- 909=>x"5300", 910=>x"8200", 911=>x"9b00", 912=>x"2900",
---- 913=>x"4c00", 914=>x"7d00", 915=>x"9900", 916=>x"2900",
---- 917=>x"4600", 918=>x"7800", 919=>x"9900", 920=>x"2500",
---- 921=>x"4b00", 922=>x"8100", 923=>x"6700", 924=>x"2800",
---- 925=>x"4900", 926=>x"7600", 927=>x"9100", 928=>x"2800",
---- 929=>x"3d00", 930=>x"6900", 931=>x"9800", 932=>x"2900",
---- 933=>x"3200", 934=>x"6800", 935=>x"9d00", 936=>x"2100",
---- 937=>x"3100", 938=>x"6b00", 939=>x"9800", 940=>x"2400",
---- 941=>x"3100", 942=>x"6800", 943=>x"9a00", 944=>x"3300",
---- 945=>x"3600", 946=>x"6800", 947=>x"9700", 948=>x"4000",
---- 949=>x"4300", 950=>x"6600", 951=>x"9200", 952=>x"4e00",
---- 953=>x"5200", 954=>x"6800", 955=>x"8a00", 956=>x"5b00",
---- 957=>x"5c00", 958=>x"7000", 959=>x"8800", 960=>x"6100",
---- 961=>x"6500", 962=>x"7700", 963=>x"8d00", 964=>x"6500",
---- 965=>x"6f00", 966=>x"7f00", 967=>x"9000", 968=>x"6e00",
---- 969=>x"7600", 970=>x"8200", 971=>x"8e00", 972=>x"7300",
---- 973=>x"7300", 974=>x"7b00", 975=>x"8a00", 976=>x"9000",
---- 977=>x"6c00", 978=>x"6b00", 979=>x"8400", 980=>x"5f00",
---- 981=>x"5f00", 982=>x"6800", 983=>x"7f00", 984=>x"5a00",
---- 985=>x"5d00", 986=>x"6700", 987=>x"7b00", 988=>x"5600",
---- 989=>x"5700", 990=>x"5e00", 991=>x"7400", 992=>x"4b00",
---- 993=>x"aa00", 994=>x"5600", 995=>x"6e00", 996=>x"4300",
---- 997=>x"4c00", 998=>x"4f00", 999=>x"6700", 1000=>x"3f00",
---- 1001=>x"3f00", 1002=>x"4400", 1003=>x"6000", 1004=>x"3c00",
---- 1005=>x"3e00", 1006=>x"4100", 1007=>x"6200", 1008=>x"3900",
---- 1009=>x"3a00", 1010=>x"3b00", 1011=>x"6500", 1012=>x"3900",
---- 1013=>x"3700", 1014=>x"3a00", 1015=>x"6100", 1016=>x"3800",
---- 1017=>x"3500", 1018=>x"3800", 1019=>x"5600", 1020=>x"3800",
---- 1021=>x"3100", 1022=>x"cd00", 1023=>x"4d00"),
----
---- 2 => (0=>x"9b00", 1=>x"a000", 2=>x"9d00", 3=>x"9b00", 4=>x"9b00",
---- 5=>x"a200", 6=>x"9c00", 7=>x"9a00", 8=>x"9a00",
---- 9=>x"9f00", 10=>x"9b00", 11=>x"9a00", 12=>x"9b00",
---- 13=>x"9b00", 14=>x"9a00", 15=>x"9700", 16=>x"9b00",
---- 17=>x"9c00", 18=>x"9b00", 19=>x"9a00", 20=>x"9b00",
---- 21=>x"9b00", 22=>x"9d00", 23=>x"9c00", 24=>x"9e00",
---- 25=>x"9d00", 26=>x"9c00", 27=>x"9c00", 28=>x"9d00",
---- 29=>x"9c00", 30=>x"9b00", 31=>x"9a00", 32=>x"9a00",
---- 33=>x"9c00", 34=>x"9c00", 35=>x"9b00", 36=>x"9d00",
---- 37=>x"9f00", 38=>x"9c00", 39=>x"9b00", 40=>x"9f00",
---- 41=>x"9f00", 42=>x"9b00", 43=>x"9c00", 44=>x"9f00",
---- 45=>x"9e00", 46=>x"9c00", 47=>x"9c00", 48=>x"9f00",
---- 49=>x"9c00", 50=>x"9c00", 51=>x"9e00", 52=>x"9e00",
---- 53=>x"9f00", 54=>x"9e00", 55=>x"9c00", 56=>x"9f00",
---- 57=>x"9f00", 58=>x"9f00", 59=>x"9e00", 60=>x"9e00",
---- 61=>x"a000", 62=>x"a000", 63=>x"a100", 64=>x"9f00",
---- 65=>x"a200", 66=>x"a000", 67=>x"a300", 68=>x"a100",
---- 69=>x"a100", 70=>x"a300", 71=>x"a500", 72=>x"a300",
---- 73=>x"a400", 74=>x"a500", 75=>x"a700", 76=>x"a300",
---- 77=>x"5900", 78=>x"a800", 79=>x"a900", 80=>x"a400",
---- 81=>x"a700", 82=>x"a900", 83=>x"a700", 84=>x"a800",
---- 85=>x"a900", 86=>x"a900", 87=>x"a200", 88=>x"ab00",
---- 89=>x"ab00", 90=>x"a700", 91=>x"a000", 92=>x"a900",
---- 93=>x"a500", 94=>x"a000", 95=>x"9c00", 96=>x"ab00",
---- 97=>x"a400", 98=>x"9e00", 99=>x"6500", 100=>x"a900",
---- 101=>x"a200", 102=>x"9c00", 103=>x"9600", 104=>x"a800",
---- 105=>x"a000", 106=>x"9900", 107=>x"6d00", 108=>x"a300",
---- 109=>x"9f00", 110=>x"9500", 111=>x"8f00", 112=>x"9e00",
---- 113=>x"9900", 114=>x"9000", 115=>x"8700", 116=>x"9b00",
---- 117=>x"9300", 118=>x"8b00", 119=>x"7e00", 120=>x"9800",
---- 121=>x"8f00", 122=>x"7f00", 123=>x"7300", 124=>x"6a00",
---- 125=>x"8700", 126=>x"7700", 127=>x"6800", 128=>x"8f00",
---- 129=>x"7d00", 130=>x"6b00", 131=>x"5c00", 132=>x"8800",
---- 133=>x"7400", 134=>x"6100", 135=>x"4f00", 136=>x"7f00",
---- 137=>x"6900", 138=>x"5300", 139=>x"4a00", 140=>x"7100",
---- 141=>x"5600", 142=>x"4a00", 143=>x"4c00", 144=>x"6600",
---- 145=>x"5000", 146=>x"b600", 147=>x"5000", 148=>x"5700",
---- 149=>x"4d00", 150=>x"4d00", 151=>x"ae00", 152=>x"5300",
---- 153=>x"5300", 154=>x"4c00", 155=>x"5100", 156=>x"5400",
---- 157=>x"5700", 158=>x"5100", 159=>x"4f00", 160=>x"5200",
---- 161=>x"5300", 162=>x"5600", 163=>x"5200", 164=>x"5300",
---- 165=>x"5400", 166=>x"5200", 167=>x"5500", 168=>x"5600",
---- 169=>x"5500", 170=>x"5300", 171=>x"5700", 172=>x"5900",
---- 173=>x"5b00", 174=>x"5400", 175=>x"5700", 176=>x"5b00",
---- 177=>x"5900", 178=>x"5300", 179=>x"5600", 180=>x"5800",
---- 181=>x"5700", 182=>x"5600", 183=>x"5700", 184=>x"5900",
---- 185=>x"5700", 186=>x"5800", 187=>x"5600", 188=>x"5900",
---- 189=>x"5900", 190=>x"5600", 191=>x"5500", 192=>x"5b00",
---- 193=>x"5800", 194=>x"5400", 195=>x"5600", 196=>x"5b00",
---- 197=>x"5b00", 198=>x"5500", 199=>x"5600", 200=>x"5c00",
---- 201=>x"5b00", 202=>x"5600", 203=>x"5500", 204=>x"5c00",
---- 205=>x"5a00", 206=>x"5700", 207=>x"5800", 208=>x"5a00",
---- 209=>x"5b00", 210=>x"5700", 211=>x"5a00", 212=>x"5d00",
---- 213=>x"5a00", 214=>x"5900", 215=>x"5b00", 216=>x"5b00",
---- 217=>x"5b00", 218=>x"5900", 219=>x"5700", 220=>x"5c00",
---- 221=>x"5700", 222=>x"5600", 223=>x"5700", 224=>x"5b00",
---- 225=>x"5a00", 226=>x"5700", 227=>x"5500", 228=>x"5600",
---- 229=>x"5500", 230=>x"5400", 231=>x"5300", 232=>x"a300",
---- 233=>x"5900", 234=>x"5400", 235=>x"5400", 236=>x"5b00",
---- 237=>x"5800", 238=>x"5300", 239=>x"5400", 240=>x"5c00",
---- 241=>x"5b00", 242=>x"5800", 243=>x"5400", 244=>x"6000",
---- 245=>x"5c00", 246=>x"5900", 247=>x"5900", 248=>x"6100",
---- 249=>x"5b00", 250=>x"5a00", 251=>x"5600", 252=>x"6100",
---- 253=>x"5f00", 254=>x"5d00", 255=>x"5500", 256=>x"6000",
---- 257=>x"6000", 258=>x"6300", 259=>x"5e00", 260=>x"6100",
---- 261=>x"9d00", 262=>x"6000", 263=>x"5f00", 264=>x"6200",
---- 265=>x"6000", 266=>x"6000", 267=>x"5d00", 268=>x"6100",
---- 269=>x"6000", 270=>x"5f00", 271=>x"5e00", 272=>x"6400",
---- 273=>x"6300", 274=>x"6000", 275=>x"6000", 276=>x"6400",
---- 277=>x"6200", 278=>x"6300", 279=>x"6100", 280=>x"6500",
---- 281=>x"6100", 282=>x"6000", 283=>x"6200", 284=>x"6600",
---- 285=>x"6300", 286=>x"6100", 287=>x"6000", 288=>x"6500",
---- 289=>x"6400", 290=>x"6200", 291=>x"6100", 292=>x"6400",
---- 293=>x"6200", 294=>x"6300", 295=>x"6400", 296=>x"6500",
---- 297=>x"6300", 298=>x"6400", 299=>x"6500", 300=>x"6100",
---- 301=>x"6100", 302=>x"6300", 303=>x"6200", 304=>x"6100",
---- 305=>x"6100", 306=>x"6100", 307=>x"5f00", 308=>x"6300",
---- 309=>x"6500", 310=>x"5e00", 311=>x"6000", 312=>x"9e00",
---- 313=>x"6200", 314=>x"6100", 315=>x"6000", 316=>x"6100",
---- 317=>x"6000", 318=>x"5f00", 319=>x"6300", 320=>x"5f00",
---- 321=>x"6000", 322=>x"6000", 323=>x"6500", 324=>x"5e00",
---- 325=>x"6000", 326=>x"5f00", 327=>x"6100", 328=>x"5d00",
---- 329=>x"6000", 330=>x"6100", 331=>x"6000", 332=>x"5d00",
---- 333=>x"5c00", 334=>x"5f00", 335=>x"6100", 336=>x"5f00",
---- 337=>x"6000", 338=>x"6200", 339=>x"6400", 340=>x"6100",
---- 341=>x"6300", 342=>x"6500", 343=>x"6900", 344=>x"6200",
---- 345=>x"6200", 346=>x"6700", 347=>x"6a00", 348=>x"6300",
---- 349=>x"6300", 350=>x"6700", 351=>x"6900", 352=>x"6600",
---- 353=>x"5f00", 354=>x"6400", 355=>x"6700", 356=>x"6700",
---- 357=>x"6500", 358=>x"6700", 359=>x"6900", 360=>x"6300",
---- 361=>x"6600", 362=>x"6a00", 363=>x"6b00", 364=>x"6400",
---- 365=>x"6400", 366=>x"6900", 367=>x"6e00", 368=>x"6200",
---- 369=>x"6900", 370=>x"6a00", 371=>x"6c00", 372=>x"5f00",
---- 373=>x"6800", 374=>x"6b00", 375=>x"6b00", 376=>x"6100",
---- 377=>x"6500", 378=>x"6a00", 379=>x"6c00", 380=>x"6300",
---- 381=>x"6300", 382=>x"6700", 383=>x"6b00", 384=>x"6500",
---- 385=>x"6400", 386=>x"9b00", 387=>x"6900", 388=>x"6200",
---- 389=>x"6200", 390=>x"6500", 391=>x"6700", 392=>x"6400",
---- 393=>x"6500", 394=>x"6700", 395=>x"6800", 396=>x"6500",
---- 397=>x"6600", 398=>x"6500", 399=>x"6600", 400=>x"6600",
---- 401=>x"6400", 402=>x"6600", 403=>x"6600", 404=>x"6400",
---- 405=>x"6100", 406=>x"6600", 407=>x"6500", 408=>x"6200",
---- 409=>x"6200", 410=>x"6200", 411=>x"6200", 412=>x"6500",
---- 413=>x"6300", 414=>x"6100", 415=>x"5f00", 416=>x"6200",
---- 417=>x"6500", 418=>x"6200", 419=>x"5f00", 420=>x"6500",
---- 421=>x"6300", 422=>x"5f00", 423=>x"5e00", 424=>x"6500",
---- 425=>x"6100", 426=>x"6100", 427=>x"5b00", 428=>x"6500",
---- 429=>x"6400", 430=>x"5f00", 431=>x"5a00", 432=>x"6200",
---- 433=>x"6200", 434=>x"5f00", 435=>x"5900", 436=>x"6300",
---- 437=>x"6300", 438=>x"5e00", 439=>x"5900", 440=>x"6200",
---- 441=>x"6200", 442=>x"5f00", 443=>x"5b00", 444=>x"6500",
---- 445=>x"6500", 446=>x"6200", 447=>x"5c00", 448=>x"6200",
---- 449=>x"6400", 450=>x"6200", 451=>x"5d00", 452=>x"6300",
---- 453=>x"6000", 454=>x"5f00", 455=>x"5e00", 456=>x"6400",
---- 457=>x"6200", 458=>x"6000", 459=>x"5e00", 460=>x"6200",
---- 461=>x"6300", 462=>x"5f00", 463=>x"5b00", 464=>x"6200",
---- 465=>x"6000", 466=>x"5c00", 467=>x"5c00", 468=>x"5e00",
---- 469=>x"5c00", 470=>x"5d00", 471=>x"5b00", 472=>x"6100",
---- 473=>x"6000", 474=>x"5c00", 475=>x"5c00", 476=>x"6200",
---- 477=>x"6300", 478=>x"6100", 479=>x"5b00", 480=>x"6000",
---- 481=>x"6200", 482=>x"6200", 483=>x"5a00", 484=>x"5e00",
---- 485=>x"6100", 486=>x"5f00", 487=>x"5a00", 488=>x"6100",
---- 489=>x"6100", 490=>x"5f00", 491=>x"5e00", 492=>x"6500",
---- 493=>x"6300", 494=>x"5f00", 495=>x"5d00", 496=>x"6200",
---- 497=>x"6400", 498=>x"6000", 499=>x"5d00", 500=>x"6500",
---- 501=>x"9d00", 502=>x"6100", 503=>x"5e00", 504=>x"6500",
---- 505=>x"6300", 506=>x"9c00", 507=>x"5b00", 508=>x"6400",
---- 509=>x"6200", 510=>x"5e00", 511=>x"5700", 512=>x"6500",
---- 513=>x"5f00", 514=>x"5c00", 515=>x"5500", 516=>x"6300",
---- 517=>x"6000", 518=>x"5c00", 519=>x"5800", 520=>x"5d00",
---- 521=>x"5f00", 522=>x"5900", 523=>x"5500", 524=>x"5d00",
---- 525=>x"5b00", 526=>x"5500", 527=>x"4e00", 528=>x"5a00",
---- 529=>x"5800", 530=>x"5300", 531=>x"5300", 532=>x"5a00",
---- 533=>x"5500", 534=>x"5200", 535=>x"4f00", 536=>x"5a00",
---- 537=>x"5700", 538=>x"5600", 539=>x"4f00", 540=>x"5a00",
---- 541=>x"5a00", 542=>x"5200", 543=>x"4d00", 544=>x"5900",
---- 545=>x"5a00", 546=>x"5300", 547=>x"4e00", 548=>x"5b00",
---- 549=>x"5900", 550=>x"5600", 551=>x"4b00", 552=>x"5b00",
---- 553=>x"5600", 554=>x"5300", 555=>x"4e00", 556=>x"5800",
---- 557=>x"5600", 558=>x"4f00", 559=>x"4e00", 560=>x"5500",
---- 561=>x"a900", 562=>x"5200", 563=>x"4a00", 564=>x"5400",
---- 565=>x"5300", 566=>x"5100", 567=>x"4b00", 568=>x"5300",
---- 569=>x"5200", 570=>x"4a00", 571=>x"4300", 572=>x"5100",
---- 573=>x"5200", 574=>x"4900", 575=>x"4200", 576=>x"5100",
---- 577=>x"4f00", 578=>x"4700", 579=>x"4100", 580=>x"4d00",
---- 581=>x"4c00", 582=>x"4600", 583=>x"3e00", 584=>x"4c00",
---- 585=>x"4b00", 586=>x"4600", 587=>x"3f00", 588=>x"4c00",
---- 589=>x"4900", 590=>x"4600", 591=>x"3f00", 592=>x"4b00",
---- 593=>x"4700", 594=>x"4300", 595=>x"3d00", 596=>x"4900",
---- 597=>x"4a00", 598=>x"4300", 599=>x"4000", 600=>x"4600",
---- 601=>x"4500", 602=>x"4100", 603=>x"3c00", 604=>x"4300",
---- 605=>x"4400", 606=>x"4000", 607=>x"3900", 608=>x"4500",
---- 609=>x"4400", 610=>x"c100", 611=>x"3900", 612=>x"4600",
---- 613=>x"4200", 614=>x"3f00", 615=>x"3500", 616=>x"4100",
---- 617=>x"4100", 618=>x"3e00", 619=>x"3500", 620=>x"4300",
---- 621=>x"3f00", 622=>x"3c00", 623=>x"3700", 624=>x"4400",
---- 625=>x"3f00", 626=>x"3500", 627=>x"3300", 628=>x"4300",
---- 629=>x"3e00", 630=>x"3600", 631=>x"3100", 632=>x"4000",
---- 633=>x"3900", 634=>x"3700", 635=>x"3100", 636=>x"4200",
---- 637=>x"3e00", 638=>x"3a00", 639=>x"3000", 640=>x"4500",
---- 641=>x"4100", 642=>x"3e00", 643=>x"3300", 644=>x"4200",
---- 645=>x"4000", 646=>x"3e00", 647=>x"3900", 648=>x"4400",
---- 649=>x"4000", 650=>x"4000", 651=>x"c300", 652=>x"4500",
---- 653=>x"4500", 654=>x"4500", 655=>x"4300", 656=>x"4300",
---- 657=>x"4100", 658=>x"4600", 659=>x"4700", 660=>x"4400",
---- 661=>x"4200", 662=>x"4800", 663=>x"4b00", 664=>x"4600",
---- 665=>x"4700", 666=>x"4300", 667=>x"4a00", 668=>x"4900",
---- 669=>x"4100", 670=>x"3c00", 671=>x"4400", 672=>x"4600",
---- 673=>x"3d00", 674=>x"3a00", 675=>x"4400", 676=>x"4000",
---- 677=>x"3d00", 678=>x"3c00", 679=>x"4500", 680=>x"4100",
---- 681=>x"4100", 682=>x"3f00", 683=>x"4800", 684=>x"4100",
---- 685=>x"3e00", 686=>x"4200", 687=>x"4b00", 688=>x"4000",
---- 689=>x"4000", 690=>x"4500", 691=>x"4300", 692=>x"4300",
---- 693=>x"3f00", 694=>x"3f00", 695=>x"4800", 696=>x"4200",
---- 697=>x"3c00", 698=>x"3d00", 699=>x"b800", 700=>x"3e00",
---- 701=>x"3d00", 702=>x"4100", 703=>x"4a00", 704=>x"3f00",
---- 705=>x"4000", 706=>x"4000", 707=>x"5000", 708=>x"3c00",
---- 709=>x"3d00", 710=>x"4600", 711=>x"5700", 712=>x"3d00",
---- 713=>x"3b00", 714=>x"4900", 715=>x"5100", 716=>x"3b00",
---- 717=>x"3700", 718=>x"4600", 719=>x"5600", 720=>x"3700",
---- 721=>x"3800", 722=>x"4600", 723=>x"ac00", 724=>x"3600",
---- 725=>x"3800", 726=>x"4700", 727=>x"5500", 728=>x"3500",
---- 729=>x"3700", 730=>x"4800", 731=>x"5c00", 732=>x"3300",
---- 733=>x"3900", 734=>x"5100", 735=>x"6000", 736=>x"2e00",
---- 737=>x"3e00", 738=>x"6200", 739=>x"6400", 740=>x"2e00",
---- 741=>x"4500", 742=>x"6400", 743=>x"6900", 744=>x"3400",
---- 745=>x"4f00", 746=>x"6500", 747=>x"6600", 748=>x"3500",
---- 749=>x"4e00", 750=>x"6500", 751=>x"6800", 752=>x"3500",
---- 753=>x"5300", 754=>x"6500", 755=>x"6d00", 756=>x"3900",
---- 757=>x"5200", 758=>x"5900", 759=>x"6100", 760=>x"3700",
---- 761=>x"4600", 762=>x"5600", 763=>x"5e00", 764=>x"3100",
---- 765=>x"3c00", 766=>x"5100", 767=>x"5e00", 768=>x"3300",
---- 769=>x"3500", 770=>x"4a00", 771=>x"5e00", 772=>x"2b00",
---- 773=>x"3800", 774=>x"4500", 775=>x"5c00", 776=>x"2700",
---- 777=>x"3400", 778=>x"4500", 779=>x"5700", 780=>x"2a00",
---- 781=>x"3300", 782=>x"4500", 783=>x"5000", 784=>x"2500",
---- 785=>x"3200", 786=>x"3f00", 787=>x"4900", 788=>x"2800",
---- 789=>x"2f00", 790=>x"3c00", 791=>x"4700", 792=>x"2f00",
---- 793=>x"3500", 794=>x"4300", 795=>x"4200", 796=>x"3300",
---- 797=>x"3d00", 798=>x"3e00", 799=>x"3900", 800=>x"3b00",
---- 801=>x"4600", 802=>x"3e00", 803=>x"3700", 804=>x"4700",
---- 805=>x"4d00", 806=>x"4500", 807=>x"3800", 808=>x"5700",
---- 809=>x"5600", 810=>x"b100", 811=>x"4200", 812=>x"6400",
---- 813=>x"5f00", 814=>x"5500", 815=>x"4800", 816=>x"7300",
---- 817=>x"6900", 818=>x"5800", 819=>x"4800", 820=>x"8100",
---- 821=>x"7500", 822=>x"6100", 823=>x"4b00", 824=>x"8500",
---- 825=>x"8300", 826=>x"7200", 827=>x"5700", 828=>x"9200",
---- 829=>x"9300", 830=>x"7e00", 831=>x"6200", 832=>x"a100",
---- 833=>x"9900", 834=>x"8500", 835=>x"6c00", 836=>x"a400",
---- 837=>x"9800", 838=>x"8a00", 839=>x"7800", 840=>x"a700",
---- 841=>x"9e00", 842=>x"8e00", 843=>x"7d00", 844=>x"ab00",
---- 845=>x"a300", 846=>x"9300", 847=>x"8500", 848=>x"ab00",
---- 849=>x"a400", 850=>x"9a00", 851=>x"8600", 852=>x"aa00",
---- 853=>x"a900", 854=>x"9c00", 855=>x"8c00", 856=>x"af00",
---- 857=>x"a900", 858=>x"a000", 859=>x"8900", 860=>x"ad00",
---- 861=>x"a800", 862=>x"9900", 863=>x"8400", 864=>x"aa00",
---- 865=>x"aa00", 866=>x"9c00", 867=>x"8500", 868=>x"ad00",
---- 869=>x"ac00", 870=>x"a000", 871=>x"8b00", 872=>x"ae00",
---- 873=>x"aa00", 874=>x"9e00", 875=>x"8c00", 876=>x"b100",
---- 877=>x"af00", 878=>x"a000", 879=>x"8d00", 880=>x"4f00",
---- 881=>x"ab00", 882=>x"a000", 883=>x"8c00", 884=>x"ac00",
---- 885=>x"aa00", 886=>x"a200", 887=>x"8e00", 888=>x"ac00",
---- 889=>x"ac00", 890=>x"a200", 891=>x"9100", 892=>x"ad00",
---- 893=>x"ad00", 894=>x"a700", 895=>x"9700", 896=>x"ac00",
---- 897=>x"ac00", 898=>x"a900", 899=>x"9800", 900=>x"a800",
---- 901=>x"ad00", 902=>x"a500", 903=>x"9700", 904=>x"a800",
---- 905=>x"ab00", 906=>x"a400", 907=>x"9900", 908=>x"aa00",
---- 909=>x"ab00", 910=>x"a700", 911=>x"9700", 912=>x"a400",
---- 913=>x"ab00", 914=>x"a700", 915=>x"9a00", 916=>x"a200",
---- 917=>x"a600", 918=>x"a300", 919=>x"9900", 920=>x"9f00",
---- 921=>x"a400", 922=>x"a300", 923=>x"9700", 924=>x"a200",
---- 925=>x"ad00", 926=>x"ac00", 927=>x"a100", 928=>x"ad00",
---- 929=>x"af00", 930=>x"af00", 931=>x"a500", 932=>x"a800",
---- 933=>x"b000", 934=>x"b000", 935=>x"5700", 936=>x"a700",
---- 937=>x"af00", 938=>x"af00", 939=>x"a900", 940=>x"a600",
---- 941=>x"af00", 942=>x"b300", 943=>x"aa00", 944=>x"a700",
---- 945=>x"b200", 946=>x"b500", 947=>x"ac00", 948=>x"aa00",
---- 949=>x"b200", 950=>x"b500", 951=>x"b300", 952=>x"a500",
---- 953=>x"b400", 954=>x"b900", 955=>x"b600", 956=>x"a400",
---- 957=>x"b200", 958=>x"b800", 959=>x"b400", 960=>x"a500",
---- 961=>x"b000", 962=>x"b700", 963=>x"b600", 964=>x"a600",
---- 965=>x"b000", 966=>x"b500", 967=>x"b700", 968=>x"a800",
---- 969=>x"b200", 970=>x"b400", 971=>x"b000", 972=>x"a300",
---- 973=>x"ad00", 974=>x"b100", 975=>x"af00", 976=>x"9c00",
---- 977=>x"aa00", 978=>x"b000", 979=>x"b000", 980=>x"9800",
---- 981=>x"a800", 982=>x"b200", 983=>x"b400", 984=>x"9400",
---- 985=>x"aa00", 986=>x"b000", 987=>x"b000", 988=>x"8f00",
---- 989=>x"a400", 990=>x"ac00", 991=>x"ae00", 992=>x"8900",
---- 993=>x"a300", 994=>x"ad00", 995=>x"b200", 996=>x"8b00",
---- 997=>x"a600", 998=>x"b600", 999=>x"bc00", 1000=>x"8d00",
---- 1001=>x"b300", 1002=>x"c500", 1003=>x"c900", 1004=>x"9200",
---- 1005=>x"c100", 1006=>x"ca00", 1007=>x"cc00", 1008=>x"9f00",
---- 1009=>x"c600", 1010=>x"c700", 1011=>x"cc00", 1012=>x"a300",
---- 1013=>x"c600", 1014=>x"c500", 1015=>x"ca00", 1016=>x"9e00",
---- 1017=>x"c600", 1018=>x"c500", 1019=>x"c700", 1020=>x"9600",
---- 1021=>x"c400", 1022=>x"c500", 1023=>x"3800"),
----
---- 3 => (0=>x"9c00", 1=>x"9a00", 2=>x"9a00", 3=>x"9b00", 4=>x"9c00",
---- 5=>x"9900", 6=>x"9a00", 7=>x"9900", 8=>x"9c00",
---- 9=>x"9a00", 10=>x"9a00", 11=>x"9a00", 12=>x"9a00",
---- 13=>x"9a00", 14=>x"9800", 15=>x"9a00", 16=>x"9b00",
---- 17=>x"9a00", 18=>x"9800", 19=>x"9a00", 20=>x"9800",
---- 21=>x"9900", 22=>x"9c00", 23=>x"9a00", 24=>x"9a00",
---- 25=>x"9900", 26=>x"6400", 27=>x"6400", 28=>x"9a00",
---- 29=>x"9a00", 30=>x"9b00", 31=>x"9c00", 32=>x"9900",
---- 33=>x"9800", 34=>x"9a00", 35=>x"a100", 36=>x"9b00",
---- 37=>x"9900", 38=>x"9d00", 39=>x"a100", 40=>x"9b00",
---- 41=>x"9b00", 42=>x"9e00", 43=>x"a000", 44=>x"9800",
---- 45=>x"9b00", 46=>x"9c00", 47=>x"a200", 48=>x"9d00",
---- 49=>x"9e00", 50=>x"a100", 51=>x"a400", 52=>x"9d00",
---- 53=>x"a100", 54=>x"a300", 55=>x"a600", 56=>x"9e00",
---- 57=>x"a200", 58=>x"a700", 59=>x"a800", 60=>x"a300",
---- 61=>x"a700", 62=>x"a700", 63=>x"a800", 64=>x"a700",
---- 65=>x"a800", 66=>x"a800", 67=>x"aa00", 68=>x"a800",
---- 69=>x"a700", 70=>x"a800", 71=>x"a800", 72=>x"a800",
---- 73=>x"a800", 74=>x"a800", 75=>x"a900", 76=>x"a700",
---- 77=>x"a800", 78=>x"a700", 79=>x"a400", 80=>x"a500",
---- 81=>x"a400", 82=>x"5e00", 83=>x"a200", 84=>x"a200",
---- 85=>x"a200", 86=>x"9e00", 87=>x"a100", 88=>x"9c00",
---- 89=>x"9e00", 90=>x"9a00", 91=>x"9d00", 92=>x"9a00",
---- 93=>x"9a00", 94=>x"9900", 95=>x"9700", 96=>x"9700",
---- 97=>x"9500", 98=>x"9400", 99=>x"9500", 100=>x"9200",
---- 101=>x"6e00", 102=>x"8e00", 103=>x"9100", 104=>x"8c00",
---- 105=>x"8c00", 106=>x"8d00", 107=>x"8a00", 108=>x"8700",
---- 109=>x"8200", 110=>x"8700", 111=>x"8a00", 112=>x"8100",
---- 113=>x"7e00", 114=>x"8000", 115=>x"8a00", 116=>x"7900",
---- 117=>x"7800", 118=>x"8000", 119=>x"8f00", 120=>x"6d00",
---- 121=>x"6f00", 122=>x"8000", 123=>x"9000", 124=>x"6100",
---- 125=>x"7000", 126=>x"8100", 127=>x"8d00", 128=>x"5a00",
---- 129=>x"7000", 130=>x"8000", 131=>x"8e00", 132=>x"5900",
---- 133=>x"7000", 134=>x"8100", 135=>x"8e00", 136=>x"5700",
---- 137=>x"6f00", 138=>x"8200", 139=>x"8e00", 140=>x"5a00",
---- 141=>x"7200", 142=>x"8000", 143=>x"8a00", 144=>x"6000",
---- 145=>x"6e00", 146=>x"8000", 147=>x"8c00", 148=>x"6000",
---- 149=>x"7200", 150=>x"8000", 151=>x"8c00", 152=>x"5f00",
---- 153=>x"7400", 154=>x"8100", 155=>x"8b00", 156=>x"5e00",
---- 157=>x"7100", 158=>x"8200", 159=>x"8c00", 160=>x"6000",
---- 161=>x"7400", 162=>x"8200", 163=>x"8e00", 164=>x"5f00",
---- 165=>x"7300", 166=>x"8400", 167=>x"8e00", 168=>x"6000",
---- 169=>x"7200", 170=>x"7f00", 171=>x"8d00", 172=>x"5f00",
---- 173=>x"7000", 174=>x"8000", 175=>x"8d00", 176=>x"6300",
---- 177=>x"8d00", 178=>x"8200", 179=>x"7200", 180=>x"9f00",
---- 181=>x"7000", 182=>x"7f00", 183=>x"8e00", 184=>x"5d00",
---- 185=>x"7000", 186=>x"7e00", 187=>x"8c00", 188=>x"5d00",
---- 189=>x"6e00", 190=>x"8000", 191=>x"8c00", 192=>x"5d00",
---- 193=>x"6f00", 194=>x"8200", 195=>x"8c00", 196=>x"6000",
---- 197=>x"6e00", 198=>x"7e00", 199=>x"8700", 200=>x"5e00",
---- 201=>x"6c00", 202=>x"7b00", 203=>x"8900", 204=>x"5f00",
---- 205=>x"6d00", 206=>x"7d00", 207=>x"8c00", 208=>x"6100",
---- 209=>x"6e00", 210=>x"8000", 211=>x"8b00", 212=>x"6300",
---- 213=>x"7100", 214=>x"8000", 215=>x"8a00", 216=>x"5f00",
---- 217=>x"7100", 218=>x"7f00", 219=>x"8a00", 220=>x"5c00",
---- 221=>x"6f00", 222=>x"7d00", 223=>x"8c00", 224=>x"5c00",
---- 225=>x"6a00", 226=>x"7d00", 227=>x"8d00", 228=>x"5c00",
---- 229=>x"6b00", 230=>x"8000", 231=>x"8c00", 232=>x"a600",
---- 233=>x"6a00", 234=>x"7a00", 235=>x"8800", 236=>x"5600",
---- 237=>x"6900", 238=>x"7b00", 239=>x"8800", 240=>x"5b00",
---- 241=>x"6c00", 242=>x"7d00", 243=>x"8700", 244=>x"5b00",
---- 245=>x"6d00", 246=>x"7c00", 247=>x"8600", 248=>x"5b00",
---- 249=>x"6c00", 250=>x"7800", 251=>x"7700", 252=>x"5e00",
---- 253=>x"6a00", 254=>x"7900", 255=>x"8800", 256=>x"6000",
---- 257=>x"6b00", 258=>x"7e00", 259=>x"8500", 260=>x"5f00",
---- 261=>x"6d00", 262=>x"7900", 263=>x"8a00", 264=>x"5f00",
---- 265=>x"6c00", 266=>x"7b00", 267=>x"8a00", 268=>x"6100",
---- 269=>x"6900", 270=>x"7b00", 271=>x"8900", 272=>x"6100",
---- 273=>x"6d00", 274=>x"7c00", 275=>x"8900", 276=>x"6600",
---- 277=>x"6e00", 278=>x"7e00", 279=>x"8a00", 280=>x"6900",
---- 281=>x"7100", 282=>x"7f00", 283=>x"8b00", 284=>x"6900",
---- 285=>x"7100", 286=>x"7e00", 287=>x"8a00", 288=>x"6600",
---- 289=>x"7200", 290=>x"7d00", 291=>x"8a00", 292=>x"6600",
---- 293=>x"7200", 294=>x"7e00", 295=>x"8900", 296=>x"6800",
---- 297=>x"7200", 298=>x"7e00", 299=>x"8800", 300=>x"6700",
---- 301=>x"6f00", 302=>x"7a00", 303=>x"8800", 304=>x"6300",
---- 305=>x"6e00", 306=>x"7900", 307=>x"8a00", 308=>x"6400",
---- 309=>x"6c00", 310=>x"7b00", 311=>x"8900", 312=>x"6700",
---- 313=>x"6f00", 314=>x"7c00", 315=>x"8900", 316=>x"6400",
---- 317=>x"6c00", 318=>x"7e00", 319=>x"8b00", 320=>x"6200",
---- 321=>x"6e00", 322=>x"7f00", 323=>x"8f00", 324=>x"6400",
---- 325=>x"7200", 326=>x"7f00", 327=>x"8c00", 328=>x"6400",
---- 329=>x"7100", 330=>x"7f00", 331=>x"8c00", 332=>x"6800",
---- 333=>x"7300", 334=>x"8200", 335=>x"8b00", 336=>x"6800",
---- 337=>x"7600", 338=>x"8100", 339=>x"8d00", 340=>x"6900",
---- 341=>x"7600", 342=>x"7f00", 343=>x"8b00", 344=>x"6b00",
---- 345=>x"7400", 346=>x"8100", 347=>x"8b00", 348=>x"9400",
---- 349=>x"7400", 350=>x"7f00", 351=>x"8d00", 352=>x"6d00",
---- 353=>x"7500", 354=>x"8400", 355=>x"8d00", 356=>x"7100",
---- 357=>x"7a00", 358=>x"8400", 359=>x"8e00", 360=>x"7000",
---- 361=>x"7800", 362=>x"8500", 363=>x"9100", 364=>x"6f00",
---- 365=>x"7600", 366=>x"8500", 367=>x"9000", 368=>x"7000",
---- 369=>x"7a00", 370=>x"8100", 371=>x"8d00", 372=>x"7100",
---- 373=>x"7a00", 374=>x"8700", 375=>x"8c00", 376=>x"6f00",
---- 377=>x"7800", 378=>x"8400", 379=>x"8e00", 380=>x"6c00",
---- 381=>x"7900", 382=>x"8300", 383=>x"8e00", 384=>x"6c00",
---- 385=>x"7800", 386=>x"8400", 387=>x"9000", 388=>x"6e00",
---- 389=>x"7600", 390=>x"8200", 391=>x"8f00", 392=>x"6d00",
---- 393=>x"7400", 394=>x"7f00", 395=>x"8d00", 396=>x"6a00",
---- 397=>x"7700", 398=>x"8300", 399=>x"8c00", 400=>x"6700",
---- 401=>x"7200", 402=>x"7d00", 403=>x"8b00", 404=>x"6600",
---- 405=>x"7400", 406=>x"7f00", 407=>x"8a00", 408=>x"6500",
---- 409=>x"7200", 410=>x"7e00", 411=>x"8800", 412=>x"9d00",
---- 413=>x"6d00", 414=>x"7c00", 415=>x"8900", 416=>x"6200",
---- 417=>x"6c00", 418=>x"7800", 419=>x"8900", 420=>x"5e00",
---- 421=>x"6800", 422=>x"7c00", 423=>x"8800", 424=>x"5d00",
---- 425=>x"6900", 426=>x"7900", 427=>x"8700", 428=>x"5a00",
---- 429=>x"6700", 430=>x"7700", 431=>x"8600", 432=>x"5c00",
---- 433=>x"6800", 434=>x"7900", 435=>x"8600", 436=>x"5900",
---- 437=>x"6400", 438=>x"7800", 439=>x"8500", 440=>x"5a00",
---- 441=>x"6400", 442=>x"7700", 443=>x"8700", 444=>x"5c00",
---- 445=>x"6900", 446=>x"7800", 447=>x"8500", 448=>x"5a00",
---- 449=>x"6600", 450=>x"7700", 451=>x"8700", 452=>x"5c00",
---- 453=>x"6400", 454=>x"7500", 455=>x"8800", 456=>x"5a00",
---- 457=>x"6600", 458=>x"7700", 459=>x"8800", 460=>x"5e00",
---- 461=>x"6800", 462=>x"7600", 463=>x"8600", 464=>x"5f00",
---- 465=>x"6500", 466=>x"7300", 467=>x"8200", 468=>x"5500",
---- 469=>x"6200", 470=>x"8900", 471=>x"8300", 472=>x"5800",
---- 473=>x"6500", 474=>x"7800", 475=>x"8600", 476=>x"5b00",
---- 477=>x"6400", 478=>x"7600", 479=>x"8500", 480=>x"5800",
---- 481=>x"6400", 482=>x"7400", 483=>x"8600", 484=>x"5900",
---- 485=>x"6400", 486=>x"7300", 487=>x"8800", 488=>x"5800",
---- 489=>x"6300", 490=>x"7200", 491=>x"8700", 492=>x"5c00",
---- 493=>x"6100", 494=>x"7400", 495=>x"8500", 496=>x"5900",
---- 497=>x"6000", 498=>x"7300", 499=>x"8500", 500=>x"5900",
---- 501=>x"6000", 502=>x"7200", 503=>x"8500", 504=>x"5900",
---- 505=>x"6000", 506=>x"7100", 507=>x"8200", 508=>x"5600",
---- 509=>x"5f00", 510=>x"7300", 511=>x"8300", 512=>x"5500",
---- 513=>x"5f00", 514=>x"7300", 515=>x"8400", 516=>x"5200",
---- 517=>x"5b00", 518=>x"7400", 519=>x"8500", 520=>x"5200",
---- 521=>x"5700", 522=>x"6f00", 523=>x"8200", 524=>x"4c00",
---- 525=>x"5500", 526=>x"6a00", 527=>x"7f00", 528=>x"4a00",
---- 529=>x"5200", 530=>x"6900", 531=>x"8100", 532=>x"4800",
---- 533=>x"ac00", 534=>x"6d00", 535=>x"8300", 536=>x"4700",
---- 537=>x"5200", 538=>x"6c00", 539=>x"8100", 540=>x"4600",
---- 541=>x"4f00", 542=>x"6800", 543=>x"8000", 544=>x"4600",
---- 545=>x"5200", 546=>x"6800", 547=>x"7e00", 548=>x"4800",
---- 549=>x"4f00", 550=>x"6900", 551=>x"8100", 552=>x"4700",
---- 553=>x"4d00", 554=>x"6900", 555=>x"8000", 556=>x"4600",
---- 557=>x"4d00", 558=>x"6600", 559=>x"7f00", 560=>x"4600",
---- 561=>x"4a00", 562=>x"6400", 563=>x"7e00", 564=>x"4100",
---- 565=>x"4900", 566=>x"6200", 567=>x"7b00", 568=>x"3800",
---- 569=>x"4000", 570=>x"6000", 571=>x"7d00", 572=>x"3c00",
---- 573=>x"4100", 574=>x"5a00", 575=>x"7b00", 576=>x"3c00",
---- 577=>x"4600", 578=>x"5b00", 579=>x"7a00", 580=>x"3b00",
---- 581=>x"4300", 582=>x"5900", 583=>x"7700", 584=>x"3900",
---- 585=>x"4200", 586=>x"6000", 587=>x"7900", 588=>x"3800",
---- 589=>x"4200", 590=>x"5f00", 591=>x"7900", 592=>x"3a00",
---- 593=>x"3e00", 594=>x"5900", 595=>x"7900", 596=>x"3900",
---- 597=>x"3f00", 598=>x"5900", 599=>x"7900", 600=>x"3700",
---- 601=>x"4000", 602=>x"5800", 603=>x"7800", 604=>x"3500",
---- 605=>x"4100", 606=>x"5400", 607=>x"7600", 608=>x"3400",
---- 609=>x"3a00", 610=>x"5700", 611=>x"7700", 612=>x"3100",
---- 613=>x"3d00", 614=>x"5c00", 615=>x"7800", 616=>x"3200",
---- 617=>x"3c00", 618=>x"5800", 619=>x"7600", 620=>x"2f00",
---- 621=>x"3600", 622=>x"5500", 623=>x"7900", 624=>x"2c00",
---- 625=>x"3100", 626=>x"5400", 627=>x"7600", 628=>x"2c00",
---- 629=>x"3000", 630=>x"5400", 631=>x"7400", 632=>x"2a00",
---- 633=>x"2f00", 634=>x"4f00", 635=>x"7300", 636=>x"2a00",
---- 637=>x"d000", 638=>x"5200", 639=>x"7600", 640=>x"2900",
---- 641=>x"3800", 642=>x"5900", 643=>x"7500", 644=>x"3000",
---- 645=>x"3e00", 646=>x"5b00", 647=>x"7800", 648=>x"3700",
---- 649=>x"4600", 650=>x"6700", 651=>x"7e00", 652=>x"4000",
---- 653=>x"4f00", 654=>x"9300", 655=>x"8200", 656=>x"4a00",
---- 657=>x"5600", 658=>x"7300", 659=>x"8600", 660=>x"4f00",
---- 661=>x"5a00", 662=>x"7600", 663=>x"8900", 664=>x"5500",
---- 665=>x"6200", 666=>x"7800", 667=>x"8b00", 668=>x"5700",
---- 669=>x"6600", 670=>x"7800", 671=>x"8b00", 672=>x"5400",
---- 673=>x"6600", 674=>x"7f00", 675=>x"8c00", 676=>x"5500",
---- 677=>x"6800", 678=>x"7e00", 679=>x"8c00", 680=>x"5100",
---- 681=>x"6400", 682=>x"7b00", 683=>x"8900", 684=>x"5000",
---- 685=>x"6000", 686=>x"7700", 687=>x"8600", 688=>x"4f00",
---- 689=>x"5f00", 690=>x"7700", 691=>x"8900", 692=>x"5100",
---- 693=>x"5e00", 694=>x"7a00", 695=>x"8900", 696=>x"4e00",
---- 697=>x"5a00", 698=>x"7800", 699=>x"8b00", 700=>x"5000",
---- 701=>x"6100", 702=>x"7700", 703=>x"8d00", 704=>x"5600",
---- 705=>x"6600", 706=>x"7a00", 707=>x"8d00", 708=>x"5b00",
---- 709=>x"6700", 710=>x"7e00", 711=>x"8d00", 712=>x"5b00",
---- 713=>x"6600", 714=>x"7b00", 715=>x"8c00", 716=>x"5b00",
---- 717=>x"6400", 718=>x"7800", 719=>x"8a00", 720=>x"5b00",
---- 721=>x"5f00", 722=>x"7600", 723=>x"8a00", 724=>x"5d00",
---- 725=>x"5e00", 726=>x"7200", 727=>x"8900", 728=>x"5800",
---- 729=>x"5700", 730=>x"7200", 731=>x"8600", 732=>x"5a00",
---- 733=>x"5800", 734=>x"6e00", 735=>x"8400", 736=>x"6100",
---- 737=>x"6300", 738=>x"7300", 739=>x"8100", 740=>x"6500",
---- 741=>x"6700", 742=>x"7700", 743=>x"8400", 744=>x"6600",
---- 745=>x"6700", 746=>x"7800", 747=>x"8300", 748=>x"6500",
---- 749=>x"6600", 750=>x"7a00", 751=>x"8400", 752=>x"6700",
---- 753=>x"6400", 754=>x"7800", 755=>x"8500", 756=>x"5f00",
---- 757=>x"6500", 758=>x"7700", 759=>x"8500", 760=>x"6200",
---- 761=>x"6900", 762=>x"7c00", 763=>x"8800", 764=>x"6500",
---- 765=>x"7000", 766=>x"8100", 767=>x"8400", 768=>x"9c00",
---- 769=>x"6a00", 770=>x"7a00", 771=>x"8300", 772=>x"6000",
---- 773=>x"5c00", 774=>x"7100", 775=>x"8300", 776=>x"5d00",
---- 777=>x"5900", 778=>x"6800", 779=>x"7e00", 780=>x"5200",
---- 781=>x"4d00", 782=>x"6400", 783=>x"7f00", 784=>x"4d00",
---- 785=>x"4a00", 786=>x"9e00", 787=>x"8000", 788=>x"4800",
---- 789=>x"4700", 790=>x"a300", 791=>x"7700", 792=>x"3b00",
---- 793=>x"3f00", 794=>x"5100", 795=>x"6b00", 796=>x"3600",
---- 797=>x"3400", 798=>x"4300", 799=>x"5f00", 800=>x"3500",
---- 801=>x"cd00", 802=>x"4000", 803=>x"5600", 804=>x"3500",
---- 805=>x"3100", 806=>x"3e00", 807=>x"5700", 808=>x"3200",
---- 809=>x"2d00", 810=>x"3c00", 811=>x"5700", 812=>x"3200",
---- 813=>x"2b00", 814=>x"3a00", 815=>x"5500", 816=>x"3800",
---- 817=>x"2b00", 818=>x"3500", 819=>x"5500", 820=>x"3c00",
---- 821=>x"2b00", 822=>x"3400", 823=>x"5700", 824=>x"4200",
---- 825=>x"2b00", 826=>x"3900", 827=>x"5200", 828=>x"4200",
---- 829=>x"2b00", 830=>x"3800", 831=>x"5600", 832=>x"4300",
---- 833=>x"2b00", 834=>x"3500", 835=>x"5500", 836=>x"5000",
---- 837=>x"2a00", 838=>x"3300", 839=>x"5200", 840=>x"5800",
---- 841=>x"2c00", 842=>x"3000", 843=>x"5000", 844=>x"5d00",
---- 845=>x"2c00", 846=>x"2b00", 847=>x"4800", 848=>x"6000",
---- 849=>x"2900", 850=>x"2500", 851=>x"3f00", 852=>x"5700",
---- 853=>x"2500", 854=>x"2600", 855=>x"4000", 856=>x"4f00",
---- 857=>x"2400", 858=>x"2700", 859=>x"4500", 860=>x"5400",
---- 861=>x"2500", 862=>x"2100", 863=>x"4000", 864=>x"5700",
---- 865=>x"2500", 866=>x"2300", 867=>x"3f00", 868=>x"5600",
---- 869=>x"2300", 870=>x"2500", 871=>x"3b00", 872=>x"5e00",
---- 873=>x"2700", 874=>x"2200", 875=>x"3800", 876=>x"9a00",
---- 877=>x"2c00", 878=>x"2300", 879=>x"3800", 880=>x"6a00",
---- 881=>x"3000", 882=>x"2300", 883=>x"3800", 884=>x"7200",
---- 885=>x"3b00", 886=>x"2400", 887=>x"3b00", 888=>x"7500",
---- 889=>x"3700", 890=>x"2300", 891=>x"3700", 892=>x"7300",
---- 893=>x"3700", 894=>x"2600", 895=>x"3b00", 896=>x"7300",
---- 897=>x"3f00", 898=>x"2500", 899=>x"3b00", 900=>x"7800",
---- 901=>x"3e00", 902=>x"2a00", 903=>x"3e00", 904=>x"7a00",
---- 905=>x"4700", 906=>x"2e00", 907=>x"3d00", 908=>x"7e00",
---- 909=>x"5100", 910=>x"3100", 911=>x"4000", 912=>x"8400",
---- 913=>x"5d00", 914=>x"3900", 915=>x"4000", 916=>x"8400",
---- 917=>x"6000", 918=>x"3700", 919=>x"3e00", 920=>x"8400",
---- 921=>x"5e00", 922=>x"3d00", 923=>x"4000", 924=>x"8800",
---- 925=>x"5a00", 926=>x"3d00", 927=>x"4300", 928=>x"9000",
---- 929=>x"6700", 930=>x"3e00", 931=>x"3d00", 932=>x"9200",
---- 933=>x"7300", 934=>x"c100", 935=>x"3a00", 936=>x"9500",
---- 937=>x"7c00", 938=>x"4700", 939=>x"3c00", 940=>x"9c00",
---- 941=>x"8300", 942=>x"4c00", 943=>x"3900", 944=>x"a300",
---- 945=>x"8800", 946=>x"4d00", 947=>x"3d00", 948=>x"ab00",
---- 949=>x"8600", 950=>x"5200", 951=>x"3e00", 952=>x"aa00",
---- 953=>x"8a00", 954=>x"5d00", 955=>x"4300", 956=>x"a800",
---- 957=>x"9100", 958=>x"6600", 959=>x"4800", 960=>x"ae00",
---- 961=>x"9600", 962=>x"7000", 963=>x"4d00", 964=>x"b000",
---- 965=>x"9900", 966=>x"7500", 967=>x"4d00", 968=>x"aa00",
---- 969=>x"9800", 970=>x"7800", 971=>x"5000", 972=>x"ab00",
---- 973=>x"9800", 974=>x"7700", 975=>x"5700", 976=>x"ab00",
---- 977=>x"9600", 978=>x"7600", 979=>x"5900", 980=>x"ae00",
---- 981=>x"9a00", 982=>x"7d00", 983=>x"5a00", 984=>x"ab00",
---- 985=>x"9c00", 986=>x"8200", 987=>x"6200", 988=>x"ab00",
---- 989=>x"9c00", 990=>x"8200", 991=>x"9300", 992=>x"ad00",
---- 993=>x"9b00", 994=>x"8500", 995=>x"7100", 996=>x"b800",
---- 997=>x"ab00", 998=>x"8f00", 999=>x"7600", 1000=>x"c600",
---- 1001=>x"c200", 1002=>x"a500", 1003=>x"7900", 1004=>x"c900",
---- 1005=>x"c800", 1006=>x"4600", 1007=>x"8900", 1008=>x"cb00",
---- 1009=>x"c500", 1010=>x"be00", 1011=>x"9d00", 1012=>x"ca00",
---- 1013=>x"c400", 1014=>x"bf00", 1015=>x"a500", 1016=>x"c600",
---- 1017=>x"c300", 1018=>x"4300", 1019=>x"a500", 1020=>x"c600",
---- 1021=>x"c100", 1022=>x"ba00", 1023=>x"9b00"),
----
---- 4 => (0=>x"9b00", 1=>x"9c00", 2=>x"a000", 3=>x"a400", 4=>x"9b00",
---- 5=>x"9c00", 6=>x"5d00", 7=>x"a400", 8=>x"9c00",
---- 9=>x"9b00", 10=>x"9f00", 11=>x"a300", 12=>x"9d00",
---- 13=>x"9900", 14=>x"9c00", 15=>x"a200", 16=>x"9b00",
---- 17=>x"9a00", 18=>x"a100", 19=>x"a400", 20=>x"9900",
---- 21=>x"9d00", 22=>x"a100", 23=>x"a600", 24=>x"9b00",
---- 25=>x"a000", 26=>x"a300", 27=>x"a600", 28=>x"9f00",
---- 29=>x"a300", 30=>x"a700", 31=>x"a800", 32=>x"a200",
---- 33=>x"a500", 34=>x"a800", 35=>x"a600", 36=>x"a200",
---- 37=>x"a700", 38=>x"a700", 39=>x"a600", 40=>x"a400",
---- 41=>x"a600", 42=>x"a400", 43=>x"a500", 44=>x"a600",
---- 45=>x"a600", 46=>x"a500", 47=>x"a200", 48=>x"a700",
---- 49=>x"a600", 50=>x"a800", 51=>x"a500", 52=>x"a600",
---- 53=>x"a700", 54=>x"a600", 55=>x"5900", 56=>x"a800",
---- 57=>x"a800", 58=>x"a600", 59=>x"a400", 60=>x"a900",
---- 61=>x"a700", 62=>x"a600", 63=>x"a300", 64=>x"aa00",
---- 65=>x"a700", 66=>x"a700", 67=>x"a200", 68=>x"a700",
---- 69=>x"a700", 70=>x"a900", 71=>x"a100", 72=>x"a600",
---- 73=>x"a600", 74=>x"a500", 75=>x"a000", 76=>x"a500",
---- 77=>x"a300", 78=>x"a200", 79=>x"a100", 80=>x"a400",
---- 81=>x"a300", 82=>x"a000", 83=>x"a000", 84=>x"a000",
---- 85=>x"9c00", 86=>x"a000", 87=>x"a300", 88=>x"9c00",
---- 89=>x"9c00", 90=>x"9d00", 91=>x"a200", 92=>x"9a00",
---- 93=>x"9b00", 94=>x"a000", 95=>x"a400", 96=>x"9500",
---- 97=>x"9a00", 98=>x"a100", 99=>x"a200", 100=>x"9200",
---- 101=>x"6500", 102=>x"a100", 103=>x"a600", 104=>x"9000",
---- 105=>x"9a00", 106=>x"a300", 107=>x"a400", 108=>x"9100",
---- 109=>x"9b00", 110=>x"a200", 111=>x"a300", 112=>x"9400",
---- 113=>x"9b00", 114=>x"a300", 115=>x"a600", 116=>x"9700",
---- 117=>x"9d00", 118=>x"a300", 119=>x"a400", 120=>x"9700",
---- 121=>x"9d00", 122=>x"a400", 123=>x"a800", 124=>x"9800",
---- 125=>x"9d00", 126=>x"a500", 127=>x"a800", 128=>x"9900",
---- 129=>x"9f00", 130=>x"a500", 131=>x"a700", 132=>x"9900",
---- 133=>x"a100", 134=>x"a600", 135=>x"a600", 136=>x"9600",
---- 137=>x"a200", 138=>x"a400", 139=>x"a800", 140=>x"9400",
---- 141=>x"a000", 142=>x"a700", 143=>x"a600", 144=>x"9600",
---- 145=>x"9f00", 146=>x"a400", 147=>x"a800", 148=>x"9800",
---- 149=>x"5f00", 150=>x"a600", 151=>x"a900", 152=>x"9800",
---- 153=>x"a000", 154=>x"a600", 155=>x"a700", 156=>x"9700",
---- 157=>x"9e00", 158=>x"a400", 159=>x"a800", 160=>x"9700",
---- 161=>x"9d00", 162=>x"a500", 163=>x"a600", 164=>x"9700",
---- 165=>x"9d00", 166=>x"a400", 167=>x"a700", 168=>x"9700",
---- 169=>x"9c00", 170=>x"a300", 171=>x"a800", 172=>x"9600",
---- 173=>x"9f00", 174=>x"a500", 175=>x"a800", 176=>x"9600",
---- 177=>x"9f00", 178=>x"a400", 179=>x"a600", 180=>x"9400",
---- 181=>x"9b00", 182=>x"a200", 183=>x"a600", 184=>x"9600",
---- 185=>x"9c00", 186=>x"a200", 187=>x"a500", 188=>x"9500",
---- 189=>x"9c00", 190=>x"a000", 191=>x"a400", 192=>x"9300",
---- 193=>x"9b00", 194=>x"a000", 195=>x"a500", 196=>x"9400",
---- 197=>x"9a00", 198=>x"a100", 199=>x"a400", 200=>x"9300",
---- 201=>x"9b00", 202=>x"a000", 203=>x"a300", 204=>x"9300",
---- 205=>x"9c00", 206=>x"a100", 207=>x"a700", 208=>x"9300",
---- 209=>x"9b00", 210=>x"9f00", 211=>x"a200", 212=>x"9200",
---- 213=>x"9b00", 214=>x"9f00", 215=>x"a400", 216=>x"9400",
---- 217=>x"9d00", 218=>x"9e00", 219=>x"a200", 220=>x"9400",
---- 221=>x"9c00", 222=>x"a000", 223=>x"a200", 224=>x"9100",
---- 225=>x"9900", 226=>x"9f00", 227=>x"a400", 228=>x"9500",
---- 229=>x"9a00", 230=>x"9f00", 231=>x"a200", 232=>x"9300",
---- 233=>x"9c00", 234=>x"a000", 235=>x"a300", 236=>x"9200",
---- 237=>x"9b00", 238=>x"a000", 239=>x"a400", 240=>x"9000",
---- 241=>x"9b00", 242=>x"a000", 243=>x"a300", 244=>x"9000",
---- 245=>x"9900", 246=>x"a000", 247=>x"a200", 248=>x"9300",
---- 249=>x"9900", 250=>x"9f00", 251=>x"a500", 252=>x"6c00",
---- 253=>x"9900", 254=>x"a000", 255=>x"a800", 256=>x"9100",
---- 257=>x"9900", 258=>x"a000", 259=>x"a400", 260=>x"9000",
---- 261=>x"9900", 262=>x"5e00", 263=>x"a700", 264=>x"9200",
---- 265=>x"9900", 266=>x"9f00", 267=>x"a600", 268=>x"9300",
---- 269=>x"9a00", 270=>x"a000", 271=>x"a300", 272=>x"9100",
---- 273=>x"9900", 274=>x"9f00", 275=>x"a400", 276=>x"9200",
---- 277=>x"9800", 278=>x"9b00", 279=>x"a400", 280=>x"9400",
---- 281=>x"9700", 282=>x"9e00", 283=>x"a600", 284=>x"9500",
---- 285=>x"9c00", 286=>x"a100", 287=>x"a500", 288=>x"9300",
---- 289=>x"9f00", 290=>x"a400", 291=>x"a500", 292=>x"9500",
---- 293=>x"9b00", 294=>x"a100", 295=>x"a800", 296=>x"9400",
---- 297=>x"9d00", 298=>x"a400", 299=>x"a900", 300=>x"9400",
---- 301=>x"9b00", 302=>x"a400", 303=>x"ab00", 304=>x"6a00",
---- 305=>x"9b00", 306=>x"a300", 307=>x"a800", 308=>x"9200",
---- 309=>x"9d00", 310=>x"a400", 311=>x"a800", 312=>x"9400",
---- 313=>x"9e00", 314=>x"a500", 315=>x"aa00", 316=>x"9900",
---- 317=>x"6100", 318=>x"a600", 319=>x"ab00", 320=>x"9800",
---- 321=>x"9e00", 322=>x"a400", 323=>x"aa00", 324=>x"9500",
---- 325=>x"9e00", 326=>x"a400", 327=>x"a800", 328=>x"9700",
---- 329=>x"9f00", 330=>x"a400", 331=>x"a900", 332=>x"9600",
---- 333=>x"9f00", 334=>x"a300", 335=>x"5500", 336=>x"9600",
---- 337=>x"6200", 338=>x"a400", 339=>x"a900", 340=>x"9700",
---- 341=>x"9f00", 342=>x"a400", 343=>x"a900", 344=>x"9300",
---- 345=>x"a000", 346=>x"a500", 347=>x"ab00", 348=>x"9600",
---- 349=>x"9e00", 350=>x"a500", 351=>x"ab00", 352=>x"9600",
---- 353=>x"9f00", 354=>x"a500", 355=>x"ac00", 356=>x"9700",
---- 357=>x"9d00", 358=>x"a500", 359=>x"ab00", 360=>x"9900",
---- 361=>x"9e00", 362=>x"a600", 363=>x"ad00", 364=>x"9800",
---- 365=>x"a100", 366=>x"a700", 367=>x"ab00", 368=>x"9800",
---- 369=>x"a000", 370=>x"a900", 371=>x"ac00", 372=>x"9800",
---- 373=>x"a000", 374=>x"a800", 375=>x"ac00", 376=>x"9600",
---- 377=>x"9d00", 378=>x"a600", 379=>x"a900", 380=>x"9600",
---- 381=>x"9d00", 382=>x"a600", 383=>x"aa00", 384=>x"9600",
---- 385=>x"9d00", 386=>x"a400", 387=>x"a900", 388=>x"9600",
---- 389=>x"9d00", 390=>x"a500", 391=>x"a800", 392=>x"9700",
---- 393=>x"9e00", 394=>x"a500", 395=>x"aa00", 396=>x"9500",
---- 397=>x"9e00", 398=>x"a500", 399=>x"aa00", 400=>x"9600",
---- 401=>x"9e00", 402=>x"a600", 403=>x"aa00", 404=>x"9600",
---- 405=>x"a000", 406=>x"a800", 407=>x"ac00", 408=>x"9400",
---- 409=>x"9f00", 410=>x"a500", 411=>x"aa00", 412=>x"9500",
---- 413=>x"9d00", 414=>x"a500", 415=>x"a700", 416=>x"9200",
---- 417=>x"9e00", 418=>x"a800", 419=>x"aa00", 420=>x"9400",
---- 421=>x"9f00", 422=>x"a400", 423=>x"5400", 424=>x"9400",
---- 425=>x"9c00", 426=>x"a200", 427=>x"a900", 428=>x"9400",
---- 429=>x"9900", 430=>x"a500", 431=>x"a900", 432=>x"9000",
---- 433=>x"9c00", 434=>x"a200", 435=>x"ab00", 436=>x"6d00",
---- 437=>x"9a00", 438=>x"a400", 439=>x"a900", 440=>x"9200",
---- 441=>x"9b00", 442=>x"a200", 443=>x"aa00", 444=>x"9200",
---- 445=>x"9b00", 446=>x"a300", 447=>x"a900", 448=>x"9200",
---- 449=>x"9b00", 450=>x"a200", 451=>x"a600", 452=>x"9400",
---- 453=>x"9b00", 454=>x"a300", 455=>x"a700", 456=>x"9100",
---- 457=>x"9b00", 458=>x"a400", 459=>x"a900", 460=>x"9100",
---- 461=>x"9a00", 462=>x"a400", 463=>x"aa00", 464=>x"8f00",
---- 465=>x"9800", 466=>x"a300", 467=>x"a800", 468=>x"9100",
---- 469=>x"9b00", 470=>x"a400", 471=>x"ab00", 472=>x"9000",
---- 473=>x"9800", 474=>x"a100", 475=>x"5500", 476=>x"9000",
---- 477=>x"9700", 478=>x"a500", 479=>x"ad00", 480=>x"9400",
---- 481=>x"9d00", 482=>x"a400", 483=>x"aa00", 484=>x"9300",
---- 485=>x"9c00", 486=>x"a300", 487=>x"a900", 488=>x"8f00",
---- 489=>x"9a00", 490=>x"5c00", 491=>x"a900", 492=>x"9000",
---- 493=>x"9c00", 494=>x"a400", 495=>x"a800", 496=>x"9300",
---- 497=>x"9c00", 498=>x"5d00", 499=>x"a900", 500=>x"9200",
---- 501=>x"9a00", 502=>x"a300", 503=>x"ab00", 504=>x"9100",
---- 505=>x"9700", 506=>x"a000", 507=>x"aa00", 508=>x"9200",
---- 509=>x"9900", 510=>x"a100", 511=>x"ab00", 512=>x"9100",
---- 513=>x"9a00", 514=>x"a200", 515=>x"ab00", 516=>x"9000",
---- 517=>x"9800", 518=>x"a200", 519=>x"aa00", 520=>x"8f00",
---- 521=>x"9a00", 522=>x"a400", 523=>x"a900", 524=>x"8f00",
---- 525=>x"9800", 526=>x"a300", 527=>x"ab00", 528=>x"8e00",
---- 529=>x"9800", 530=>x"a400", 531=>x"ac00", 532=>x"8e00",
---- 533=>x"9a00", 534=>x"a400", 535=>x"ad00", 536=>x"8d00",
---- 537=>x"9a00", 538=>x"a400", 539=>x"ac00", 540=>x"8d00",
---- 541=>x"9a00", 542=>x"a400", 543=>x"aa00", 544=>x"8f00",
---- 545=>x"9900", 546=>x"a200", 547=>x"ac00", 548=>x"9000",
---- 549=>x"9800", 550=>x"a400", 551=>x"aa00", 552=>x"8d00",
---- 553=>x"9b00", 554=>x"a400", 555=>x"ab00", 556=>x"6e00",
---- 557=>x"9c00", 558=>x"a300", 559=>x"ab00", 560=>x"8e00",
---- 561=>x"9900", 562=>x"a300", 563=>x"ab00", 564=>x"8c00",
---- 565=>x"9700", 566=>x"a500", 567=>x"ab00", 568=>x"8c00",
---- 569=>x"9800", 570=>x"a200", 571=>x"a900", 572=>x"8d00",
---- 573=>x"9700", 574=>x"a100", 575=>x"a900", 576=>x"8b00",
---- 577=>x"9600", 578=>x"a100", 579=>x"aa00", 580=>x"8900",
---- 581=>x"9700", 582=>x"a200", 583=>x"aa00", 584=>x"8a00",
---- 585=>x"9700", 586=>x"a200", 587=>x"a900", 588=>x"8b00",
---- 589=>x"9600", 590=>x"a200", 591=>x"aa00", 592=>x"8b00",
---- 593=>x"9800", 594=>x"a200", 595=>x"ab00", 596=>x"8800",
---- 597=>x"9700", 598=>x"a100", 599=>x"a800", 600=>x"8a00",
---- 601=>x"9600", 602=>x"5f00", 603=>x"a900", 604=>x"8c00",
---- 605=>x"9600", 606=>x"9f00", 607=>x"a800", 608=>x"8c00",
---- 609=>x"9900", 610=>x"9f00", 611=>x"a800", 612=>x"8a00",
---- 613=>x"9500", 614=>x"9f00", 615=>x"a500", 616=>x"8900",
---- 617=>x"9400", 618=>x"9f00", 619=>x"a600", 620=>x"8900",
---- 621=>x"9600", 622=>x"9f00", 623=>x"a700", 624=>x"8700",
---- 625=>x"9600", 626=>x"a000", 627=>x"a700", 628=>x"8600",
---- 629=>x"9700", 630=>x"9f00", 631=>x"a700", 632=>x"8400",
---- 633=>x"9500", 634=>x"a000", 635=>x"a800", 636=>x"8600",
---- 637=>x"9600", 638=>x"a100", 639=>x"a800", 640=>x"8600",
---- 641=>x"9400", 642=>x"a200", 643=>x"a900", 644=>x"7500",
---- 645=>x"6b00", 646=>x"a100", 647=>x"a800", 648=>x"8e00",
---- 649=>x"9700", 650=>x"9f00", 651=>x"a600", 652=>x"9300",
---- 653=>x"9a00", 654=>x"a200", 655=>x"a800", 656=>x"9200",
---- 657=>x"9b00", 658=>x"a300", 659=>x"a500", 660=>x"9400",
---- 661=>x"9d00", 662=>x"a300", 663=>x"a700", 664=>x"9800",
---- 665=>x"9c00", 666=>x"a100", 667=>x"a800", 668=>x"9700",
---- 669=>x"9d00", 670=>x"a200", 671=>x"a600", 672=>x"9700",
---- 673=>x"9e00", 674=>x"a300", 675=>x"a700", 676=>x"9700",
---- 677=>x"9d00", 678=>x"a400", 679=>x"a700", 680=>x"9600",
---- 681=>x"9e00", 682=>x"a300", 683=>x"a500", 684=>x"9500",
---- 685=>x"9d00", 686=>x"a200", 687=>x"a600", 688=>x"9500",
---- 689=>x"9b00", 690=>x"a200", 691=>x"a800", 692=>x"9700",
---- 693=>x"9f00", 694=>x"a300", 695=>x"a700", 696=>x"9700",
---- 697=>x"a100", 698=>x"a600", 699=>x"a900", 700=>x"9800",
---- 701=>x"9d00", 702=>x"a400", 703=>x"ad00", 704=>x"9700",
---- 705=>x"9e00", 706=>x"a500", 707=>x"ac00", 708=>x"9700",
---- 709=>x"9f00", 710=>x"a600", 711=>x"ab00", 712=>x"9700",
---- 713=>x"9e00", 714=>x"a300", 715=>x"ab00", 716=>x"9700",
---- 717=>x"9c00", 718=>x"a200", 719=>x"aa00", 720=>x"9600",
---- 721=>x"9e00", 722=>x"a200", 723=>x"aa00", 724=>x"9300",
---- 725=>x"9e00", 726=>x"a200", 727=>x"a800", 728=>x"9100",
---- 729=>x"9900", 730=>x"a000", 731=>x"a700", 732=>x"9000",
---- 733=>x"9600", 734=>x"9d00", 735=>x"a700", 736=>x"8c00",
---- 737=>x"9400", 738=>x"9c00", 739=>x"a600", 740=>x"8a00",
---- 741=>x"9200", 742=>x"9a00", 743=>x"a500", 744=>x"8d00",
---- 745=>x"9200", 746=>x"9a00", 747=>x"a800", 748=>x"8a00",
---- 749=>x"9500", 750=>x"9c00", 751=>x"a500", 752=>x"8a00",
---- 753=>x"9300", 754=>x"9e00", 755=>x"a600", 756=>x"8a00",
---- 757=>x"9300", 758=>x"9c00", 759=>x"a700", 760=>x"8b00",
---- 761=>x"9500", 762=>x"9f00", 763=>x"a800", 764=>x"8b00",
---- 765=>x"9600", 766=>x"9e00", 767=>x"a700", 768=>x"8f00",
---- 769=>x"9900", 770=>x"a000", 771=>x"a600", 772=>x"8d00",
---- 773=>x"9900", 774=>x"a000", 775=>x"a600", 776=>x"8b00",
---- 777=>x"9600", 778=>x"a000", 779=>x"a600", 780=>x"8c00",
---- 781=>x"9600", 782=>x"9e00", 783=>x"a600", 784=>x"8900",
---- 785=>x"9400", 786=>x"9d00", 787=>x"a800", 788=>x"8500",
---- 789=>x"8f00", 790=>x"9c00", 791=>x"a400", 792=>x"7e00",
---- 793=>x"8d00", 794=>x"9c00", 795=>x"a500", 796=>x"7700",
---- 797=>x"8900", 798=>x"9a00", 799=>x"a400", 800=>x"7100",
---- 801=>x"8700", 802=>x"9800", 803=>x"a300", 804=>x"7100",
---- 805=>x"8900", 806=>x"9900", 807=>x"a200", 808=>x"6f00",
---- 809=>x"8500", 810=>x"9a00", 811=>x"a300", 812=>x"7200",
---- 813=>x"8800", 814=>x"9900", 815=>x"a400", 816=>x"7500",
---- 817=>x"8a00", 818=>x"9900", 819=>x"a700", 820=>x"7000",
---- 821=>x"8800", 822=>x"9b00", 823=>x"a500", 824=>x"6f00",
---- 825=>x"8800", 826=>x"6500", 827=>x"a400", 828=>x"7000",
---- 829=>x"8900", 830=>x"9900", 831=>x"a500", 832=>x"7100",
---- 833=>x"8a00", 834=>x"9d00", 835=>x"a600", 836=>x"7100",
---- 837=>x"8c00", 838=>x"9c00", 839=>x"a500", 840=>x"7200",
---- 841=>x"8d00", 842=>x"9c00", 843=>x"a600", 844=>x"7100",
---- 845=>x"8e00", 846=>x"9c00", 847=>x"a600", 848=>x"6f00",
---- 849=>x"8c00", 850=>x"9a00", 851=>x"a500", 852=>x"7000",
---- 853=>x"8d00", 854=>x"9a00", 855=>x"a500", 856=>x"6f00",
---- 857=>x"8e00", 858=>x"9a00", 859=>x"a500", 860=>x"6f00",
---- 861=>x"8b00", 862=>x"9a00", 863=>x"a800", 864=>x"6c00",
---- 865=>x"8a00", 866=>x"9c00", 867=>x"a700", 868=>x"6b00",
---- 869=>x"8b00", 870=>x"9d00", 871=>x"a800", 872=>x"6c00",
---- 873=>x"8a00", 874=>x"9c00", 875=>x"a800", 876=>x"6700",
---- 877=>x"8900", 878=>x"9a00", 879=>x"a700", 880=>x"6400",
---- 881=>x"8a00", 882=>x"9d00", 883=>x"a800", 884=>x"6300",
---- 885=>x"8800", 886=>x"9b00", 887=>x"a800", 888=>x"5f00",
---- 889=>x"8500", 890=>x"9c00", 891=>x"a700", 892=>x"6300",
---- 893=>x"8600", 894=>x"9b00", 895=>x"a800", 896=>x"9e00",
---- 897=>x"8500", 898=>x"9800", 899=>x"a700", 900=>x"6100",
---- 901=>x"8500", 902=>x"9600", 903=>x"a600", 904=>x"5d00",
---- 905=>x"8400", 906=>x"9800", 907=>x"a300", 908=>x"5e00",
---- 909=>x"8400", 910=>x"9600", 911=>x"a500", 912=>x"5d00",
---- 913=>x"8300", 914=>x"9600", 915=>x"a600", 916=>x"5c00",
---- 917=>x"8000", 918=>x"9500", 919=>x"a200", 920=>x"5b00",
---- 921=>x"7e00", 922=>x"9200", 923=>x"a000", 924=>x"5c00",
---- 925=>x"7e00", 926=>x"9500", 927=>x"a100", 928=>x"5500",
---- 929=>x"7d00", 930=>x"9100", 931=>x"9e00", 932=>x"5800",
---- 933=>x"7b00", 934=>x"8e00", 935=>x"9e00", 936=>x"5700",
---- 937=>x"7800", 938=>x"8f00", 939=>x"9e00", 940=>x"5500",
---- 941=>x"7600", 942=>x"9000", 943=>x"9f00", 944=>x"5900",
---- 945=>x"7a00", 946=>x"9200", 947=>x"9f00", 948=>x"5a00",
---- 949=>x"7700", 950=>x"8f00", 951=>x"9d00", 952=>x"5900",
---- 953=>x"7600", 954=>x"8e00", 955=>x"9d00", 956=>x"5b00",
---- 957=>x"8a00", 958=>x"8e00", 959=>x"9d00", 960=>x"5e00",
---- 961=>x"7300", 962=>x"8d00", 963=>x"9c00", 964=>x"5c00",
---- 965=>x"7400", 966=>x"8a00", 967=>x"9d00", 968=>x"5c00",
---- 969=>x"7500", 970=>x"8b00", 971=>x"9c00", 972=>x"5c00",
---- 973=>x"7500", 974=>x"8c00", 975=>x"9b00", 976=>x"6000",
---- 977=>x"7100", 978=>x"8b00", 979=>x"9a00", 980=>x"5c00",
---- 981=>x"7200", 982=>x"8800", 983=>x"9900", 984=>x"5d00",
---- 985=>x"7100", 986=>x"8800", 987=>x"9900", 988=>x"6100",
---- 989=>x"7300", 990=>x"8500", 991=>x"9700", 992=>x"6300",
---- 993=>x"7300", 994=>x"8300", 995=>x"9600", 996=>x"6400",
---- 997=>x"7100", 998=>x"8600", 999=>x"9800", 1000=>x"6600",
---- 1001=>x"7600", 1002=>x"8700", 1003=>x"9a00", 1004=>x"6900",
---- 1005=>x"7700", 1006=>x"8500", 1007=>x"9800", 1008=>x"6a00",
---- 1009=>x"7500", 1010=>x"8500", 1011=>x"9700", 1012=>x"6c00",
---- 1013=>x"7400", 1014=>x"8600", 1015=>x"9800", 1016=>x"6e00",
---- 1017=>x"7300", 1018=>x"8800", 1019=>x"9a00", 1020=>x"6a00",
---- 1021=>x"7800", 1022=>x"8900", 1023=>x"9900"),
----
---- 5 => (0=>x"a600", 1=>x"a700", 2=>x"ae00", 3=>x"ad00", 4=>x"a600",
---- 5=>x"a700", 6=>x"ad00", 7=>x"ad00", 8=>x"a400",
---- 9=>x"a700", 10=>x"ac00", 11=>x"ad00", 12=>x"a600",
---- 13=>x"a900", 14=>x"ab00", 15=>x"ac00", 16=>x"a800",
---- 17=>x"ab00", 18=>x"ac00", 19=>x"ac00", 20=>x"a800",
---- 21=>x"a800", 22=>x"ab00", 23=>x"ab00", 24=>x"a900",
---- 25=>x"a900", 26=>x"a900", 27=>x"a800", 28=>x"a900",
---- 29=>x"a800", 30=>x"a900", 31=>x"a800", 32=>x"a700",
---- 33=>x"a900", 34=>x"a500", 35=>x"a700", 36=>x"a700",
---- 37=>x"a400", 38=>x"a600", 39=>x"a400", 40=>x"a700",
---- 41=>x"a400", 42=>x"a500", 43=>x"a200", 44=>x"a600",
---- 45=>x"a500", 46=>x"a400", 47=>x"a300", 48=>x"5b00",
---- 49=>x"a400", 50=>x"a300", 51=>x"9f00", 52=>x"a100",
---- 53=>x"a100", 54=>x"a100", 55=>x"9e00", 56=>x"a000",
---- 57=>x"9e00", 58=>x"9e00", 59=>x"9e00", 60=>x"a000",
---- 61=>x"9f00", 62=>x"9d00", 63=>x"9d00", 64=>x"9f00",
---- 65=>x"9f00", 66=>x"9e00", 67=>x"9e00", 68=>x"a000",
---- 69=>x"a100", 70=>x"9d00", 71=>x"9e00", 72=>x"9c00",
---- 73=>x"9e00", 74=>x"9e00", 75=>x"9f00", 76=>x"9e00",
---- 77=>x"9e00", 78=>x"a000", 79=>x"a100", 80=>x"9f00",
---- 81=>x"9f00", 82=>x"a100", 83=>x"a100", 84=>x"a000",
---- 85=>x"9e00", 86=>x"a000", 87=>x"a000", 88=>x"a100",
---- 89=>x"9f00", 90=>x"9f00", 91=>x"9f00", 92=>x"a500",
---- 93=>x"a300", 94=>x"a000", 95=>x"a100", 96=>x"a200",
---- 97=>x"a100", 98=>x"9f00", 99=>x"a100", 100=>x"a300",
---- 101=>x"a100", 102=>x"a100", 103=>x"a100", 104=>x"a400",
---- 105=>x"a200", 106=>x"a200", 107=>x"a200", 108=>x"a400",
---- 109=>x"a200", 110=>x"a200", 111=>x"5c00", 112=>x"a400",
---- 113=>x"a300", 114=>x"a200", 115=>x"a600", 116=>x"a500",
---- 117=>x"a600", 118=>x"a400", 119=>x"a400", 120=>x"a400",
---- 121=>x"a700", 122=>x"a400", 123=>x"a300", 124=>x"a500",
---- 125=>x"a500", 126=>x"a600", 127=>x"a500", 128=>x"a600",
---- 129=>x"a500", 130=>x"a400", 131=>x"a500", 132=>x"a500",
---- 133=>x"a600", 134=>x"a900", 135=>x"a300", 136=>x"a700",
---- 137=>x"a400", 138=>x"a500", 139=>x"a300", 140=>x"a800",
---- 141=>x"a400", 142=>x"a400", 143=>x"a600", 144=>x"ab00",
---- 145=>x"a600", 146=>x"a600", 147=>x"a500", 148=>x"a700",
---- 149=>x"a600", 150=>x"5900", 151=>x"a400", 152=>x"a600",
---- 153=>x"a800", 154=>x"a700", 155=>x"a400", 156=>x"a800",
---- 157=>x"a900", 158=>x"a800", 159=>x"a600", 160=>x"a800",
---- 161=>x"a800", 162=>x"a700", 163=>x"a700", 164=>x"a700",
---- 165=>x"a700", 166=>x"a900", 167=>x"a700", 168=>x"a800",
---- 169=>x"a800", 170=>x"5700", 171=>x"a600", 172=>x"a700",
---- 173=>x"a800", 174=>x"a700", 175=>x"a600", 176=>x"a800",
---- 177=>x"a600", 178=>x"a600", 179=>x"a500", 180=>x"a700",
---- 181=>x"a800", 182=>x"a400", 183=>x"a600", 184=>x"a500",
---- 185=>x"a800", 186=>x"a600", 187=>x"a400", 188=>x"a700",
---- 189=>x"a700", 190=>x"a600", 191=>x"a600", 192=>x"a500",
---- 193=>x"a700", 194=>x"a800", 195=>x"a700", 196=>x"a500",
---- 197=>x"a700", 198=>x"a500", 199=>x"a600", 200=>x"a600",
---- 201=>x"a600", 202=>x"a500", 203=>x"a500", 204=>x"a500",
---- 205=>x"a500", 206=>x"a800", 207=>x"a700", 208=>x"a600",
---- 209=>x"a600", 210=>x"a700", 211=>x"a600", 212=>x"a400",
---- 213=>x"a200", 214=>x"a400", 215=>x"a600", 216=>x"a500",
---- 217=>x"a300", 218=>x"a300", 219=>x"a300", 220=>x"a500",
---- 221=>x"a500", 222=>x"a600", 223=>x"a300", 224=>x"a500",
---- 225=>x"a500", 226=>x"a500", 227=>x"a400", 228=>x"a500",
---- 229=>x"a300", 230=>x"a300", 231=>x"a200", 232=>x"a600",
---- 233=>x"a300", 234=>x"a400", 235=>x"a400", 236=>x"a300",
---- 237=>x"a500", 238=>x"a400", 239=>x"a200", 240=>x"a500",
---- 241=>x"a400", 242=>x"a400", 243=>x"a300", 244=>x"a500",
---- 245=>x"a700", 246=>x"a700", 247=>x"a600", 248=>x"a600",
---- 249=>x"a800", 250=>x"a600", 251=>x"a500", 252=>x"a900",
---- 253=>x"a400", 254=>x"a800", 255=>x"a700", 256=>x"a700",
---- 257=>x"a700", 258=>x"a900", 259=>x"a800", 260=>x"a800",
---- 261=>x"a800", 262=>x"aa00", 263=>x"a800", 264=>x"a600",
---- 265=>x"a500", 266=>x"a700", 267=>x"a800", 268=>x"a700",
---- 269=>x"a600", 270=>x"a700", 271=>x"a600", 272=>x"a700",
---- 273=>x"a600", 274=>x"a900", 275=>x"a800", 276=>x"a400",
---- 277=>x"a700", 278=>x"aa00", 279=>x"aa00", 280=>x"a600",
---- 281=>x"a900", 282=>x"a900", 283=>x"ac00", 284=>x"a700",
---- 285=>x"ab00", 286=>x"ac00", 287=>x"ad00", 288=>x"a900",
---- 289=>x"ab00", 290=>x"ac00", 291=>x"ac00", 292=>x"aa00",
---- 293=>x"ab00", 294=>x"5100", 295=>x"ad00", 296=>x"ab00",
---- 297=>x"ac00", 298=>x"b000", 299=>x"b000", 300=>x"ab00",
---- 301=>x"ad00", 302=>x"af00", 303=>x"ae00", 304=>x"ac00",
---- 305=>x"ae00", 306=>x"ad00", 307=>x"ad00", 308=>x"ab00",
---- 309=>x"ac00", 310=>x"ae00", 311=>x"ab00", 312=>x"ad00",
---- 313=>x"ac00", 314=>x"ad00", 315=>x"ae00", 316=>x"ab00",
---- 317=>x"ad00", 318=>x"ac00", 319=>x"ac00", 320=>x"ab00",
---- 321=>x"a900", 322=>x"ab00", 323=>x"ac00", 324=>x"aa00",
---- 325=>x"ac00", 326=>x"ac00", 327=>x"ac00", 328=>x"ac00",
---- 329=>x"aa00", 330=>x"ac00", 331=>x"ab00", 332=>x"a900",
---- 333=>x"aa00", 334=>x"ab00", 335=>x"a800", 336=>x"ab00",
---- 337=>x"ad00", 338=>x"ae00", 339=>x"ad00", 340=>x"ac00",
---- 341=>x"ac00", 342=>x"ab00", 343=>x"ae00", 344=>x"ab00",
---- 345=>x"ac00", 346=>x"ad00", 347=>x"ad00", 348=>x"a900",
---- 349=>x"ad00", 350=>x"ac00", 351=>x"ac00", 352=>x"ac00",
---- 353=>x"ad00", 354=>x"af00", 355=>x"af00", 356=>x"ae00",
---- 357=>x"ab00", 358=>x"ae00", 359=>x"af00", 360=>x"ac00",
---- 361=>x"ac00", 362=>x"ae00", 363=>x"af00", 364=>x"ac00",
---- 365=>x"ad00", 366=>x"ac00", 367=>x"ad00", 368=>x"ac00",
---- 369=>x"ab00", 370=>x"ad00", 371=>x"ad00", 372=>x"ac00",
---- 373=>x"aa00", 374=>x"ac00", 375=>x"ac00", 376=>x"ac00",
---- 377=>x"ab00", 378=>x"aa00", 379=>x"b000", 380=>x"ac00",
---- 381=>x"ac00", 382=>x"ab00", 383=>x"ab00", 384=>x"ab00",
---- 385=>x"aa00", 386=>x"aa00", 387=>x"aa00", 388=>x"a900",
---- 389=>x"5400", 390=>x"aa00", 391=>x"ac00", 392=>x"ad00",
---- 393=>x"ac00", 394=>x"a900", 395=>x"ac00", 396=>x"ac00",
---- 397=>x"aa00", 398=>x"ad00", 399=>x"ad00", 400=>x"ac00",
---- 401=>x"aa00", 402=>x"ac00", 403=>x"aa00", 404=>x"ab00",
---- 405=>x"5400", 406=>x"ac00", 407=>x"ac00", 408=>x"ac00",
---- 409=>x"ab00", 410=>x"ac00", 411=>x"af00", 412=>x"ac00",
---- 413=>x"ab00", 414=>x"ad00", 415=>x"ae00", 416=>x"ab00",
---- 417=>x"ad00", 418=>x"ad00", 419=>x"ac00", 420=>x"ae00",
---- 421=>x"ac00", 422=>x"ad00", 423=>x"ad00", 424=>x"ad00",
---- 425=>x"ae00", 426=>x"ad00", 427=>x"ac00", 428=>x"ab00",
---- 429=>x"ad00", 430=>x"ab00", 431=>x"ab00", 432=>x"ae00",
---- 433=>x"ab00", 434=>x"ac00", 435=>x"af00", 436=>x"aa00",
---- 437=>x"5200", 438=>x"ad00", 439=>x"ae00", 440=>x"ab00",
---- 441=>x"ac00", 442=>x"ae00", 443=>x"ae00", 444=>x"ae00",
---- 445=>x"ac00", 446=>x"aa00", 447=>x"af00", 448=>x"ab00",
---- 449=>x"ad00", 450=>x"5200", 451=>x"ac00", 452=>x"ab00",
---- 453=>x"af00", 454=>x"ad00", 455=>x"ad00", 456=>x"ac00",
---- 457=>x"ac00", 458=>x"ae00", 459=>x"af00", 460=>x"ab00",
---- 461=>x"ae00", 462=>x"ad00", 463=>x"5100", 464=>x"ab00",
---- 465=>x"ad00", 466=>x"ae00", 467=>x"b000", 468=>x"ad00",
---- 469=>x"ae00", 470=>x"ae00", 471=>x"b000", 472=>x"ac00",
---- 473=>x"ad00", 474=>x"af00", 475=>x"ad00", 476=>x"ad00",
---- 477=>x"ad00", 478=>x"b000", 479=>x"ad00", 480=>x"aa00",
---- 481=>x"ae00", 482=>x"b000", 483=>x"af00", 484=>x"ac00",
---- 485=>x"ac00", 486=>x"b000", 487=>x"af00", 488=>x"ac00",
---- 489=>x"ae00", 490=>x"af00", 491=>x"af00", 492=>x"ad00",
---- 493=>x"b000", 494=>x"b100", 495=>x"b200", 496=>x"ad00",
---- 497=>x"ad00", 498=>x"b100", 499=>x"b200", 500=>x"ae00",
---- 501=>x"ad00", 502=>x"b000", 503=>x"af00", 504=>x"ae00",
---- 505=>x"ac00", 506=>x"b000", 507=>x"af00", 508=>x"af00",
---- 509=>x"af00", 510=>x"ae00", 511=>x"af00", 512=>x"af00",
---- 513=>x"b100", 514=>x"af00", 515=>x"b000", 516=>x"ae00",
---- 517=>x"b000", 518=>x"b000", 519=>x"b300", 520=>x"ac00",
---- 521=>x"b100", 522=>x"b000", 523=>x"b100", 524=>x"ae00",
---- 525=>x"b000", 526=>x"ae00", 527=>x"b100", 528=>x"b000",
---- 529=>x"ae00", 530=>x"b000", 531=>x"b200", 532=>x"b000",
---- 533=>x"b200", 534=>x"af00", 535=>x"b100", 536=>x"b000",
---- 537=>x"b000", 538=>x"b100", 539=>x"b200", 540=>x"b200",
---- 541=>x"b100", 542=>x"b100", 543=>x"b600", 544=>x"b100",
---- 545=>x"b200", 546=>x"b400", 547=>x"b300", 548=>x"b000",
---- 549=>x"b300", 550=>x"b400", 551=>x"b400", 552=>x"af00",
---- 553=>x"b200", 554=>x"b400", 555=>x"b500", 556=>x"ae00",
---- 557=>x"b100", 558=>x"b300", 559=>x"b600", 560=>x"b100",
---- 561=>x"b300", 562=>x"b300", 563=>x"b600", 564=>x"b000",
---- 565=>x"b200", 566=>x"b300", 567=>x"b600", 568=>x"ae00",
---- 569=>x"4e00", 570=>x"b500", 571=>x"b400", 572=>x"af00",
---- 573=>x"b300", 574=>x"b500", 575=>x"b500", 576=>x"ad00",
---- 577=>x"b200", 578=>x"b400", 579=>x"b400", 580=>x"af00",
---- 581=>x"b300", 582=>x"b200", 583=>x"b200", 584=>x"af00",
---- 585=>x"b200", 586=>x"b400", 587=>x"b500", 588=>x"af00",
---- 589=>x"b000", 590=>x"b200", 591=>x"b300", 592=>x"af00",
---- 593=>x"b100", 594=>x"b200", 595=>x"b300", 596=>x"ae00",
---- 597=>x"b000", 598=>x"b200", 599=>x"b400", 600=>x"ac00",
---- 601=>x"ae00", 602=>x"b200", 603=>x"b100", 604=>x"ab00",
---- 605=>x"ae00", 606=>x"b000", 607=>x"ae00", 608=>x"ad00",
---- 609=>x"af00", 610=>x"ac00", 611=>x"ac00", 612=>x"ac00",
---- 613=>x"ae00", 614=>x"ac00", 615=>x"ac00", 616=>x"ac00",
---- 617=>x"ae00", 618=>x"ac00", 619=>x"ac00", 620=>x"ab00",
---- 621=>x"ad00", 622=>x"ad00", 623=>x"ab00", 624=>x"ab00",
---- 625=>x"ad00", 626=>x"af00", 627=>x"4f00", 628=>x"ab00",
---- 629=>x"ad00", 630=>x"b000", 631=>x"b000", 632=>x"ac00",
---- 633=>x"ae00", 634=>x"af00", 635=>x"af00", 636=>x"ac00",
---- 637=>x"ae00", 638=>x"af00", 639=>x"b000", 640=>x"ad00",
---- 641=>x"ac00", 642=>x"ae00", 643=>x"ad00", 644=>x"a900",
---- 645=>x"ac00", 646=>x"ad00", 647=>x"ae00", 648=>x"aa00",
---- 649=>x"ad00", 650=>x"af00", 651=>x"af00", 652=>x"ab00",
---- 653=>x"ae00", 654=>x"ac00", 655=>x"ae00", 656=>x"aa00",
---- 657=>x"ab00", 658=>x"ab00", 659=>x"ad00", 660=>x"a800",
---- 661=>x"aa00", 662=>x"aa00", 663=>x"ab00", 664=>x"a700",
---- 665=>x"a900", 666=>x"ab00", 667=>x"ad00", 668=>x"a700",
---- 669=>x"a900", 670=>x"ab00", 671=>x"b000", 672=>x"a700",
---- 673=>x"ac00", 674=>x"ab00", 675=>x"ac00", 676=>x"aa00",
---- 677=>x"a900", 678=>x"a900", 679=>x"ac00", 680=>x"a800",
---- 681=>x"ab00", 682=>x"ab00", 683=>x"af00", 684=>x"a800",
---- 685=>x"5500", 686=>x"ac00", 687=>x"af00", 688=>x"a900",
---- 689=>x"ab00", 690=>x"ad00", 691=>x"b000", 692=>x"ab00",
---- 693=>x"ac00", 694=>x"ac00", 695=>x"ae00", 696=>x"ad00",
---- 697=>x"ad00", 698=>x"ae00", 699=>x"af00", 700=>x"af00",
---- 701=>x"ad00", 702=>x"b000", 703=>x"b200", 704=>x"af00",
---- 705=>x"b000", 706=>x"b200", 707=>x"b100", 708=>x"b000",
---- 709=>x"af00", 710=>x"b000", 711=>x"af00", 712=>x"af00",
---- 713=>x"b000", 714=>x"b200", 715=>x"b200", 716=>x"ae00",
---- 717=>x"b000", 718=>x"b200", 719=>x"b000", 720=>x"ad00",
---- 721=>x"b100", 722=>x"b200", 723=>x"b300", 724=>x"af00",
---- 725=>x"b200", 726=>x"b300", 727=>x"b300", 728=>x"b000",
---- 729=>x"b300", 730=>x"b300", 731=>x"b300", 732=>x"af00",
---- 733=>x"b300", 734=>x"b200", 735=>x"b200", 736=>x"ae00",
---- 737=>x"af00", 738=>x"b200", 739=>x"b100", 740=>x"af00",
---- 741=>x"b000", 742=>x"b100", 743=>x"b100", 744=>x"ad00",
---- 745=>x"af00", 746=>x"b200", 747=>x"b000", 748=>x"ae00",
---- 749=>x"af00", 750=>x"b000", 751=>x"b000", 752=>x"af00",
---- 753=>x"b000", 754=>x"af00", 755=>x"b000", 756=>x"ae00",
---- 757=>x"b000", 758=>x"af00", 759=>x"af00", 760=>x"ac00",
---- 761=>x"af00", 762=>x"ad00", 763=>x"af00", 764=>x"ad00",
---- 765=>x"ae00", 766=>x"ac00", 767=>x"af00", 768=>x"ac00",
---- 769=>x"ad00", 770=>x"ac00", 771=>x"ae00", 772=>x"ad00",
---- 773=>x"ac00", 774=>x"ad00", 775=>x"ad00", 776=>x"ab00",
---- 777=>x"ae00", 778=>x"ac00", 779=>x"ac00", 780=>x"ab00",
---- 781=>x"ad00", 782=>x"ad00", 783=>x"ad00", 784=>x"ab00",
---- 785=>x"ad00", 786=>x"ac00", 787=>x"ae00", 788=>x"aa00",
---- 789=>x"ac00", 790=>x"ab00", 791=>x"aa00", 792=>x"ab00",
---- 793=>x"ab00", 794=>x"aa00", 795=>x"a900", 796=>x"aa00",
---- 797=>x"a900", 798=>x"ac00", 799=>x"aa00", 800=>x"aa00",
---- 801=>x"a900", 802=>x"ad00", 803=>x"ad00", 804=>x"a800",
---- 805=>x"aa00", 806=>x"a900", 807=>x"ac00", 808=>x"a700",
---- 809=>x"a800", 810=>x"5400", 811=>x"aa00", 812=>x"a800",
---- 813=>x"a900", 814=>x"ab00", 815=>x"aa00", 816=>x"5600",
---- 817=>x"ad00", 818=>x"ad00", 819=>x"ab00", 820=>x"ac00",
---- 821=>x"ae00", 822=>x"ae00", 823=>x"ad00", 824=>x"ab00",
---- 825=>x"b100", 826=>x"af00", 827=>x"ad00", 828=>x"ae00",
---- 829=>x"b100", 830=>x"b000", 831=>x"af00", 832=>x"ae00",
---- 833=>x"b100", 834=>x"b100", 835=>x"b000", 836=>x"af00",
---- 837=>x"b300", 838=>x"b000", 839=>x"af00", 840=>x"ae00",
---- 841=>x"b200", 842=>x"b200", 843=>x"b200", 844=>x"b000",
---- 845=>x"af00", 846=>x"b000", 847=>x"b000", 848=>x"ad00",
---- 849=>x"b100", 850=>x"b100", 851=>x"ae00", 852=>x"ae00",
---- 853=>x"b300", 854=>x"b300", 855=>x"b000", 856=>x"b000",
---- 857=>x"b500", 858=>x"b400", 859=>x"b200", 860=>x"b000",
---- 861=>x"b200", 862=>x"b100", 863=>x"b000", 864=>x"af00",
---- 865=>x"b300", 866=>x"b100", 867=>x"b300", 868=>x"af00",
---- 869=>x"b400", 870=>x"b300", 871=>x"b200", 872=>x"b300",
---- 873=>x"b500", 874=>x"b300", 875=>x"b100", 876=>x"af00",
---- 877=>x"b200", 878=>x"b300", 879=>x"b100", 880=>x"b000",
---- 881=>x"b100", 882=>x"b100", 883=>x"b100", 884=>x"af00",
---- 885=>x"b000", 886=>x"ad00", 887=>x"ac00", 888=>x"b000",
---- 889=>x"b300", 890=>x"b000", 891=>x"af00", 892=>x"af00",
---- 893=>x"b000", 894=>x"b100", 895=>x"b100", 896=>x"ae00",
---- 897=>x"4d00", 898=>x"b200", 899=>x"b100", 900=>x"ae00",
---- 901=>x"b100", 902=>x"b200", 903=>x"b100", 904=>x"ac00",
---- 905=>x"b000", 906=>x"b100", 907=>x"b100", 908=>x"ae00",
---- 909=>x"b100", 910=>x"b100", 911=>x"b100", 912=>x"ad00",
---- 913=>x"b100", 914=>x"b000", 915=>x"af00", 916=>x"aa00",
---- 917=>x"b100", 918=>x"af00", 919=>x"ad00", 920=>x"a900",
---- 921=>x"af00", 922=>x"b000", 923=>x"b000", 924=>x"aa00",
---- 925=>x"ac00", 926=>x"af00", 927=>x"af00", 928=>x"a800",
---- 929=>x"ab00", 930=>x"ae00", 931=>x"ae00", 932=>x"a700",
---- 933=>x"ad00", 934=>x"ae00", 935=>x"af00", 936=>x"a700",
---- 937=>x"ac00", 938=>x"ad00", 939=>x"af00", 940=>x"a600",
---- 941=>x"ab00", 942=>x"ae00", 943=>x"b100", 944=>x"a700",
---- 945=>x"ac00", 946=>x"b000", 947=>x"af00", 948=>x"a500",
---- 949=>x"ab00", 950=>x"b000", 951=>x"b000", 952=>x"a600",
---- 953=>x"ae00", 954=>x"b100", 955=>x"b100", 956=>x"a700",
---- 957=>x"ad00", 958=>x"b000", 959=>x"b100", 960=>x"a800",
---- 961=>x"ad00", 962=>x"b100", 963=>x"b400", 964=>x"a800",
---- 965=>x"ac00", 966=>x"b000", 967=>x"b200", 968=>x"a600",
---- 969=>x"ab00", 970=>x"b000", 971=>x"b000", 972=>x"a700",
---- 973=>x"ad00", 974=>x"ad00", 975=>x"af00", 976=>x"a600",
---- 977=>x"ad00", 978=>x"af00", 979=>x"b100", 980=>x"a500",
---- 981=>x"ae00", 982=>x"b200", 983=>x"b200", 984=>x"a300",
---- 985=>x"ab00", 986=>x"b000", 987=>x"b200", 988=>x"a500",
---- 989=>x"ad00", 990=>x"b000", 991=>x"b300", 992=>x"a400",
---- 993=>x"ac00", 994=>x"b000", 995=>x"b300", 996=>x"a500",
---- 997=>x"ae00", 998=>x"4d00", 999=>x"b300", 1000=>x"a500",
---- 1001=>x"ae00", 1002=>x"b200", 1003=>x"b200", 1004=>x"a400",
---- 1005=>x"ad00", 1006=>x"b300", 1007=>x"b200", 1008=>x"a200",
---- 1009=>x"ad00", 1010=>x"af00", 1011=>x"b000", 1012=>x"a200",
---- 1013=>x"ae00", 1014=>x"b300", 1015=>x"b000", 1016=>x"a300",
---- 1017=>x"ac00", 1018=>x"b200", 1019=>x"b200", 1020=>x"a200",
---- 1021=>x"a900", 1022=>x"b200", 1023=>x"b400"),
----
---- 6 => (0=>x"ab00", 1=>x"ab00", 2=>x"a900", 3=>x"a200", 4=>x"5400",
---- 5=>x"ab00", 6=>x"a900", 7=>x"a300", 8=>x"ab00",
---- 9=>x"ac00", 10=>x"a900", 11=>x"a200", 12=>x"ad00",
---- 13=>x"ab00", 14=>x"a600", 15=>x"a000", 16=>x"ac00",
---- 17=>x"a900", 18=>x"a600", 19=>x"9e00", 20=>x"aa00",
---- 21=>x"a900", 22=>x"a700", 23=>x"9d00", 24=>x"a800",
---- 25=>x"a700", 26=>x"a600", 27=>x"9d00", 28=>x"a700",
---- 29=>x"a500", 30=>x"9f00", 31=>x"9b00", 32=>x"a600",
---- 33=>x"a300", 34=>x"9f00", 35=>x"9b00", 36=>x"a500",
---- 37=>x"a300", 38=>x"9e00", 39=>x"9800", 40=>x"a200",
---- 41=>x"a300", 42=>x"9d00", 43=>x"9a00", 44=>x"9f00",
---- 45=>x"a100", 46=>x"9f00", 47=>x"9a00", 48=>x"9f00",
---- 49=>x"a200", 50=>x"9f00", 51=>x"9900", 52=>x"a000",
---- 53=>x"a100", 54=>x"a000", 55=>x"9900", 56=>x"a000",
---- 57=>x"a200", 58=>x"a100", 59=>x"9c00", 60=>x"a000",
---- 61=>x"a400", 62=>x"a300", 63=>x"a000", 64=>x"a000",
---- 65=>x"a100", 66=>x"a100", 67=>x"9d00", 68=>x"a000",
---- 69=>x"a300", 70=>x"a200", 71=>x"9b00", 72=>x"9f00",
---- 73=>x"a100", 74=>x"a100", 75=>x"9c00", 76=>x"5d00",
---- 77=>x"a100", 78=>x"a000", 79=>x"9a00", 80=>x"a100",
---- 81=>x"a100", 82=>x"9f00", 83=>x"9b00", 84=>x"5f00",
---- 85=>x"a100", 86=>x"a000", 87=>x"9a00", 88=>x"a000",
---- 89=>x"a200", 90=>x"a000", 91=>x"9900", 92=>x"a200",
---- 93=>x"a400", 94=>x"a100", 95=>x"9a00", 96=>x"a400",
---- 97=>x"5d00", 98=>x"a000", 99=>x"9c00", 100=>x"a400",
---- 101=>x"a400", 102=>x"a100", 103=>x"9c00", 104=>x"a500",
---- 105=>x"a400", 106=>x"a200", 107=>x"9b00", 108=>x"a600",
---- 109=>x"a400", 110=>x"a200", 111=>x"9d00", 112=>x"a600",
---- 113=>x"a500", 114=>x"a400", 115=>x"9f00", 116=>x"a500",
---- 117=>x"a400", 118=>x"a000", 119=>x"9c00", 120=>x"a400",
---- 121=>x"a500", 122=>x"a100", 123=>x"9f00", 124=>x"a600",
---- 125=>x"a500", 126=>x"a300", 127=>x"9d00", 128=>x"a600",
---- 129=>x"a600", 130=>x"a400", 131=>x"9d00", 132=>x"a300",
---- 133=>x"a300", 134=>x"a200", 135=>x"9b00", 136=>x"a300",
---- 137=>x"a300", 138=>x"a100", 139=>x"9a00", 140=>x"a600",
---- 141=>x"a500", 142=>x"a000", 143=>x"9b00", 144=>x"a200",
---- 145=>x"a200", 146=>x"a000", 147=>x"9a00", 148=>x"a500",
---- 149=>x"a300", 150=>x"a000", 151=>x"9900", 152=>x"a400",
---- 153=>x"a300", 154=>x"a000", 155=>x"9900", 156=>x"a300",
---- 157=>x"a100", 158=>x"a000", 159=>x"9c00", 160=>x"a400",
---- 161=>x"a300", 162=>x"5f00", 163=>x"9a00", 164=>x"a600",
---- 165=>x"a300", 166=>x"9f00", 167=>x"9a00", 168=>x"a600",
---- 169=>x"a200", 170=>x"9d00", 171=>x"9800", 172=>x"a600",
---- 173=>x"a500", 174=>x"9e00", 175=>x"9800", 176=>x"a800",
---- 177=>x"a500", 178=>x"9e00", 179=>x"9800", 180=>x"a700",
---- 181=>x"a400", 182=>x"9f00", 183=>x"9800", 184=>x"a400",
---- 185=>x"a300", 186=>x"a000", 187=>x"9a00", 188=>x"a600",
---- 189=>x"a200", 190=>x"9f00", 191=>x"9b00", 192=>x"a300",
---- 193=>x"a400", 194=>x"9e00", 195=>x"9a00", 196=>x"a200",
---- 197=>x"a200", 198=>x"a000", 199=>x"9900", 200=>x"a600",
---- 201=>x"a300", 202=>x"a100", 203=>x"9800", 204=>x"a600",
---- 205=>x"a300", 206=>x"a000", 207=>x"9a00", 208=>x"a400",
---- 209=>x"a300", 210=>x"9f00", 211=>x"6500", 212=>x"a000",
---- 213=>x"a200", 214=>x"9f00", 215=>x"9a00", 216=>x"a300",
---- 217=>x"a300", 218=>x"a100", 219=>x"9c00", 220=>x"a200",
---- 221=>x"a400", 222=>x"a400", 223=>x"9b00", 224=>x"a300",
---- 225=>x"a500", 226=>x"a400", 227=>x"9d00", 228=>x"a300",
---- 229=>x"a300", 230=>x"a400", 231=>x"9b00", 232=>x"a300",
---- 233=>x"a200", 234=>x"a100", 235=>x"9900", 236=>x"a200",
---- 237=>x"a400", 238=>x"a100", 239=>x"9a00", 240=>x"a400",
---- 241=>x"a500", 242=>x"a200", 243=>x"9a00", 244=>x"a300",
---- 245=>x"a200", 246=>x"a000", 247=>x"9c00", 248=>x"a400",
---- 249=>x"a400", 250=>x"a100", 251=>x"9a00", 252=>x"a600",
---- 253=>x"a700", 254=>x"a000", 255=>x"9900", 256=>x"a700",
---- 257=>x"a700", 258=>x"a100", 259=>x"9b00", 260=>x"a500",
---- 261=>x"a500", 262=>x"a400", 263=>x"9e00", 264=>x"a700",
---- 265=>x"a700", 266=>x"a700", 267=>x"9e00", 268=>x"a800",
---- 269=>x"aa00", 270=>x"a600", 271=>x"9e00", 272=>x"a800",
---- 273=>x"a800", 274=>x"a500", 275=>x"a100", 276=>x"a900",
---- 277=>x"a900", 278=>x"aa00", 279=>x"a000", 280=>x"ab00",
---- 281=>x"ac00", 282=>x"aa00", 283=>x"a300", 284=>x"ab00",
---- 285=>x"ad00", 286=>x"aa00", 287=>x"a300", 288=>x"ae00",
---- 289=>x"af00", 290=>x"ac00", 291=>x"a600", 292=>x"ad00",
---- 293=>x"ad00", 294=>x"ac00", 295=>x"a600", 296=>x"ad00",
---- 297=>x"af00", 298=>x"aa00", 299=>x"a500", 300=>x"ab00",
---- 301=>x"ae00", 302=>x"ab00", 303=>x"a500", 304=>x"ae00",
---- 305=>x"b000", 306=>x"ab00", 307=>x"a500", 308=>x"ac00",
---- 309=>x"ae00", 310=>x"aa00", 311=>x"a400", 312=>x"5300",
---- 313=>x"ad00", 314=>x"ac00", 315=>x"a300", 316=>x"aa00",
---- 317=>x"ab00", 318=>x"a900", 319=>x"a400", 320=>x"aa00",
---- 321=>x"ab00", 322=>x"a700", 323=>x"a300", 324=>x"ac00",
---- 325=>x"ac00", 326=>x"aa00", 327=>x"a400", 328=>x"ad00",
---- 329=>x"ab00", 330=>x"ab00", 331=>x"a500", 332=>x"ad00",
---- 333=>x"ab00", 334=>x"aa00", 335=>x"a600", 336=>x"ad00",
---- 337=>x"ad00", 338=>x"a900", 339=>x"a400", 340=>x"ab00",
---- 341=>x"ab00", 342=>x"a800", 343=>x"a300", 344=>x"aa00",
---- 345=>x"ab00", 346=>x"aa00", 347=>x"a700", 348=>x"ae00",
---- 349=>x"ad00", 350=>x"ab00", 351=>x"a800", 352=>x"ad00",
---- 353=>x"ac00", 354=>x"ab00", 355=>x"a600", 356=>x"ac00",
---- 357=>x"ad00", 358=>x"ac00", 359=>x"a500", 360=>x"ae00",
---- 361=>x"ae00", 362=>x"ac00", 363=>x"a700", 364=>x"ac00",
---- 365=>x"ad00", 366=>x"ad00", 367=>x"a600", 368=>x"ae00",
---- 369=>x"ad00", 370=>x"ad00", 371=>x"a600", 372=>x"ad00",
---- 373=>x"ac00", 374=>x"aa00", 375=>x"a700", 376=>x"ac00",
---- 377=>x"ac00", 378=>x"ac00", 379=>x"a600", 380=>x"ac00",
---- 381=>x"ac00", 382=>x"ab00", 383=>x"a700", 384=>x"aa00",
---- 385=>x"aa00", 386=>x"aa00", 387=>x"a600", 388=>x"ab00",
---- 389=>x"ab00", 390=>x"ab00", 391=>x"a700", 392=>x"ab00",
---- 393=>x"ac00", 394=>x"ab00", 395=>x"a800", 396=>x"ac00",
---- 397=>x"ab00", 398=>x"aa00", 399=>x"a600", 400=>x"aa00",
---- 401=>x"ab00", 402=>x"ad00", 403=>x"a800", 404=>x"ac00",
---- 405=>x"ab00", 406=>x"ae00", 407=>x"a500", 408=>x"ae00",
---- 409=>x"ad00", 410=>x"ac00", 411=>x"a500", 412=>x"ae00",
---- 413=>x"ad00", 414=>x"ab00", 415=>x"a800", 416=>x"af00",
---- 417=>x"b100", 418=>x"ae00", 419=>x"a900", 420=>x"ae00",
---- 421=>x"ae00", 422=>x"ae00", 423=>x"aa00", 424=>x"af00",
---- 425=>x"ae00", 426=>x"ac00", 427=>x"a800", 428=>x"ae00",
---- 429=>x"ae00", 430=>x"ad00", 431=>x"a900", 432=>x"af00",
---- 433=>x"ae00", 434=>x"af00", 435=>x"aa00", 436=>x"ac00",
---- 437=>x"ae00", 438=>x"ae00", 439=>x"a800", 440=>x"ad00",
---- 441=>x"ac00", 442=>x"ac00", 443=>x"a800", 444=>x"ae00",
---- 445=>x"ad00", 446=>x"ad00", 447=>x"a700", 448=>x"ae00",
---- 449=>x"ad00", 450=>x"ad00", 451=>x"aa00", 452=>x"b000",
---- 453=>x"ad00", 454=>x"ad00", 455=>x"ad00", 456=>x"ae00",
---- 457=>x"ae00", 458=>x"ad00", 459=>x"ab00", 460=>x"ad00",
---- 461=>x"b000", 462=>x"ae00", 463=>x"aa00", 464=>x"af00",
---- 465=>x"5100", 466=>x"af00", 467=>x"ab00", 468=>x"b000",
---- 469=>x"ad00", 470=>x"ad00", 471=>x"aa00", 472=>x"4e00",
---- 473=>x"ae00", 474=>x"ac00", 475=>x"a700", 476=>x"b100",
---- 477=>x"b000", 478=>x"af00", 479=>x"ab00", 480=>x"b100",
---- 481=>x"af00", 482=>x"ad00", 483=>x"ab00", 484=>x"af00",
---- 485=>x"b000", 486=>x"b100", 487=>x"ac00", 488=>x"b100",
---- 489=>x"af00", 490=>x"ae00", 491=>x"aa00", 492=>x"b100",
---- 493=>x"b000", 494=>x"ad00", 495=>x"ab00", 496=>x"b100",
---- 497=>x"b100", 498=>x"b100", 499=>x"ac00", 500=>x"b100",
---- 501=>x"b400", 502=>x"b000", 503=>x"ab00", 504=>x"b000",
---- 505=>x"b200", 506=>x"b200", 507=>x"ac00", 508=>x"b000",
---- 509=>x"b100", 510=>x"b300", 511=>x"ae00", 512=>x"b000",
---- 513=>x"af00", 514=>x"af00", 515=>x"aa00", 516=>x"b100",
---- 517=>x"b100", 518=>x"b000", 519=>x"ab00", 520=>x"b300",
---- 521=>x"b000", 522=>x"b000", 523=>x"aa00", 524=>x"b100",
---- 525=>x"b000", 526=>x"b000", 527=>x"aa00", 528=>x"b100",
---- 529=>x"b000", 530=>x"b100", 531=>x"aa00", 532=>x"b200",
---- 533=>x"b300", 534=>x"b400", 535=>x"b000", 536=>x"b300",
---- 537=>x"b400", 538=>x"b400", 539=>x"ae00", 540=>x"4900",
---- 541=>x"b400", 542=>x"b200", 543=>x"ae00", 544=>x"b500",
---- 545=>x"b300", 546=>x"b300", 547=>x"af00", 548=>x"b500",
---- 549=>x"b400", 550=>x"b400", 551=>x"4f00", 552=>x"b500",
---- 553=>x"b600", 554=>x"b500", 555=>x"b100", 556=>x"b800",
---- 557=>x"b700", 558=>x"b700", 559=>x"b100", 560=>x"b700",
---- 561=>x"b700", 562=>x"b900", 563=>x"b000", 564=>x"b800",
---- 565=>x"b800", 566=>x"b500", 567=>x"b200", 568=>x"b500",
---- 569=>x"b700", 570=>x"b700", 571=>x"b400", 572=>x"b700",
---- 573=>x"b600", 574=>x"b700", 575=>x"b300", 576=>x"b700",
---- 577=>x"b600", 578=>x"b600", 579=>x"b200", 580=>x"b600",
---- 581=>x"b600", 582=>x"b500", 583=>x"b000", 584=>x"b400",
---- 585=>x"b600", 586=>x"b600", 587=>x"b200", 588=>x"b300",
---- 589=>x"b700", 590=>x"b600", 591=>x"b100", 592=>x"b600",
---- 593=>x"b600", 594=>x"b400", 595=>x"af00", 596=>x"b500",
---- 597=>x"b300", 598=>x"b400", 599=>x"b000", 600=>x"4d00",
---- 601=>x"b100", 602=>x"b100", 603=>x"ae00", 604=>x"af00",
---- 605=>x"b200", 606=>x"b000", 607=>x"ad00", 608=>x"af00",
---- 609=>x"af00", 610=>x"b200", 611=>x"ac00", 612=>x"b000",
---- 613=>x"b300", 614=>x"b100", 615=>x"ac00", 616=>x"ad00",
---- 617=>x"b000", 618=>x"b000", 619=>x"ab00", 620=>x"ac00",
---- 621=>x"b000", 622=>x"b100", 623=>x"ac00", 624=>x"ae00",
---- 625=>x"b000", 626=>x"b200", 627=>x"ae00", 628=>x"b000",
---- 629=>x"b200", 630=>x"b400", 631=>x"ad00", 632=>x"b000",
---- 633=>x"b100", 634=>x"b500", 635=>x"b000", 636=>x"4f00",
---- 637=>x"b200", 638=>x"b400", 639=>x"af00", 640=>x"b100",
---- 641=>x"b200", 642=>x"b300", 643=>x"af00", 644=>x"af00",
---- 645=>x"b100", 646=>x"b300", 647=>x"b100", 648=>x"5000",
---- 649=>x"b100", 650=>x"b400", 651=>x"af00", 652=>x"b000",
---- 653=>x"b200", 654=>x"b300", 655=>x"b000", 656=>x"ae00",
---- 657=>x"b100", 658=>x"b400", 659=>x"b300", 660=>x"af00",
---- 661=>x"b000", 662=>x"b400", 663=>x"b300", 664=>x"ad00",
---- 665=>x"b100", 666=>x"b100", 667=>x"b200", 668=>x"b000",
---- 669=>x"b300", 670=>x"b600", 671=>x"b200", 672=>x"af00",
---- 673=>x"b400", 674=>x"b200", 675=>x"b000", 676=>x"af00",
---- 677=>x"b300", 678=>x"b600", 679=>x"b100", 680=>x"ae00",
---- 681=>x"b000", 682=>x"b400", 683=>x"b300", 684=>x"b000",
---- 685=>x"b100", 686=>x"b400", 687=>x"b200", 688=>x"b100",
---- 689=>x"b300", 690=>x"b600", 691=>x"b200", 692=>x"b000",
---- 693=>x"b400", 694=>x"b500", 695=>x"b300", 696=>x"b100",
---- 697=>x"b500", 698=>x"b500", 699=>x"b300", 700=>x"b300",
---- 701=>x"b300", 702=>x"b200", 703=>x"b300", 704=>x"b200",
---- 705=>x"b300", 706=>x"b500", 707=>x"4c00", 708=>x"b300",
---- 709=>x"b600", 710=>x"b600", 711=>x"b300", 712=>x"b500",
---- 713=>x"b600", 714=>x"b600", 715=>x"b200", 716=>x"b200",
---- 717=>x"b400", 718=>x"b400", 719=>x"b000", 720=>x"b600",
---- 721=>x"b600", 722=>x"b700", 723=>x"b300", 724=>x"b400",
---- 725=>x"b400", 726=>x"b600", 727=>x"4b00", 728=>x"b300",
---- 729=>x"b500", 730=>x"b500", 731=>x"b300", 732=>x"b300",
---- 733=>x"b600", 734=>x"b600", 735=>x"b200", 736=>x"b200",
---- 737=>x"b400", 738=>x"b500", 739=>x"b200", 740=>x"b100",
---- 741=>x"b300", 742=>x"b500", 743=>x"b200", 744=>x"b000",
---- 745=>x"b300", 746=>x"b500", 747=>x"b000", 748=>x"b000",
---- 749=>x"b200", 750=>x"b300", 751=>x"b200", 752=>x"4e00",
---- 753=>x"b100", 754=>x"b100", 755=>x"b200", 756=>x"b100",
---- 757=>x"b000", 758=>x"b300", 759=>x"b200", 760=>x"b300",
---- 761=>x"b100", 762=>x"b300", 763=>x"b200", 764=>x"b000",
---- 765=>x"b200", 766=>x"b300", 767=>x"b200", 768=>x"b100",
---- 769=>x"b200", 770=>x"4d00", 771=>x"b000", 772=>x"b000",
---- 773=>x"b000", 774=>x"b400", 775=>x"b200", 776=>x"af00",
---- 777=>x"af00", 778=>x"b100", 779=>x"af00", 780=>x"ad00",
---- 781=>x"ac00", 782=>x"ae00", 783=>x"b000", 784=>x"ad00",
---- 785=>x"ae00", 786=>x"af00", 787=>x"af00", 788=>x"ab00",
---- 789=>x"ad00", 790=>x"af00", 791=>x"ad00", 792=>x"ab00",
---- 793=>x"ac00", 794=>x"ae00", 795=>x"ad00", 796=>x"ab00",
---- 797=>x"ab00", 798=>x"ac00", 799=>x"b200", 800=>x"ac00",
---- 801=>x"ab00", 802=>x"b000", 803=>x"bb00", 804=>x"ac00",
---- 805=>x"a800", 806=>x"b000", 807=>x"b100", 808=>x"ab00",
---- 809=>x"ab00", 810=>x"ab00", 811=>x"ac00", 812=>x"ab00",
---- 813=>x"ae00", 814=>x"ae00", 815=>x"ae00", 816=>x"ac00",
---- 817=>x"ac00", 818=>x"af00", 819=>x"af00", 820=>x"ad00",
---- 821=>x"ac00", 822=>x"b100", 823=>x"b000", 824=>x"ad00",
---- 825=>x"af00", 826=>x"b100", 827=>x"ae00", 828=>x"af00",
---- 829=>x"ae00", 830=>x"4d00", 831=>x"b000", 832=>x"ae00",
---- 833=>x"b100", 834=>x"b400", 835=>x"b100", 836=>x"b000",
---- 837=>x"b300", 838=>x"b400", 839=>x"b000", 840=>x"b100",
---- 841=>x"b200", 842=>x"b300", 843=>x"b000", 844=>x"b200",
---- 845=>x"b100", 846=>x"b300", 847=>x"b100", 848=>x"af00",
---- 849=>x"b200", 850=>x"b200", 851=>x"b200", 852=>x"af00",
---- 853=>x"b300", 854=>x"b300", 855=>x"b200", 856=>x"b200",
---- 857=>x"b300", 858=>x"b500", 859=>x"b200", 860=>x"b100",
---- 861=>x"b200", 862=>x"b600", 863=>x"b500", 864=>x"b300",
---- 865=>x"b100", 866=>x"b500", 867=>x"b600", 868=>x"b200",
---- 869=>x"b400", 870=>x"b600", 871=>x"b300", 872=>x"b300",
---- 873=>x"4b00", 874=>x"b500", 875=>x"b400", 876=>x"b300",
---- 877=>x"b300", 878=>x"b400", 879=>x"b400", 880=>x"b100",
---- 881=>x"b200", 882=>x"b100", 883=>x"b200", 884=>x"ac00",
---- 885=>x"a900", 886=>x"a900", 887=>x"ad00", 888=>x"ad00",
---- 889=>x"ab00", 890=>x"af00", 891=>x"b100", 892=>x"b200",
---- 893=>x"b100", 894=>x"b300", 895=>x"b200", 896=>x"b200",
---- 897=>x"b200", 898=>x"b500", 899=>x"b300", 900=>x"b200",
---- 901=>x"b200", 902=>x"b300", 903=>x"b300", 904=>x"b200",
---- 905=>x"b100", 906=>x"b200", 907=>x"b300", 908=>x"b000",
---- 909=>x"b100", 910=>x"b100", 911=>x"b200", 912=>x"b000",
---- 913=>x"b100", 914=>x"b200", 915=>x"b200", 916=>x"b100",
---- 917=>x"b100", 918=>x"b200", 919=>x"b300", 920=>x"b000",
---- 921=>x"b000", 922=>x"b100", 923=>x"b100", 924=>x"b000",
---- 925=>x"b200", 926=>x"b300", 927=>x"b300", 928=>x"b000",
---- 929=>x"b200", 930=>x"b300", 931=>x"b500", 932=>x"b200",
---- 933=>x"b000", 934=>x"b100", 935=>x"b200", 936=>x"b100",
---- 937=>x"af00", 938=>x"b100", 939=>x"b500", 940=>x"b000",
---- 941=>x"b000", 942=>x"b200", 943=>x"b500", 944=>x"af00",
---- 945=>x"ae00", 946=>x"b300", 947=>x"b600", 948=>x"ac00",
---- 949=>x"ae00", 950=>x"b400", 951=>x"b700", 952=>x"ae00",
---- 953=>x"ad00", 954=>x"b300", 955=>x"b700", 956=>x"b100",
---- 957=>x"b000", 958=>x"b500", 959=>x"ba00", 960=>x"b100",
---- 961=>x"b000", 962=>x"b500", 963=>x"b900", 964=>x"b200",
---- 965=>x"b300", 966=>x"b600", 967=>x"b800", 968=>x"b200",
---- 969=>x"b500", 970=>x"b700", 971=>x"b800", 972=>x"b100",
---- 973=>x"b300", 974=>x"b600", 975=>x"b800", 976=>x"b200",
---- 977=>x"b300", 978=>x"b600", 979=>x"b700", 980=>x"b400",
---- 981=>x"b400", 982=>x"b600", 983=>x"b700", 984=>x"b500",
---- 985=>x"b400", 986=>x"4800", 987=>x"b900", 988=>x"b400",
---- 989=>x"b400", 990=>x"b600", 991=>x"b900", 992=>x"b400",
---- 993=>x"b500", 994=>x"b500", 995=>x"b800", 996=>x"b500",
---- 997=>x"b500", 998=>x"b900", 999=>x"b900", 1000=>x"b500",
---- 1001=>x"b600", 1002=>x"ba00", 1003=>x"bb00", 1004=>x"b600",
---- 1005=>x"b400", 1006=>x"b700", 1007=>x"b800", 1008=>x"b300",
---- 1009=>x"b200", 1010=>x"b500", 1011=>x"b500", 1012=>x"b300",
---- 1013=>x"b300", 1014=>x"b400", 1015=>x"b700", 1016=>x"b400",
---- 1017=>x"b400", 1018=>x"b400", 1019=>x"b700", 1020=>x"b400",
---- 1021=>x"b400", 1022=>x"b500", 1023=>x"b600"),
----
---- 7 => (0=>x"9700", 1=>x"9600", 2=>x"8200", 3=>x"7300", 4=>x"9700",
---- 5=>x"9700", 6=>x"8300", 7=>x"7200", 8=>x"9800",
---- 9=>x"9500", 10=>x"8000", 11=>x"7000", 12=>x"9700",
---- 13=>x"8b00", 14=>x"7c00", 15=>x"7100", 16=>x"9500",
---- 17=>x"8b00", 18=>x"7d00", 19=>x"7300", 20=>x"9100",
---- 21=>x"8800", 22=>x"8000", 23=>x"7000", 24=>x"8e00",
---- 25=>x"8900", 26=>x"7d00", 27=>x"6c00", 28=>x"9300",
---- 29=>x"8800", 30=>x"7d00", 31=>x"7200", 32=>x"9000",
---- 33=>x"8800", 34=>x"7c00", 35=>x"6d00", 36=>x"9000",
---- 37=>x"8a00", 38=>x"7f00", 39=>x"6f00", 40=>x"9100",
---- 41=>x"8b00", 42=>x"8400", 43=>x"7900", 44=>x"9300",
---- 45=>x"8900", 46=>x"8200", 47=>x"7100", 48=>x"9500",
---- 49=>x"8b00", 50=>x"8000", 51=>x"7200", 52=>x"9400",
---- 53=>x"8b00", 54=>x"7b00", 55=>x"6c00", 56=>x"9400",
---- 57=>x"8a00", 58=>x"7b00", 59=>x"6d00", 60=>x"9400",
---- 61=>x"8900", 62=>x"7e00", 63=>x"6e00", 64=>x"9600",
---- 65=>x"8c00", 66=>x"8000", 67=>x"6f00", 68=>x"9300",
---- 69=>x"8800", 70=>x"7c00", 71=>x"6c00", 72=>x"9200",
---- 73=>x"8700", 74=>x"7f00", 75=>x"6d00", 76=>x"9100",
---- 77=>x"8900", 78=>x"7f00", 79=>x"6d00", 80=>x"9400",
---- 81=>x"8700", 82=>x"7b00", 83=>x"6900", 84=>x"9100",
---- 85=>x"8900", 86=>x"7b00", 87=>x"6900", 88=>x"9400",
---- 89=>x"8900", 90=>x"7c00", 91=>x"6a00", 92=>x"9500",
---- 93=>x"8b00", 94=>x"7d00", 95=>x"6b00", 96=>x"9500",
---- 97=>x"8a00", 98=>x"8200", 99=>x"7000", 100=>x"9500",
---- 101=>x"8900", 102=>x"8100", 103=>x"6c00", 104=>x"9300",
---- 105=>x"8a00", 106=>x"7f00", 107=>x"6c00", 108=>x"9100",
---- 109=>x"8d00", 110=>x"7e00", 111=>x"6c00", 112=>x"9500",
---- 113=>x"8b00", 114=>x"8000", 115=>x"6c00", 116=>x"6900",
---- 117=>x"8b00", 118=>x"7e00", 119=>x"6800", 120=>x"9600",
---- 121=>x"8d00", 122=>x"8000", 123=>x"6b00", 124=>x"9600",
---- 125=>x"8b00", 126=>x"8000", 127=>x"6e00", 128=>x"9600",
---- 129=>x"8b00", 130=>x"7d00", 131=>x"6a00", 132=>x"9400",
---- 133=>x"8b00", 134=>x"7e00", 135=>x"6d00", 136=>x"9100",
---- 137=>x"8800", 138=>x"7f00", 139=>x"6b00", 140=>x"8f00",
---- 141=>x"8800", 142=>x"7d00", 143=>x"6b00", 144=>x"9100",
---- 145=>x"8900", 146=>x"7c00", 147=>x"6a00", 148=>x"9200",
---- 149=>x"8700", 150=>x"8200", 151=>x"6c00", 152=>x"9300",
---- 153=>x"8900", 154=>x"7a00", 155=>x"6700", 156=>x"9400",
---- 157=>x"8a00", 158=>x"7b00", 159=>x"6b00", 160=>x"9300",
---- 161=>x"8900", 162=>x"7900", 163=>x"6800", 164=>x"9100",
---- 165=>x"8600", 166=>x"7900", 167=>x"6700", 168=>x"8f00",
---- 169=>x"8600", 170=>x"7500", 171=>x"6b00", 172=>x"9000",
---- 173=>x"8600", 174=>x"7900", 175=>x"6a00", 176=>x"9000",
---- 177=>x"8300", 178=>x"7c00", 179=>x"6b00", 180=>x"9000",
---- 181=>x"8400", 182=>x"7700", 183=>x"6a00", 184=>x"9000",
---- 185=>x"8500", 186=>x"7900", 187=>x"6800", 188=>x"9100",
---- 189=>x"8400", 190=>x"7600", 191=>x"6700", 192=>x"9200",
---- 193=>x"8800", 194=>x"7800", 195=>x"6c00", 196=>x"8e00",
---- 197=>x"8500", 198=>x"7a00", 199=>x"6800", 200=>x"9000",
---- 201=>x"8600", 202=>x"7800", 203=>x"6a00", 204=>x"9100",
---- 205=>x"8500", 206=>x"7a00", 207=>x"6b00", 208=>x"9200",
---- 209=>x"8600", 210=>x"7a00", 211=>x"6800", 212=>x"9200",
---- 213=>x"8900", 214=>x"7900", 215=>x"6900", 216=>x"6f00",
---- 217=>x"8800", 218=>x"7900", 219=>x"6a00", 220=>x"9300",
---- 221=>x"8800", 222=>x"7b00", 223=>x"6a00", 224=>x"9200",
---- 225=>x"8700", 226=>x"7800", 227=>x"6c00", 228=>x"9200",
---- 229=>x"8900", 230=>x"7d00", 231=>x"7000", 232=>x"9300",
---- 233=>x"8600", 234=>x"7b00", 235=>x"6c00", 236=>x"9100",
---- 237=>x"8800", 238=>x"7800", 239=>x"6800", 240=>x"9100",
---- 241=>x"8600", 242=>x"7a00", 243=>x"6a00", 244=>x"9300",
---- 245=>x"8600", 246=>x"7b00", 247=>x"6500", 248=>x"9300",
---- 249=>x"8600", 250=>x"7700", 251=>x"6600", 252=>x"9300",
---- 253=>x"8600", 254=>x"7a00", 255=>x"6900", 256=>x"9500",
---- 257=>x"8a00", 258=>x"7700", 259=>x"6800", 260=>x"9600",
---- 261=>x"8b00", 262=>x"7a00", 263=>x"6b00", 264=>x"9800",
---- 265=>x"8d00", 266=>x"7a00", 267=>x"6a00", 268=>x"9600",
---- 269=>x"8c00", 270=>x"7900", 271=>x"6900", 272=>x"9800",
---- 273=>x"8c00", 274=>x"7b00", 275=>x"6e00", 276=>x"9800",
---- 277=>x"8b00", 278=>x"7b00", 279=>x"6f00", 280=>x"9900",
---- 281=>x"8d00", 282=>x"7e00", 283=>x"6c00", 284=>x"6400",
---- 285=>x"8e00", 286=>x"7e00", 287=>x"6900", 288=>x"9b00",
---- 289=>x"8e00", 290=>x"7e00", 291=>x"6a00", 292=>x"9a00",
---- 293=>x"9000", 294=>x"7d00", 295=>x"6e00", 296=>x"9b00",
---- 297=>x"8f00", 298=>x"7c00", 299=>x"6e00", 300=>x"9a00",
---- 301=>x"8d00", 302=>x"7c00", 303=>x"6e00", 304=>x"9800",
---- 305=>x"8d00", 306=>x"7f00", 307=>x"7000", 308=>x"9a00",
---- 309=>x"8e00", 310=>x"8100", 311=>x"6f00", 312=>x"9a00",
---- 313=>x"8f00", 314=>x"7e00", 315=>x"6c00", 316=>x"9b00",
---- 317=>x"8f00", 318=>x"8100", 319=>x"6c00", 320=>x"9a00",
---- 321=>x"8f00", 322=>x"7f00", 323=>x"6c00", 324=>x"9b00",
---- 325=>x"9300", 326=>x"8000", 327=>x"6c00", 328=>x"9a00",
---- 329=>x"9100", 330=>x"8300", 331=>x"6c00", 332=>x"9a00",
---- 333=>x"9200", 334=>x"8300", 335=>x"6d00", 336=>x"9c00",
---- 337=>x"9400", 338=>x"8400", 339=>x"7200", 340=>x"9d00",
---- 341=>x"9400", 342=>x"8600", 343=>x"6d00", 344=>x"9d00",
---- 345=>x"9100", 346=>x"8300", 347=>x"6c00", 348=>x"9f00",
---- 349=>x"9400", 350=>x"8500", 351=>x"6e00", 352=>x"9f00",
---- 353=>x"9400", 354=>x"8300", 355=>x"6f00", 356=>x"9f00",
---- 357=>x"9300", 358=>x"8300", 359=>x"6e00", 360=>x"9e00",
---- 361=>x"9200", 362=>x"8500", 363=>x"7000", 364=>x"9e00",
---- 365=>x"9500", 366=>x"8500", 367=>x"7200", 368=>x"9f00",
---- 369=>x"9400", 370=>x"8700", 371=>x"6e00", 372=>x"a100",
---- 373=>x"9300", 374=>x"8400", 375=>x"6f00", 376=>x"a000",
---- 377=>x"9400", 378=>x"8600", 379=>x"6f00", 380=>x"a000",
---- 381=>x"9400", 382=>x"8500", 383=>x"6f00", 384=>x"9e00",
---- 385=>x"9600", 386=>x"8600", 387=>x"7200", 388=>x"9f00",
---- 389=>x"9400", 390=>x"8700", 391=>x"7100", 392=>x"9e00",
---- 393=>x"9200", 394=>x"8700", 395=>x"7100", 396=>x"9d00",
---- 397=>x"9400", 398=>x"8600", 399=>x"8b00", 400=>x"a000",
---- 401=>x"9500", 402=>x"8b00", 403=>x"7600", 404=>x"9f00",
---- 405=>x"6b00", 406=>x"8800", 407=>x"7600", 408=>x"9f00",
---- 409=>x"9600", 410=>x"8800", 411=>x"7400", 412=>x"9f00",
---- 413=>x"6900", 414=>x"8800", 415=>x"7500", 416=>x"9f00",
---- 417=>x"6b00", 418=>x"8700", 419=>x"7400", 420=>x"9e00",
---- 421=>x"9600", 422=>x"8b00", 423=>x"7400", 424=>x"a000",
---- 425=>x"9600", 426=>x"8900", 427=>x"7700", 428=>x"a100",
---- 429=>x"9500", 430=>x"8900", 431=>x"7800", 432=>x"9f00",
---- 433=>x"9700", 434=>x"8a00", 435=>x"7800", 436=>x"9e00",
---- 437=>x"9800", 438=>x"8900", 439=>x"7400", 440=>x"a100",
---- 441=>x"9500", 442=>x"8a00", 443=>x"7500", 444=>x"a000",
---- 445=>x"9a00", 446=>x"8b00", 447=>x"7600", 448=>x"a100",
---- 449=>x"6600", 450=>x"8c00", 451=>x"7a00", 452=>x"a100",
---- 453=>x"9600", 454=>x"8a00", 455=>x"7900", 456=>x"a200",
---- 457=>x"9700", 458=>x"8900", 459=>x"7700", 460=>x"a000",
---- 461=>x"9600", 462=>x"8a00", 463=>x"7800", 464=>x"a100",
---- 465=>x"9600", 466=>x"8b00", 467=>x"7600", 468=>x"a100",
---- 469=>x"9400", 470=>x"8b00", 471=>x"7700", 472=>x"a100",
---- 473=>x"9900", 474=>x"8e00", 475=>x"7700", 476=>x"a000",
---- 477=>x"9800", 478=>x"8b00", 479=>x"7500", 480=>x"a100",
---- 481=>x"9500", 482=>x"8900", 483=>x"7500", 484=>x"a100",
---- 485=>x"9700", 486=>x"8b00", 487=>x"7600", 488=>x"a300",
---- 489=>x"9900", 490=>x"8b00", 491=>x"7700", 492=>x"a200",
---- 493=>x"9800", 494=>x"8a00", 495=>x"7700", 496=>x"a200",
---- 497=>x"6500", 498=>x"8c00", 499=>x"7500", 500=>x"a300",
---- 501=>x"9800", 502=>x"8e00", 503=>x"7a00", 504=>x"a200",
---- 505=>x"9600", 506=>x"8c00", 507=>x"7a00", 508=>x"a200",
---- 509=>x"9b00", 510=>x"8e00", 511=>x"7a00", 512=>x"a400",
---- 513=>x"9c00", 514=>x"9200", 515=>x"7c00", 516=>x"a300",
---- 517=>x"9a00", 518=>x"8d00", 519=>x"7c00", 520=>x"a000",
---- 521=>x"9700", 522=>x"8e00", 523=>x"7b00", 524=>x"a000",
---- 525=>x"9a00", 526=>x"8c00", 527=>x"7a00", 528=>x"a000",
---- 529=>x"9700", 530=>x"8b00", 531=>x"7800", 532=>x"a100",
---- 533=>x"9700", 534=>x"8b00", 535=>x"7900", 536=>x"a400",
---- 537=>x"9700", 538=>x"8a00", 539=>x"7b00", 540=>x"a500",
---- 541=>x"9600", 542=>x"8900", 543=>x"7b00", 544=>x"a500",
---- 545=>x"9a00", 546=>x"8900", 547=>x"7800", 548=>x"a400",
---- 549=>x"9b00", 550=>x"8a00", 551=>x"7e00", 552=>x"a500",
---- 553=>x"9d00", 554=>x"8e00", 555=>x"7e00", 556=>x"a900",
---- 557=>x"9f00", 558=>x"8e00", 559=>x"7e00", 560=>x"aa00",
---- 561=>x"9f00", 562=>x"8f00", 563=>x"7e00", 564=>x"aa00",
---- 565=>x"9e00", 566=>x"9000", 567=>x"8000", 568=>x"a700",
---- 569=>x"9d00", 570=>x"9000", 571=>x"8200", 572=>x"a800",
---- 573=>x"9f00", 574=>x"8f00", 575=>x"7f00", 576=>x"a800",
---- 577=>x"9f00", 578=>x"9000", 579=>x"8000", 580=>x"a800",
---- 581=>x"9e00", 582=>x"9000", 583=>x"7e00", 584=>x"a600",
---- 585=>x"9e00", 586=>x"8d00", 587=>x"8000", 588=>x"a700",
---- 589=>x"9e00", 590=>x"9100", 591=>x"7f00", 592=>x"a800",
---- 593=>x"9b00", 594=>x"9100", 595=>x"7e00", 596=>x"a700",
---- 597=>x"9900", 598=>x"9200", 599=>x"7f00", 600=>x"a400",
---- 601=>x"9d00", 602=>x"9000", 603=>x"8000", 604=>x"a600",
---- 605=>x"9c00", 606=>x"9000", 607=>x"8100", 608=>x"a400",
---- 609=>x"9900", 610=>x"9100", 611=>x"8100", 612=>x"a300",
---- 613=>x"9a00", 614=>x"9000", 615=>x"7f00", 616=>x"a400",
---- 617=>x"9a00", 618=>x"8f00", 619=>x"7f00", 620=>x"a400",
---- 621=>x"9a00", 622=>x"9000", 623=>x"8000", 624=>x"a500",
---- 625=>x"9d00", 626=>x"9100", 627=>x"7e00", 628=>x"a600",
---- 629=>x"9d00", 630=>x"9100", 631=>x"7f00", 632=>x"a900",
---- 633=>x"9e00", 634=>x"9000", 635=>x"7f00", 636=>x"a800",
---- 637=>x"9d00", 638=>x"9200", 639=>x"7f00", 640=>x"a900",
---- 641=>x"9e00", 642=>x"8f00", 643=>x"7f00", 644=>x"a800",
---- 645=>x"9b00", 646=>x"9000", 647=>x"8300", 648=>x"aa00",
---- 649=>x"9e00", 650=>x"9000", 651=>x"8500", 652=>x"aa00",
---- 653=>x"a000", 654=>x"9100", 655=>x"8300", 656=>x"a900",
---- 657=>x"9e00", 658=>x"9200", 659=>x"8400", 660=>x"ab00",
---- 661=>x"9e00", 662=>x"9200", 663=>x"8400", 664=>x"ab00",
---- 665=>x"a000", 666=>x"9400", 667=>x"8200", 668=>x"ab00",
---- 669=>x"a100", 670=>x"9400", 671=>x"8700", 672=>x"aa00",
---- 673=>x"a000", 674=>x"9400", 675=>x"8400", 676=>x"ab00",
---- 677=>x"a100", 678=>x"9400", 679=>x"8500", 680=>x"aa00",
---- 681=>x"a200", 682=>x"9400", 683=>x"8400", 684=>x"ad00",
---- 685=>x"5c00", 686=>x"9700", 687=>x"8600", 688=>x"ae00",
---- 689=>x"a400", 690=>x"9400", 691=>x"8600", 692=>x"ae00",
---- 693=>x"a400", 694=>x"9700", 695=>x"8400", 696=>x"ad00",
---- 697=>x"a100", 698=>x"9500", 699=>x"8300", 700=>x"ac00",
---- 701=>x"a300", 702=>x"9400", 703=>x"8000", 704=>x"aa00",
---- 705=>x"a100", 706=>x"9200", 707=>x"8100", 708=>x"a800",
---- 709=>x"9f00", 710=>x"9400", 711=>x"8200", 712=>x"a900",
---- 713=>x"5e00", 714=>x"9500", 715=>x"7d00", 716=>x"a900",
---- 717=>x"a800", 718=>x"9b00", 719=>x"8300", 720=>x"aa00",
---- 721=>x"a800", 722=>x"ae00", 723=>x"9900", 724=>x"ac00",
---- 725=>x"a100", 726=>x"9900", 727=>x"8400", 728=>x"ac00",
---- 729=>x"9f00", 730=>x"9300", 731=>x"8000", 732=>x"aa00",
---- 733=>x"a000", 734=>x"9400", 735=>x"8200", 736=>x"ab00",
---- 737=>x"a200", 738=>x"6900", 739=>x"8600", 740=>x"aa00",
---- 741=>x"a300", 742=>x"9800", 743=>x"8500", 744=>x"a900",
---- 745=>x"a000", 746=>x"9500", 747=>x"8400", 748=>x"aa00",
---- 749=>x"a200", 750=>x"9600", 751=>x"7b00", 752=>x"a900",
---- 753=>x"a100", 754=>x"9400", 755=>x"8100", 756=>x"aa00",
---- 757=>x"a200", 758=>x"9400", 759=>x"8500", 760=>x"aa00",
---- 761=>x"a300", 762=>x"9800", 763=>x"8300", 764=>x"ae00",
---- 765=>x"a300", 766=>x"9700", 767=>x"8600", 768=>x"ab00",
---- 769=>x"a300", 770=>x"9400", 771=>x"8400", 772=>x"a800",
---- 773=>x"a000", 774=>x"9200", 775=>x"7f00", 776=>x"a800",
---- 777=>x"9e00", 778=>x"9100", 779=>x"7a00", 780=>x"a800",
---- 781=>x"9d00", 782=>x"8d00", 783=>x"7800", 784=>x"a800",
---- 785=>x"9900", 786=>x"8c00", 787=>x"7b00", 788=>x"a600",
---- 789=>x"9b00", 790=>x"9000", 791=>x"a800", 792=>x"a600",
---- 793=>x"a000", 794=>x"b600", 795=>x"c300", 796=>x"b900",
---- 797=>x"b600", 798=>x"ac00", 799=>x"8600", 800=>x"bd00",
---- 801=>x"a800", 802=>x"9500", 803=>x"8100", 804=>x"a900",
---- 805=>x"a200", 806=>x"9700", 807=>x"8500", 808=>x"a900",
---- 809=>x"a200", 810=>x"9600", 811=>x"7f00", 812=>x"a800",
---- 813=>x"9f00", 814=>x"9300", 815=>x"7d00", 816=>x"a800",
---- 817=>x"a000", 818=>x"8f00", 819=>x"8800", 820=>x"a800",
---- 821=>x"a100", 822=>x"8d00", 823=>x"9800", 824=>x"a700",
---- 825=>x"9e00", 826=>x"8f00", 827=>x"a300", 828=>x"a900",
---- 829=>x"a100", 830=>x"9100", 831=>x"9400", 832=>x"a900",
---- 833=>x"a200", 834=>x"9200", 835=>x"9400", 836=>x"aa00",
---- 837=>x"9e00", 838=>x"9400", 839=>x"9e00", 840=>x"a900",
---- 841=>x"a200", 842=>x"9400", 843=>x"9300", 844=>x"a900",
---- 845=>x"a200", 846=>x"9800", 847=>x"8800", 848=>x"ac00",
---- 849=>x"a400", 850=>x"9a00", 851=>x"8a00", 852=>x"ac00",
---- 853=>x"a500", 854=>x"9b00", 855=>x"8a00", 856=>x"ad00",
---- 857=>x"a600", 858=>x"9c00", 859=>x"8d00", 860=>x"af00",
---- 861=>x"a700", 862=>x"9c00", 863=>x"8800", 864=>x"af00",
---- 865=>x"a600", 866=>x"9c00", 867=>x"8700", 868=>x"ac00",
---- 869=>x"a500", 870=>x"9b00", 871=>x"8900", 872=>x"ad00",
---- 873=>x"a600", 874=>x"9c00", 875=>x"8900", 876=>x"b000",
---- 877=>x"a700", 878=>x"9e00", 879=>x"8c00", 880=>x"ac00",
---- 881=>x"a300", 882=>x"9c00", 883=>x"9200", 884=>x"a800",
---- 885=>x"a000", 886=>x"9900", 887=>x"8f00", 888=>x"aa00",
---- 889=>x"a300", 890=>x"9900", 891=>x"8b00", 892=>x"ac00",
---- 893=>x"a600", 894=>x"9900", 895=>x"9200", 896=>x"ae00",
---- 897=>x"a600", 898=>x"9c00", 899=>x"8d00", 900=>x"b000",
---- 901=>x"a600", 902=>x"9800", 903=>x"8f00", 904=>x"ae00",
---- 905=>x"a800", 906=>x"9500", 907=>x"9800", 908=>x"aa00",
---- 909=>x"a500", 910=>x"9800", 911=>x"9000", 912=>x"ad00",
---- 913=>x"a400", 914=>x"9800", 915=>x"8c00", 916=>x"ad00",
---- 917=>x"a700", 918=>x"9c00", 919=>x"8700", 920=>x"ad00",
---- 921=>x"a700", 922=>x"9d00", 923=>x"8500", 924=>x"ae00",
---- 925=>x"5a00", 926=>x"9e00", 927=>x"8a00", 928=>x"af00",
---- 929=>x"a900", 930=>x"9e00", 931=>x"8e00", 932=>x"af00",
---- 933=>x"a800", 934=>x"9d00", 935=>x"6d00", 936=>x"b100",
---- 937=>x"a600", 938=>x"9e00", 939=>x"9500", 940=>x"b200",
---- 941=>x"ab00", 942=>x"a100", 943=>x"8e00", 944=>x"b300",
---- 945=>x"ac00", 946=>x"a400", 947=>x"8500", 948=>x"b100",
---- 949=>x"aa00", 950=>x"a500", 951=>x"7e00", 952=>x"b100",
---- 953=>x"ab00", 954=>x"a000", 955=>x"7600", 956=>x"b100",
---- 957=>x"ae00", 958=>x"9d00", 959=>x"7700", 960=>x"b300",
---- 961=>x"ac00", 962=>x"9d00", 963=>x"7000", 964=>x"b200",
---- 965=>x"af00", 966=>x"a100", 967=>x"6400", 968=>x"b100",
---- 969=>x"ac00", 970=>x"a400", 971=>x"6100", 972=>x"b200",
---- 973=>x"ab00", 974=>x"a400", 975=>x"6900", 976=>x"b300",
---- 977=>x"ab00", 978=>x"a700", 979=>x"6c00", 980=>x"b100",
---- 981=>x"aa00", 982=>x"a700", 983=>x"7a00", 984=>x"4900",
---- 985=>x"ad00", 986=>x"a800", 987=>x"8700", 988=>x"b500",
---- 989=>x"a800", 990=>x"a600", 991=>x"9000", 992=>x"b300",
---- 993=>x"a900", 994=>x"5900", 995=>x"8f00", 996=>x"b400",
---- 997=>x"ad00", 998=>x"a300", 999=>x"7200", 1000=>x"b600",
---- 1001=>x"ac00", 1002=>x"8100", 1003=>x"4900", 1004=>x"b400",
---- 1005=>x"aa00", 1006=>x"8700", 1007=>x"6500", 1008=>x"b200",
---- 1009=>x"ae00", 1010=>x"9600", 1011=>x"8000", 1012=>x"b300",
---- 1013=>x"ac00", 1014=>x"8800", 1015=>x"7500", 1016=>x"b400",
---- 1017=>x"ad00", 1018=>x"7700", 1019=>x"5a00", 1020=>x"b200",
---- 1021=>x"b200", 1022=>x"7800", 1023=>x"5500"),
----
---- 8 => (0=>x"6300", 1=>x"5d00", 2=>x"5b00", 3=>x"6400", 4=>x"6300",
---- 5=>x"5e00", 6=>x"5b00", 7=>x"6500", 8=>x"6400",
---- 9=>x"5e00", 10=>x"5c00", 11=>x"6300", 12=>x"6300",
---- 13=>x"5b00", 14=>x"5a00", 15=>x"5e00", 16=>x"6300",
---- 17=>x"5a00", 18=>x"5800", 19=>x"5a00", 20=>x"6000",
---- 21=>x"5b00", 22=>x"5900", 23=>x"5b00", 24=>x"6300",
---- 25=>x"5900", 26=>x"5900", 27=>x"5b00", 28=>x"6400",
---- 29=>x"5a00", 30=>x"5c00", 31=>x"5b00", 32=>x"6100",
---- 33=>x"5900", 34=>x"5700", 35=>x"5b00", 36=>x"6100",
---- 37=>x"5b00", 38=>x"5700", 39=>x"5d00", 40=>x"6600",
---- 41=>x"a300", 42=>x"5700", 43=>x"5d00", 44=>x"6100",
---- 45=>x"5a00", 46=>x"5b00", 47=>x"5f00", 48=>x"6300",
---- 49=>x"5800", 50=>x"5600", 51=>x"5d00", 52=>x"5c00",
---- 53=>x"5800", 54=>x"5200", 55=>x"5600", 56=>x"5f00",
---- 57=>x"5700", 58=>x"5500", 59=>x"5700", 60=>x"6100",
---- 61=>x"5a00", 62=>x"5600", 63=>x"5a00", 64=>x"6100",
---- 65=>x"5a00", 66=>x"5700", 67=>x"5e00", 68=>x"5f00",
---- 69=>x"5800", 70=>x"5a00", 71=>x"5d00", 72=>x"6000",
---- 73=>x"5600", 74=>x"5600", 75=>x"5a00", 76=>x"5b00",
---- 77=>x"5300", 78=>x"5300", 79=>x"5700", 80=>x"5d00",
---- 81=>x"5400", 82=>x"5100", 83=>x"5b00", 84=>x"5d00",
---- 85=>x"5400", 86=>x"5300", 87=>x"5900", 88=>x"5d00",
---- 89=>x"5300", 90=>x"5300", 91=>x"5b00", 92=>x"5e00",
---- 93=>x"5400", 94=>x"5100", 95=>x"5b00", 96=>x"6100",
---- 97=>x"5800", 98=>x"5300", 99=>x"5900", 100=>x"5c00",
---- 101=>x"5600", 102=>x"5500", 103=>x"5900", 104=>x"5e00",
---- 105=>x"5200", 106=>x"ae00", 107=>x"5700", 108=>x"5c00",
---- 109=>x"5100", 110=>x"5500", 111=>x"5800", 112=>x"5900",
---- 113=>x"4f00", 114=>x"5000", 115=>x"5600", 116=>x"5900",
---- 117=>x"4c00", 118=>x"4e00", 119=>x"5300", 120=>x"a600",
---- 121=>x"5100", 122=>x"4e00", 123=>x"5300", 124=>x"5900",
---- 125=>x"5200", 126=>x"4d00", 127=>x"5000", 128=>x"5a00",
---- 129=>x"4c00", 130=>x"4c00", 131=>x"5100", 132=>x"5700",
---- 133=>x"4b00", 134=>x"4900", 135=>x"5100", 136=>x"5900",
---- 137=>x"4e00", 138=>x"4700", 139=>x"5000", 140=>x"5500",
---- 141=>x"4b00", 142=>x"4700", 143=>x"5000", 144=>x"5300",
---- 145=>x"4b00", 146=>x"4800", 147=>x"5000", 148=>x"5300",
---- 149=>x"4b00", 150=>x"4800", 151=>x"5000", 152=>x"5400",
---- 153=>x"4900", 154=>x"4b00", 155=>x"5100", 156=>x"5700",
---- 157=>x"4a00", 158=>x"4e00", 159=>x"5100", 160=>x"5600",
---- 161=>x"4d00", 162=>x"4700", 163=>x"5000", 164=>x"5400",
---- 165=>x"4d00", 166=>x"4a00", 167=>x"5000", 168=>x"5900",
---- 169=>x"4c00", 170=>x"4a00", 171=>x"5000", 172=>x"5b00",
---- 173=>x"5000", 174=>x"4f00", 175=>x"5300", 176=>x"5900",
---- 177=>x"4f00", 178=>x"4a00", 179=>x"5000", 180=>x"5800",
---- 181=>x"4b00", 182=>x"4900", 183=>x"5200", 184=>x"5a00",
---- 185=>x"4c00", 186=>x"4b00", 187=>x"5300", 188=>x"a500",
---- 189=>x"4d00", 190=>x"4e00", 191=>x"5200", 192=>x"5c00",
---- 193=>x"4900", 194=>x"4e00", 195=>x"5300", 196=>x"5a00",
---- 197=>x"4d00", 198=>x"4c00", 199=>x"4d00", 200=>x"5900",
---- 201=>x"4c00", 202=>x"4b00", 203=>x"4d00", 204=>x"5e00",
---- 205=>x"4e00", 206=>x"b700", 207=>x"4f00", 208=>x"5e00",
---- 209=>x"4e00", 210=>x"4900", 211=>x"5000", 212=>x"5900",
---- 213=>x"5000", 214=>x"4c00", 215=>x"4e00", 216=>x"5e00",
---- 217=>x"4f00", 218=>x"4b00", 219=>x"5100", 220=>x"a400",
---- 221=>x"4e00", 222=>x"4a00", 223=>x"5200", 224=>x"5900",
---- 225=>x"4c00", 226=>x"4a00", 227=>x"5100", 228=>x"5c00",
---- 229=>x"5000", 230=>x"4b00", 231=>x"5000", 232=>x"5c00",
---- 233=>x"4900", 234=>x"4700", 235=>x"4f00", 236=>x"5600",
---- 237=>x"4600", 238=>x"4700", 239=>x"4f00", 240=>x"5300",
---- 241=>x"4800", 242=>x"4600", 243=>x"4b00", 244=>x"5600",
---- 245=>x"4700", 246=>x"4500", 247=>x"4a00", 248=>x"5500",
---- 249=>x"4d00", 250=>x"4900", 251=>x"4c00", 252=>x"5300",
---- 253=>x"4a00", 254=>x"4b00", 255=>x"4d00", 256=>x"5700",
---- 257=>x"4900", 258=>x"4b00", 259=>x"4d00", 260=>x"5900",
---- 261=>x"5000", 262=>x"4c00", 263=>x"5000", 264=>x"5900",
---- 265=>x"4f00", 266=>x"4c00", 267=>x"5100", 268=>x"5800",
---- 269=>x"4d00", 270=>x"4e00", 271=>x"5300", 272=>x"5b00",
---- 273=>x"4b00", 274=>x"4d00", 275=>x"5000", 276=>x"a700",
---- 277=>x"4d00", 278=>x"4e00", 279=>x"5100", 280=>x"5900",
---- 281=>x"4c00", 282=>x"4c00", 283=>x"4f00", 284=>x"5800",
---- 285=>x"4e00", 286=>x"4d00", 287=>x"5000", 288=>x"5b00",
---- 289=>x"4d00", 290=>x"4e00", 291=>x"5200", 292=>x"5b00",
---- 293=>x"4d00", 294=>x"4b00", 295=>x"4d00", 296=>x"5900",
---- 297=>x"4e00", 298=>x"4c00", 299=>x"4f00", 300=>x"5900",
---- 301=>x"4b00", 302=>x"4900", 303=>x"5000", 304=>x"5a00",
---- 305=>x"4c00", 306=>x"4b00", 307=>x"5100", 308=>x"5a00",
---- 309=>x"4f00", 310=>x"4d00", 311=>x"5100", 312=>x"5900",
---- 313=>x"5100", 314=>x"4d00", 315=>x"5200", 316=>x"5900",
---- 317=>x"5000", 318=>x"4c00", 319=>x"5000", 320=>x"5b00",
---- 321=>x"4f00", 322=>x"4f00", 323=>x"4f00", 324=>x"5b00",
---- 325=>x"4b00", 326=>x"4d00", 327=>x"5000", 328=>x"5e00",
---- 329=>x"5000", 330=>x"4d00", 331=>x"5300", 332=>x"5d00",
---- 333=>x"4f00", 334=>x"4c00", 335=>x"5300", 336=>x"6200",
---- 337=>x"4c00", 338=>x"4b00", 339=>x"5000", 340=>x"5a00",
---- 341=>x"4d00", 342=>x"4b00", 343=>x"4d00", 344=>x"5a00",
---- 345=>x"4f00", 346=>x"4700", 347=>x"5000", 348=>x"5a00",
---- 349=>x"4f00", 350=>x"4600", 351=>x"4c00", 352=>x"5900",
---- 353=>x"4900", 354=>x"4700", 355=>x"4e00", 356=>x"5b00",
---- 357=>x"4a00", 358=>x"4800", 359=>x"4d00", 360=>x"5b00",
---- 361=>x"4e00", 362=>x"4700", 363=>x"4c00", 364=>x"5800",
---- 365=>x"4b00", 366=>x"4700", 367=>x"4f00", 368=>x"5700",
---- 369=>x"4d00", 370=>x"4800", 371=>x"5100", 372=>x"5a00",
---- 373=>x"4b00", 374=>x"4900", 375=>x"5100", 376=>x"5900",
---- 377=>x"4e00", 378=>x"4d00", 379=>x"4e00", 380=>x"5c00",
---- 381=>x"4f00", 382=>x"4700", 383=>x"4d00", 384=>x"5d00",
---- 385=>x"4d00", 386=>x"4900", 387=>x"4e00", 388=>x"5c00",
---- 389=>x"4d00", 390=>x"4900", 391=>x"4c00", 392=>x"5c00",
---- 393=>x"4e00", 394=>x"4700", 395=>x"5000", 396=>x"a100",
---- 397=>x"4e00", 398=>x"4800", 399=>x"4e00", 400=>x"5c00",
---- 401=>x"4a00", 402=>x"4500", 403=>x"4b00", 404=>x"5b00",
---- 405=>x"4b00", 406=>x"4400", 407=>x"4c00", 408=>x"5900",
---- 409=>x"4d00", 410=>x"4900", 411=>x"4d00", 412=>x"5a00",
---- 413=>x"4900", 414=>x"4800", 415=>x"4d00", 416=>x"5b00",
---- 417=>x"4c00", 418=>x"4600", 419=>x"4b00", 420=>x"5900",
---- 421=>x"4b00", 422=>x"4400", 423=>x"4900", 424=>x"6000",
---- 425=>x"4a00", 426=>x"4300", 427=>x"4a00", 428=>x"5d00",
---- 429=>x"4900", 430=>x"4300", 431=>x"4e00", 432=>x"5c00",
---- 433=>x"4a00", 434=>x"4600", 435=>x"4b00", 436=>x"5e00",
---- 437=>x"4c00", 438=>x"4900", 439=>x"4900", 440=>x"5f00",
---- 441=>x"4d00", 442=>x"4800", 443=>x"4c00", 444=>x"6000",
---- 445=>x"4c00", 446=>x"4500", 447=>x"4d00", 448=>x"6200",
---- 449=>x"4d00", 450=>x"4600", 451=>x"4d00", 452=>x"6300",
---- 453=>x"5100", 454=>x"4900", 455=>x"4d00", 456=>x"6300",
---- 457=>x"5000", 458=>x"4700", 459=>x"4c00", 460=>x"6400",
---- 461=>x"5300", 462=>x"4a00", 463=>x"5300", 464=>x"6200",
---- 465=>x"5200", 466=>x"4f00", 467=>x"5400", 468=>x"6200",
---- 469=>x"4e00", 470=>x"4c00", 471=>x"4e00", 472=>x"5f00",
---- 473=>x"4d00", 474=>x"4b00", 475=>x"4e00", 476=>x"5e00",
---- 477=>x"5100", 478=>x"4d00", 479=>x"4f00", 480=>x"6200",
---- 481=>x"5100", 482=>x"4a00", 483=>x"4e00", 484=>x"6100",
---- 485=>x"5000", 486=>x"4a00", 487=>x"4d00", 488=>x"5f00",
---- 489=>x"5100", 490=>x"4900", 491=>x"5100", 492=>x"6100",
---- 493=>x"5200", 494=>x"4a00", 495=>x"5000", 496=>x"5e00",
---- 497=>x"4f00", 498=>x"4a00", 499=>x"4f00", 500=>x"5f00",
---- 501=>x"4e00", 502=>x"4c00", 503=>x"5000", 504=>x"5e00",
---- 505=>x"4e00", 506=>x"5100", 507=>x"5300", 508=>x"6400",
---- 509=>x"5000", 510=>x"4a00", 511=>x"5100", 512=>x"6000",
---- 513=>x"4e00", 514=>x"4a00", 515=>x"4f00", 516=>x"6300",
---- 517=>x"5100", 518=>x"4c00", 519=>x"4b00", 520=>x"6100",
---- 521=>x"5400", 522=>x"4800", 523=>x"4b00", 524=>x"6200",
---- 525=>x"4a00", 526=>x"4700", 527=>x"4900", 528=>x"6200",
---- 529=>x"4d00", 530=>x"4900", 531=>x"4a00", 532=>x"6100",
---- 533=>x"4c00", 534=>x"4900", 535=>x"5000", 536=>x"6500",
---- 537=>x"4f00", 538=>x"4900", 539=>x"5000", 540=>x"6500",
---- 541=>x"5300", 542=>x"4e00", 543=>x"5300", 544=>x"6900",
---- 545=>x"5300", 546=>x"5000", 547=>x"5400", 548=>x"6600",
---- 549=>x"5600", 550=>x"5400", 551=>x"5600", 552=>x"6600",
---- 553=>x"5700", 554=>x"5200", 555=>x"5600", 556=>x"6a00",
---- 557=>x"aa00", 558=>x"5000", 559=>x"5700", 560=>x"6c00",
---- 561=>x"5500", 562=>x"4f00", 563=>x"5600", 564=>x"6900",
---- 565=>x"5200", 566=>x"4c00", 567=>x"ac00", 568=>x"6800",
---- 569=>x"5300", 570=>x"5000", 571=>x"5500", 572=>x"6700",
---- 573=>x"5600", 574=>x"4d00", 575=>x"5500", 576=>x"6900",
---- 577=>x"5700", 578=>x"4f00", 579=>x"5300", 580=>x"6700",
---- 581=>x"5600", 582=>x"4e00", 583=>x"5200", 584=>x"6900",
---- 585=>x"5200", 586=>x"4d00", 587=>x"5300", 588=>x"6600",
---- 589=>x"5100", 590=>x"4e00", 591=>x"5000", 592=>x"9800",
---- 593=>x"5600", 594=>x"4c00", 595=>x"5300", 596=>x"6800",
---- 597=>x"5500", 598=>x"4c00", 599=>x"5500", 600=>x"6900",
---- 601=>x"5300", 602=>x"4d00", 603=>x"5200", 604=>x"6800",
---- 605=>x"5100", 606=>x"4c00", 607=>x"5400", 608=>x"9700",
---- 609=>x"5200", 610=>x"4800", 611=>x"4e00", 612=>x"6900",
---- 613=>x"4f00", 614=>x"4a00", 615=>x"4900", 616=>x"6500",
---- 617=>x"4d00", 618=>x"4800", 619=>x"4800", 620=>x"6500",
---- 621=>x"4f00", 622=>x"4800", 623=>x"4a00", 624=>x"6400",
---- 625=>x"4f00", 626=>x"4a00", 627=>x"4a00", 628=>x"6700",
---- 629=>x"5100", 630=>x"4900", 631=>x"4d00", 632=>x"6b00",
---- 633=>x"4f00", 634=>x"4400", 635=>x"4800", 636=>x"6800",
---- 637=>x"4e00", 638=>x"4700", 639=>x"5800", 640=>x"6d00",
---- 641=>x"5a00", 642=>x"6600", 643=>x"7800", 644=>x"6f00",
---- 645=>x"6500", 646=>x"5700", 647=>x"5100", 648=>x"7200",
---- 649=>x"5700", 650=>x"4600", 651=>x"4b00", 652=>x"6d00",
---- 653=>x"5300", 654=>x"4900", 655=>x"5000", 656=>x"6d00",
---- 657=>x"5500", 658=>x"4800", 659=>x"4e00", 660=>x"6c00",
---- 661=>x"5500", 662=>x"4a00", 663=>x"4e00", 664=>x"6d00",
---- 665=>x"5500", 666=>x"4b00", 667=>x"5000", 668=>x"6f00",
---- 669=>x"5500", 670=>x"4a00", 671=>x"4e00", 672=>x"6e00",
---- 673=>x"5600", 674=>x"4a00", 675=>x"4d00", 676=>x"6d00",
---- 677=>x"5700", 678=>x"4700", 679=>x"4a00", 680=>x"6d00",
---- 681=>x"5500", 682=>x"4600", 683=>x"4b00", 684=>x"7000",
---- 685=>x"5300", 686=>x"4500", 687=>x"4c00", 688=>x"7200",
---- 689=>x"5300", 690=>x"4500", 691=>x"4b00", 692=>x"6d00",
---- 693=>x"5300", 694=>x"4800", 695=>x"4900", 696=>x"6c00",
---- 697=>x"5200", 698=>x"4500", 699=>x"4900", 700=>x"6d00",
---- 701=>x"5200", 702=>x"3f00", 703=>x"6b00", 704=>x"6e00",
---- 705=>x"5000", 706=>x"5b00", 707=>x"9500", 708=>x"6800",
---- 709=>x"6600", 710=>x"9800", 711=>x"7f00", 712=>x"7800",
---- 713=>x"9800", 714=>x"8500", 715=>x"4e00", 716=>x"9000",
---- 717=>x"7c00", 718=>x"4c00", 719=>x"4400", 720=>x"7b00",
---- 721=>x"5300", 722=>x"3e00", 723=>x"4600", 724=>x"6900",
---- 725=>x"4d00", 726=>x"4400", 727=>x"4800", 728=>x"6900",
---- 729=>x"4f00", 730=>x"4300", 731=>x"4200", 732=>x"6a00",
---- 733=>x"b000", 734=>x"4100", 735=>x"4300", 736=>x"6e00",
---- 737=>x"4f00", 738=>x"4000", 739=>x"4200", 740=>x"6d00",
---- 741=>x"5100", 742=>x"4100", 743=>x"4300", 744=>x"6e00",
---- 745=>x"5800", 746=>x"4500", 747=>x"4400", 748=>x"6c00",
---- 749=>x"5500", 750=>x"4300", 751=>x"4400", 752=>x"6c00",
---- 753=>x"5200", 754=>x"4100", 755=>x"4900", 756=>x"6f00",
---- 757=>x"5200", 758=>x"4300", 759=>x"4800", 760=>x"6c00",
---- 761=>x"4f00", 762=>x"4200", 763=>x"4600", 764=>x"6c00",
---- 765=>x"4d00", 766=>x"3e00", 767=>x"4200", 768=>x"6a00",
---- 769=>x"4d00", 770=>x"3900", 771=>x"3b00", 772=>x"6600",
---- 773=>x"4500", 774=>x"3800", 775=>x"6900", 776=>x"5f00",
---- 777=>x"4800", 778=>x"7900", 779=>x"cf00", 780=>x"6100",
---- 781=>x"8800", 782=>x"d700", 783=>x"9900", 784=>x"9c00",
---- 785=>x"d400", 786=>x"9100", 787=>x"3e00", 788=>x"c400",
---- 789=>x"7a00", 790=>x"3700", 791=>x"5100", 792=>x"7a00",
---- 793=>x"4000", 794=>x"4100", 795=>x"4f00", 796=>x"6300",
---- 797=>x"4c00", 798=>x"4100", 799=>x"5700", 800=>x"6c00",
---- 801=>x"4c00", 802=>x"5400", 803=>x"7100", 804=>x"6700",
---- 805=>x"5600", 806=>x"7500", 807=>x"8200", 808=>x"7200",
---- 809=>x"7c00", 810=>x"8600", 811=>x"7d00", 812=>x"8900",
---- 813=>x"ae00", 814=>x"8000", 815=>x"7300", 816=>x"4400",
---- 817=>x"c200", 818=>x"5e00", 819=>x"6100", 820=>x"de00",
---- 821=>x"a700", 822=>x"5b00", 823=>x"5700", 824=>x"de00",
---- 825=>x"9000", 826=>x"8200", 827=>x"9200", 828=>x"cd00",
---- 829=>x"7700", 830=>x"5b00", 831=>x"9e00", 832=>x"a800",
---- 833=>x"7600", 834=>x"4f00", 835=>x"4c00", 836=>x"b300",
---- 837=>x"7800", 838=>x"5a00", 839=>x"3a00", 840=>x"c000",
---- 841=>x"7700", 842=>x"5600", 843=>x"5a00", 844=>x"8100",
---- 845=>x"9200", 846=>x"6d00", 847=>x"6500", 848=>x"6d00",
---- 849=>x"ab00", 850=>x"a200", 851=>x"3700", 852=>x"6d00",
---- 853=>x"7100", 854=>x"7700", 855=>x"4100", 856=>x"7800",
---- 857=>x"8e00", 858=>x"9200", 859=>x"3d00", 860=>x"9800",
---- 861=>x"9100", 862=>x"6700", 863=>x"2b00", 864=>x"9e00",
---- 865=>x"8c00", 866=>x"5c00", 867=>x"2c00", 868=>x"9500",
---- 869=>x"7d00", 870=>x"3300", 871=>x"2a00", 872=>x"8d00",
---- 873=>x"7600", 874=>x"2a00", 875=>x"2d00", 876=>x"8400",
---- 877=>x"7000", 878=>x"3500", 879=>x"3800", 880=>x"7e00",
---- 881=>x"6900", 882=>x"4300", 883=>x"3e00", 884=>x"8000",
---- 885=>x"7f00", 886=>x"5100", 887=>x"3100", 888=>x"8a00",
---- 889=>x"8a00", 890=>x"4c00", 891=>x"3f00", 892=>x"9400",
---- 893=>x"6f00", 894=>x"4400", 895=>x"3d00", 896=>x"9100",
---- 897=>x"6900", 898=>x"3d00", 899=>x"2f00", 900=>x"9800",
---- 901=>x"6d00", 902=>x"4000", 903=>x"3500", 904=>x"9c00",
---- 905=>x"7e00", 906=>x"4600", 907=>x"3700", 908=>x"9f00",
---- 909=>x"8600", 910=>x"4000", 911=>x"4a00", 912=>x"a400",
---- 913=>x"8700", 914=>x"4300", 915=>x"5800", 916=>x"9b00",
---- 917=>x"9100", 918=>x"4500", 919=>x"5800", 920=>x"8d00",
---- 921=>x"8c00", 922=>x"4500", 923=>x"5100", 924=>x"8100",
---- 925=>x"7f00", 926=>x"5000", 927=>x"5600", 928=>x"7f00",
---- 929=>x"7300", 930=>x"5400", 931=>x"5200", 932=>x"8100",
---- 933=>x"7200", 934=>x"5800", 935=>x"5000", 936=>x"6e00",
---- 937=>x"7100", 938=>x"6300", 939=>x"5400", 940=>x"5100",
---- 941=>x"7000", 942=>x"6700", 943=>x"5500", 944=>x"5000",
---- 945=>x"7500", 946=>x"6100", 947=>x"4400", 948=>x"5700",
---- 949=>x"7d00", 950=>x"6c00", 951=>x"3900", 952=>x"5f00",
---- 953=>x"8100", 954=>x"7200", 955=>x"3f00", 956=>x"6700",
---- 957=>x"7d00", 958=>x"6a00", 959=>x"4c00", 960=>x"6700",
---- 961=>x"7a00", 962=>x"6300", 963=>x"4e00", 964=>x"6a00",
---- 965=>x"8500", 966=>x"6000", 967=>x"4400", 968=>x"6d00",
---- 969=>x"7a00", 970=>x"5b00", 971=>x"3800", 972=>x"6400",
---- 973=>x"7a00", 974=>x"6400", 975=>x"3200", 976=>x"5600",
---- 977=>x"7300", 978=>x"5c00", 979=>x"2d00", 980=>x"5400",
---- 981=>x"6400", 982=>x"5100", 983=>x"2900", 984=>x"4900",
---- 985=>x"5100", 986=>x"3d00", 987=>x"2b00", 988=>x"4500",
---- 989=>x"4900", 990=>x"3400", 991=>x"d500", 992=>x"4600",
---- 993=>x"4700", 994=>x"3900", 995=>x"3200", 996=>x"4100",
---- 997=>x"4100", 998=>x"4300", 999=>x"3d00", 1000=>x"3400",
---- 1001=>x"3b00", 1002=>x"3a00", 1003=>x"3600", 1004=>x"4700",
---- 1005=>x"3a00", 1006=>x"3300", 1007=>x"3200", 1008=>x"5c00",
---- 1009=>x"3a00", 1010=>x"2e00", 1011=>x"3100", 1012=>x"5500",
---- 1013=>x"3300", 1014=>x"3200", 1015=>x"2e00", 1016=>x"4700",
---- 1017=>x"3600", 1018=>x"3c00", 1019=>x"2b00", 1020=>x"4600",
---- 1021=>x"3900", 1022=>x"3800", 1023=>x"2800"),
----
---- 9 => (0=>x"6400", 1=>x"6700", 2=>x"6900", 3=>x"6900", 4=>x"6400",
---- 5=>x"6700", 6=>x"6900", 7=>x"6900", 8=>x"9c00",
---- 9=>x"6600", 10=>x"6900", 11=>x"6900", 12=>x"6100",
---- 13=>x"6000", 14=>x"6900", 15=>x"6c00", 16=>x"5f00",
---- 17=>x"6400", 18=>x"6600", 19=>x"6800", 20=>x"6200",
---- 21=>x"6100", 22=>x"6300", 23=>x"6700", 24=>x"5d00",
---- 25=>x"6000", 26=>x"6300", 27=>x"6900", 28=>x"5d00",
---- 29=>x"6500", 30=>x"6500", 31=>x"6600", 32=>x"5c00",
---- 33=>x"6500", 34=>x"9700", 35=>x"6200", 36=>x"5f00",
---- 37=>x"6400", 38=>x"6600", 39=>x"6200", 40=>x"5e00",
---- 41=>x"6100", 42=>x"6700", 43=>x"6700", 44=>x"6100",
---- 45=>x"6200", 46=>x"6400", 47=>x"6600", 48=>x"6000",
---- 49=>x"6000", 50=>x"6300", 51=>x"6800", 52=>x"5d00",
---- 53=>x"6000", 54=>x"6500", 55=>x"6700", 56=>x"5f00",
---- 57=>x"6200", 58=>x"6400", 59=>x"6700", 60=>x"6100",
---- 61=>x"6200", 62=>x"6200", 63=>x"6800", 64=>x"5f00",
---- 65=>x"6000", 66=>x"6400", 67=>x"6400", 68=>x"5f00",
---- 69=>x"6400", 70=>x"6200", 71=>x"6700", 72=>x"6100",
---- 73=>x"6100", 74=>x"6500", 75=>x"6600", 76=>x"5f00",
---- 77=>x"5f00", 78=>x"6400", 79=>x"6500", 80=>x"5e00",
---- 81=>x"6000", 82=>x"6800", 83=>x"6800", 84=>x"5c00",
---- 85=>x"6200", 86=>x"6700", 87=>x"6700", 88=>x"5e00",
---- 89=>x"6200", 90=>x"6400", 91=>x"6500", 92=>x"5d00",
---- 93=>x"5f00", 94=>x"6200", 95=>x"6600", 96=>x"5e00",
---- 97=>x"6000", 98=>x"6200", 99=>x"6500", 100=>x"5c00",
---- 101=>x"6000", 102=>x"6100", 103=>x"6300", 104=>x"5e00",
---- 105=>x"5c00", 106=>x"6200", 107=>x"6500", 108=>x"5d00",
---- 109=>x"5e00", 110=>x"6300", 111=>x"6200", 112=>x"5600",
---- 113=>x"5b00", 114=>x"6000", 115=>x"6000", 116=>x"5a00",
---- 117=>x"5f00", 118=>x"9c00", 119=>x"6000", 120=>x"5f00",
---- 121=>x"5b00", 122=>x"5e00", 123=>x"6100", 124=>x"5700",
---- 125=>x"5600", 126=>x"5a00", 127=>x"5c00", 128=>x"5300",
---- 129=>x"5600", 130=>x"5b00", 131=>x"5e00", 132=>x"5200",
---- 133=>x"5700", 134=>x"5b00", 135=>x"5d00", 136=>x"5200",
---- 137=>x"5a00", 138=>x"5e00", 139=>x"5d00", 140=>x"5700",
---- 141=>x"5800", 142=>x"5900", 143=>x"5d00", 144=>x"5600",
---- 145=>x"5800", 146=>x"5b00", 147=>x"5f00", 148=>x"5600",
---- 149=>x"5a00", 150=>x"5e00", 151=>x"6000", 152=>x"5400",
---- 153=>x"5800", 154=>x"5c00", 155=>x"6000", 156=>x"5800",
---- 157=>x"5600", 158=>x"5c00", 159=>x"6200", 160=>x"5500",
---- 161=>x"5900", 162=>x"5f00", 163=>x"6100", 164=>x"5800",
---- 165=>x"5a00", 166=>x"5e00", 167=>x"5f00", 168=>x"5600",
---- 169=>x"5a00", 170=>x"6100", 171=>x"5f00", 172=>x"5800",
---- 173=>x"5a00", 174=>x"5c00", 175=>x"5c00", 176=>x"5500",
---- 177=>x"5b00", 178=>x"5c00", 179=>x"5e00", 180=>x"5800",
---- 181=>x"5b00", 182=>x"5d00", 183=>x"6200", 184=>x"5800",
---- 185=>x"5a00", 186=>x"6000", 187=>x"6100", 188=>x"5800",
---- 189=>x"5f00", 190=>x"6200", 191=>x"6100", 192=>x"5900",
---- 193=>x"5b00", 194=>x"6200", 195=>x"5d00", 196=>x"5600",
---- 197=>x"5c00", 198=>x"6000", 199=>x"6100", 200=>x"5600",
---- 201=>x"5900", 202=>x"5e00", 203=>x"6100", 204=>x"5600",
---- 205=>x"5800", 206=>x"5e00", 207=>x"5f00", 208=>x"5500",
---- 209=>x"5a00", 210=>x"5e00", 211=>x"5e00", 212=>x"5500",
---- 213=>x"5b00", 214=>x"5e00", 215=>x"5f00", 216=>x"5500",
---- 217=>x"5a00", 218=>x"5c00", 219=>x"5b00", 220=>x"5500",
---- 221=>x"5400", 222=>x"5a00", 223=>x"5d00", 224=>x"5600",
---- 225=>x"5600", 226=>x"5c00", 227=>x"6000", 228=>x"5400",
---- 229=>x"5a00", 230=>x"5d00", 231=>x"5f00", 232=>x"5000",
---- 233=>x"5600", 234=>x"5800", 235=>x"5800", 236=>x"5300",
---- 237=>x"5500", 238=>x"5800", 239=>x"5800", 240=>x"4f00",
---- 241=>x"5300", 242=>x"5900", 243=>x"5c00", 244=>x"4d00",
---- 245=>x"5200", 246=>x"5b00", 247=>x"5f00", 248=>x"4900",
---- 249=>x"5300", 250=>x"5800", 251=>x"5f00", 252=>x"4f00",
---- 253=>x"5500", 254=>x"5b00", 255=>x"5e00", 256=>x"5000",
---- 257=>x"5700", 258=>x"5b00", 259=>x"5c00", 260=>x"5200",
---- 261=>x"5700", 262=>x"5b00", 263=>x"a100", 264=>x"5400",
---- 265=>x"5c00", 266=>x"6000", 267=>x"5f00", 268=>x"5500",
---- 269=>x"5700", 270=>x"5d00", 271=>x"5f00", 272=>x"5600",
---- 273=>x"5400", 274=>x"5d00", 275=>x"5f00", 276=>x"5500",
---- 277=>x"5a00", 278=>x"5d00", 279=>x"5f00", 280=>x"5600",
---- 281=>x"5d00", 282=>x"5d00", 283=>x"5e00", 284=>x"5900",
---- 285=>x"5b00", 286=>x"5d00", 287=>x"6000", 288=>x"5c00",
---- 289=>x"6200", 290=>x"5a00", 291=>x"5d00", 292=>x"5400",
---- 293=>x"5800", 294=>x"a500", 295=>x"5d00", 296=>x"5400",
---- 297=>x"5a00", 298=>x"5d00", 299=>x"5e00", 300=>x"5400",
---- 301=>x"5900", 302=>x"5b00", 303=>x"6000", 304=>x"5500",
---- 305=>x"5b00", 306=>x"5e00", 307=>x"6000", 308=>x"5800",
---- 309=>x"a500", 310=>x"5f00", 311=>x"5e00", 312=>x"5a00",
---- 313=>x"5d00", 314=>x"6000", 315=>x"5f00", 316=>x"5500",
---- 317=>x"5e00", 318=>x"6000", 319=>x"5f00", 320=>x"5500",
---- 321=>x"5c00", 322=>x"5e00", 323=>x"6100", 324=>x"5500",
---- 325=>x"5c00", 326=>x"5e00", 327=>x"6100", 328=>x"5700",
---- 329=>x"5d00", 330=>x"5e00", 331=>x"6100", 332=>x"5900",
---- 333=>x"5b00", 334=>x"5c00", 335=>x"6200", 336=>x"5600",
---- 337=>x"5900", 338=>x"5c00", 339=>x"5f00", 340=>x"5300",
---- 341=>x"5a00", 342=>x"5f00", 343=>x"6000", 344=>x"5400",
---- 345=>x"5800", 346=>x"a300", 347=>x"6200", 348=>x"5600",
---- 349=>x"5900", 350=>x"5b00", 351=>x"6100", 352=>x"5300",
---- 353=>x"5600", 354=>x"5c00", 355=>x"5f00", 356=>x"5100",
---- 357=>x"5600", 358=>x"5e00", 359=>x"5e00", 360=>x"5300",
---- 361=>x"5500", 362=>x"6000", 363=>x"5e00", 364=>x"5300",
---- 365=>x"5600", 366=>x"5e00", 367=>x"5f00", 368=>x"5300",
---- 369=>x"5900", 370=>x"5d00", 371=>x"6100", 372=>x"5100",
---- 373=>x"5a00", 374=>x"5e00", 375=>x"6000", 376=>x"5100",
---- 377=>x"5800", 378=>x"5e00", 379=>x"5d00", 380=>x"5400",
---- 381=>x"5b00", 382=>x"5c00", 383=>x"6000", 384=>x"5300",
---- 385=>x"5500", 386=>x"5c00", 387=>x"5e00", 388=>x"5200",
---- 389=>x"ac00", 390=>x"5b00", 391=>x"5e00", 392=>x"aa00",
---- 393=>x"5800", 394=>x"5d00", 395=>x"5e00", 396=>x"a900",
---- 397=>x"a600", 398=>x"5d00", 399=>x"5e00", 400=>x"5300",
---- 401=>x"5900", 402=>x"5b00", 403=>x"5b00", 404=>x"5300",
---- 405=>x"5700", 406=>x"5b00", 407=>x"5b00", 408=>x"5400",
---- 409=>x"5400", 410=>x"5a00", 411=>x"5d00", 412=>x"5200",
---- 413=>x"5300", 414=>x"5800", 415=>x"5d00", 416=>x"5000",
---- 417=>x"5500", 418=>x"5700", 419=>x"5b00", 420=>x"5000",
---- 421=>x"5400", 422=>x"5900", 423=>x"5a00", 424=>x"5100",
---- 425=>x"5200", 426=>x"5800", 427=>x"5900", 428=>x"4f00",
---- 429=>x"5200", 430=>x"5a00", 431=>x"5c00", 432=>x"5100",
---- 433=>x"5400", 434=>x"5c00", 435=>x"5a00", 436=>x"5200",
---- 437=>x"5800", 438=>x"5e00", 439=>x"5c00", 440=>x"5000",
---- 441=>x"5400", 442=>x"5d00", 443=>x"5f00", 444=>x"5100",
---- 445=>x"5400", 446=>x"5e00", 447=>x"5c00", 448=>x"4f00",
---- 449=>x"5400", 450=>x"5b00", 451=>x"5e00", 452=>x"4f00",
---- 453=>x"5300", 454=>x"5b00", 455=>x"5b00", 456=>x"5100",
---- 457=>x"5700", 458=>x"5d00", 459=>x"5e00", 460=>x"5300",
---- 461=>x"5700", 462=>x"5e00", 463=>x"6100", 464=>x"5800",
---- 465=>x"5a00", 466=>x"5f00", 467=>x"5e00", 468=>x"5900",
---- 469=>x"5c00", 470=>x"5e00", 471=>x"6000", 472=>x"5800",
---- 473=>x"5b00", 474=>x"5f00", 475=>x"5f00", 476=>x"5500",
---- 477=>x"5700", 478=>x"5e00", 479=>x"5f00", 480=>x"5500",
---- 481=>x"5600", 482=>x"5c00", 483=>x"6000", 484=>x"5200",
---- 485=>x"5900", 486=>x"5d00", 487=>x"6000", 488=>x"5400",
---- 489=>x"5700", 490=>x"5c00", 491=>x"5e00", 492=>x"5600",
---- 493=>x"5600", 494=>x"5b00", 495=>x"5d00", 496=>x"5500",
---- 497=>x"5300", 498=>x"5e00", 499=>x"6000", 500=>x"5500",
---- 501=>x"5800", 502=>x"5b00", 503=>x"6000", 504=>x"5500",
---- 505=>x"5900", 506=>x"5e00", 507=>x"6100", 508=>x"5700",
---- 509=>x"5900", 510=>x"5e00", 511=>x"6000", 512=>x"5300",
---- 513=>x"5300", 514=>x"5c00", 515=>x"6100", 516=>x"5200",
---- 517=>x"5500", 518=>x"5a00", 519=>x"5e00", 520=>x"5300",
---- 521=>x"5500", 522=>x"5900", 523=>x"5900", 524=>x"5100",
---- 525=>x"5600", 526=>x"5900", 527=>x"a500", 528=>x"5300",
---- 529=>x"5800", 530=>x"5d00", 531=>x"5f00", 532=>x"5600",
---- 533=>x"5a00", 534=>x"6000", 535=>x"6100", 536=>x"5500",
---- 537=>x"5b00", 538=>x"6200", 539=>x"6200", 540=>x"5600",
---- 541=>x"5c00", 542=>x"6200", 543=>x"6100", 544=>x"5a00",
---- 545=>x"5e00", 546=>x"6700", 547=>x"6600", 548=>x"5a00",
---- 549=>x"5e00", 550=>x"6300", 551=>x"6600", 552=>x"5d00",
---- 553=>x"6000", 554=>x"6600", 555=>x"6900", 556=>x"5c00",
---- 557=>x"6300", 558=>x"6600", 559=>x"6900", 560=>x"5b00",
---- 561=>x"6100", 562=>x"6500", 563=>x"9600", 564=>x"5c00",
---- 565=>x"5e00", 566=>x"6300", 567=>x"6700", 568=>x"5c00",
---- 569=>x"5d00", 570=>x"6300", 571=>x"6900", 572=>x"5900",
---- 573=>x"5f00", 574=>x"6400", 575=>x"6800", 576=>x"5a00",
---- 577=>x"5e00", 578=>x"6300", 579=>x"6800", 580=>x"5b00",
---- 581=>x"5c00", 582=>x"6200", 583=>x"6300", 584=>x"5900",
---- 585=>x"5a00", 586=>x"6100", 587=>x"6300", 588=>x"5400",
---- 589=>x"5a00", 590=>x"6300", 591=>x"7500", 592=>x"5a00",
---- 593=>x"5d00", 594=>x"6600", 595=>x"7200", 596=>x"5900",
---- 597=>x"5f00", 598=>x"6400", 599=>x"6800", 600=>x"5600",
---- 601=>x"5b00", 602=>x"6200", 603=>x"6800", 604=>x"5b00",
---- 605=>x"6100", 606=>x"6000", 607=>x"6300", 608=>x"5d00",
---- 609=>x"7e00", 610=>x"6b00", 611=>x"6100", 612=>x"6100",
---- 613=>x"8800", 614=>x"6200", 615=>x"5c00", 616=>x"5800",
---- 617=>x"8b00", 618=>x"7300", 619=>x"6000", 620=>x"b200",
---- 621=>x"7200", 622=>x"9500", 623=>x"8600", 624=>x"4f00",
---- 625=>x"5b00", 626=>x"6e00", 627=>x"7800", 628=>x"5200",
---- 629=>x"5800", 630=>x"5c00", 631=>x"6f00", 632=>x"5500",
---- 633=>x"6b00", 634=>x"8000", 635=>x"7d00", 636=>x"7800",
---- 637=>x"8c00", 638=>x"7d00", 639=>x"6700", 640=>x"7800",
---- 641=>x"6a00", 642=>x"5f00", 643=>x"6300", 644=>x"5200",
---- 645=>x"5700", 646=>x"5f00", 647=>x"6500", 648=>x"5500",
---- 649=>x"5b00", 650=>x"5e00", 651=>x"6500", 652=>x"5600",
---- 653=>x"5b00", 654=>x"6100", 655=>x"6400", 656=>x"5600",
---- 657=>x"5c00", 658=>x"6100", 659=>x"6400", 660=>x"5500",
---- 661=>x"5a00", 662=>x"5f00", 663=>x"6000", 664=>x"5600",
---- 665=>x"5a00", 666=>x"5d00", 667=>x"6200", 668=>x"5600",
---- 669=>x"5d00", 670=>x"5e00", 671=>x"6300", 672=>x"5200",
---- 673=>x"5900", 674=>x"5f00", 675=>x"5e00", 676=>x"af00",
---- 677=>x"5800", 678=>x"5d00", 679=>x"9b00", 680=>x"ac00",
---- 681=>x"5500", 682=>x"5800", 683=>x"7c00", 684=>x"5300",
---- 685=>x"5400", 686=>x"7200", 687=>x"9100", 688=>x"4e00",
---- 689=>x"6400", 690=>x"9000", 691=>x"7100", 692=>x"5100",
---- 693=>x"8500", 694=>x"7e00", 695=>x"5900", 696=>x"7000",
---- 697=>x"8800", 698=>x"5e00", 699=>x"5a00", 700=>x"9300",
---- 701=>x"6900", 702=>x"5500", 703=>x"5900", 704=>x"7600",
---- 705=>x"5200", 706=>x"5300", 707=>x"5e00", 708=>x"4d00",
---- 709=>x"5000", 710=>x"5700", 711=>x"7300", 712=>x"4c00",
---- 713=>x"5100", 714=>x"5d00", 715=>x"8900", 716=>x"4c00",
---- 717=>x"5100", 718=>x"6d00", 719=>x"9600", 720=>x"4b00",
---- 721=>x"5c00", 722=>x"9100", 723=>x"8900", 724=>x"5000",
---- 725=>x"8100", 726=>x"9900", 727=>x"6900", 728=>x"5d00",
---- 729=>x"9900", 730=>x"7700", 731=>x"5f00", 732=>x"6600",
---- 733=>x"9800", 734=>x"6400", 735=>x"6200", 736=>x"6800",
---- 737=>x"9400", 738=>x"6200", 739=>x"6000", 740=>x"5e00",
---- 741=>x"8900", 742=>x"6d00", 743=>x"6100", 744=>x"5300",
---- 745=>x"7600", 746=>x"7600", 747=>x"6b00", 748=>x"5300",
---- 749=>x"6700", 750=>x"6c00", 751=>x"6600", 752=>x"5400",
---- 753=>x"6500", 754=>x"6600", 755=>x"6600", 756=>x"5300",
---- 757=>x"6200", 758=>x"6600", 759=>x"5c00", 760=>x"5200",
---- 761=>x"5f00", 762=>x"7600", 763=>x"4800", 764=>x"4700",
---- 765=>x"6a00", 766=>x"6200", 767=>x"3500", 768=>x"6100",
---- 769=>x"8200", 770=>x"5200", 771=>x"5600", 772=>x"b800",
---- 773=>x"8b00", 774=>x"5f00", 775=>x"9000", 776=>x"9a00",
---- 777=>x"4500", 778=>x"6000", 779=>x"9100", 780=>x"5300",
---- 781=>x"4000", 782=>x"6300", 783=>x"8400", 784=>x"5600",
---- 785=>x"3c00", 786=>x"5800", 787=>x"5c00", 788=>x"4100",
---- 789=>x"3400", 790=>x"8700", 791=>x"4700", 792=>x"3900",
---- 793=>x"7100", 794=>x"9700", 795=>x"3000", 796=>x"6600",
---- 797=>x"9700", 798=>x"5a00", 799=>x"2400", 800=>x"a800",
---- 801=>x"7100", 802=>x"2a00", 803=>x"2800", 804=>x"bd00",
---- 805=>x"3f00", 806=>x"2900", 807=>x"2a00", 808=>x"9200",
---- 809=>x"2900", 810=>x"2b00", 811=>x"2a00", 812=>x"5d00",
---- 813=>x"2700", 814=>x"2c00", 815=>x"2d00", 816=>x"5700",
---- 817=>x"3800", 818=>x"2e00", 819=>x"2800", 820=>x"4200",
---- 821=>x"3c00", 822=>x"3800", 823=>x"2e00", 824=>x"3000",
---- 825=>x"2500", 826=>x"2d00", 827=>x"2f00", 828=>x"2b00",
---- 829=>x"2300", 830=>x"2900", 831=>x"2d00", 832=>x"2500",
---- 833=>x"2700", 834=>x"2f00", 835=>x"2c00", 836=>x"2a00",
---- 837=>x"2900", 838=>x"2b00", 839=>x"2c00", 840=>x"2700",
---- 841=>x"2700", 842=>x"2c00", 843=>x"2900", 844=>x"1f00",
---- 845=>x"2600", 846=>x"3100", 847=>x"2a00", 848=>x"2700",
---- 849=>x"2d00", 850=>x"2f00", 851=>x"2900", 852=>x"2200",
---- 853=>x"3100", 854=>x"2e00", 855=>x"2900", 856=>x"2d00",
---- 857=>x"3300", 858=>x"2f00", 859=>x"2c00", 860=>x"3500",
---- 861=>x"3100", 862=>x"2600", 863=>x"3200", 864=>x"3500",
---- 865=>x"2d00", 866=>x"2b00", 867=>x"4000", 868=>x"3400",
---- 869=>x"2f00", 870=>x"3800", 871=>x"3b00", 872=>x"3800",
---- 873=>x"3c00", 874=>x"3d00", 875=>x"2a00", 876=>x"4300",
---- 877=>x"3500", 878=>x"3000", 879=>x"2800", 880=>x"4000",
---- 881=>x"2d00", 882=>x"2b00", 883=>x"2b00", 884=>x"3500",
---- 885=>x"2d00", 886=>x"2d00", 887=>x"2e00", 888=>x"2c00",
---- 889=>x"2b00", 890=>x"2e00", 891=>x"2e00", 892=>x"2d00",
---- 893=>x"3100", 894=>x"2b00", 895=>x"3400", 896=>x"2e00",
---- 897=>x"3900", 898=>x"3100", 899=>x"2e00", 900=>x"2e00",
---- 901=>x"3800", 902=>x"3000", 903=>x"2b00", 904=>x"3200",
---- 905=>x"3200", 906=>x"2f00", 907=>x"2b00", 908=>x"3b00",
---- 909=>x"3100", 910=>x"2a00", 911=>x"2900", 912=>x"4000",
---- 913=>x"2e00", 914=>x"2600", 915=>x"2900", 916=>x"4000",
---- 917=>x"3000", 918=>x"2c00", 919=>x"2e00", 920=>x"3d00",
---- 921=>x"3600", 922=>x"2b00", 923=>x"2a00", 924=>x"4400",
---- 925=>x"3200", 926=>x"d800", 927=>x"2d00", 928=>x"5200",
---- 929=>x"2b00", 930=>x"2600", 931=>x"2d00", 932=>x"5a00",
---- 933=>x"2d00", 934=>x"2800", 935=>x"3000", 936=>x"5700",
---- 937=>x"2800", 938=>x"2600", 939=>x"3500", 940=>x"5400",
---- 941=>x"2600", 942=>x"2e00", 943=>x"3800", 944=>x"4200",
---- 945=>x"2800", 946=>x"3300", 947=>x"3100", 948=>x"3800",
---- 949=>x"2c00", 950=>x"3200", 951=>x"2e00", 952=>x"3200",
---- 953=>x"2b00", 954=>x"3500", 955=>x"3100", 956=>x"2700",
---- 957=>x"2a00", 958=>x"2f00", 959=>x"3500", 960=>x"3000",
---- 961=>x"2c00", 962=>x"3100", 963=>x"2e00", 964=>x"2b00",
---- 965=>x"3300", 966=>x"2f00", 967=>x"2d00", 968=>x"2700",
---- 969=>x"3500", 970=>x"2f00", 971=>x"3300", 972=>x"2a00",
---- 973=>x"3100", 974=>x"2a00", 975=>x"3600", 976=>x"2600",
---- 977=>x"2e00", 978=>x"2c00", 979=>x"3500", 980=>x"2c00",
---- 981=>x"2c00", 982=>x"3200", 983=>x"3500", 984=>x"3100",
---- 985=>x"2900", 986=>x"2a00", 987=>x"3000", 988=>x"3000",
---- 989=>x"2b00", 990=>x"3600", 991=>x"3200", 992=>x"3000",
---- 993=>x"2f00", 994=>x"3b00", 995=>x"3600", 996=>x"3000",
---- 997=>x"2e00", 998=>x"2f00", 999=>x"3000", 1000=>x"2d00",
---- 1001=>x"3300", 1002=>x"3600", 1003=>x"2d00", 1004=>x"3a00",
---- 1005=>x"2e00", 1006=>x"3300", 1007=>x"2d00", 1008=>x"3e00",
---- 1009=>x"2f00", 1010=>x"3800", 1011=>x"2f00", 1012=>x"3100",
---- 1013=>x"2b00", 1014=>x"3700", 1015=>x"3300", 1016=>x"2800",
---- 1017=>x"2e00", 1018=>x"3e00", 1019=>x"2e00", 1020=>x"2600",
---- 1021=>x"3300", 1022=>x"4400", 1023=>x"2700"),
----
---- 10 => (0=>x"6d00", 1=>x"6a00", 2=>x"6900", 3=>x"6d00", 4=>x"6e00",
---- 5=>x"6a00", 6=>x"6900", 7=>x"6e00", 8=>x"6d00",
---- 9=>x"6a00", 10=>x"6800", 11=>x"6c00", 12=>x"6700",
---- 13=>x"6800", 14=>x"6700", 15=>x"6800", 16=>x"9500",
---- 17=>x"6900", 18=>x"6500", 19=>x"6a00", 20=>x"9b00",
---- 21=>x"6600", 22=>x"6700", 23=>x"6700", 24=>x"6600",
---- 25=>x"6900", 26=>x"6a00", 27=>x"6b00", 28=>x"6900",
---- 29=>x"6e00", 30=>x"6b00", 31=>x"6b00", 32=>x"6a00",
---- 33=>x"6a00", 34=>x"6900", 35=>x"6a00", 36=>x"6600",
---- 37=>x"6700", 38=>x"6a00", 39=>x"6b00", 40=>x"6b00",
---- 41=>x"6c00", 42=>x"6b00", 43=>x"6c00", 44=>x"7000",
---- 45=>x"6700", 46=>x"6700", 47=>x"6700", 48=>x"6a00",
---- 49=>x"6800", 50=>x"6900", 51=>x"6600", 52=>x"6900",
---- 53=>x"6900", 54=>x"6900", 55=>x"6900", 56=>x"6700",
---- 57=>x"6800", 58=>x"6800", 59=>x"6b00", 60=>x"6b00",
---- 61=>x"6b00", 62=>x"6c00", 63=>x"6700", 64=>x"6900",
---- 65=>x"6b00", 66=>x"6c00", 67=>x"6c00", 68=>x"6800",
---- 69=>x"6900", 70=>x"6800", 71=>x"6a00", 72=>x"6800",
---- 73=>x"6700", 74=>x"6600", 75=>x"6500", 76=>x"6600",
---- 77=>x"6900", 78=>x"6500", 79=>x"6500", 80=>x"6700",
---- 81=>x"6700", 82=>x"6400", 83=>x"6700", 84=>x"6700",
---- 85=>x"9a00", 86=>x"6600", 87=>x"6700", 88=>x"6700",
---- 89=>x"6600", 90=>x"6900", 91=>x"6700", 92=>x"6800",
---- 93=>x"6900", 94=>x"6900", 95=>x"6b00", 96=>x"6700",
---- 97=>x"6900", 98=>x"6900", 99=>x"6c00", 100=>x"6700",
---- 101=>x"6700", 102=>x"6600", 103=>x"6700", 104=>x"6800",
---- 105=>x"6900", 106=>x"6700", 107=>x"6800", 108=>x"6500",
---- 109=>x"6900", 110=>x"6500", 111=>x"6500", 112=>x"6300",
---- 113=>x"6400", 114=>x"6800", 115=>x"6300", 116=>x"5f00",
---- 117=>x"6100", 118=>x"6300", 119=>x"6600", 120=>x"6500",
---- 121=>x"6500", 122=>x"6400", 123=>x"9d00", 124=>x"6100",
---- 125=>x"6400", 126=>x"6100", 127=>x"5f00", 128=>x"5f00",
---- 129=>x"5e00", 130=>x"5d00", 131=>x"6200", 132=>x"5e00",
---- 133=>x"5f00", 134=>x"5f00", 135=>x"6200", 136=>x"5f00",
---- 137=>x"6100", 138=>x"6200", 139=>x"6100", 140=>x"6400",
---- 141=>x"6700", 142=>x"6600", 143=>x"6900", 144=>x"6400",
---- 145=>x"6500", 146=>x"6000", 147=>x"6700", 148=>x"6100",
---- 149=>x"6200", 150=>x"6100", 151=>x"6600", 152=>x"6500",
---- 153=>x"6200", 154=>x"6200", 155=>x"6400", 156=>x"6900",
---- 157=>x"6200", 158=>x"6300", 159=>x"6400", 160=>x"6100",
---- 161=>x"6000", 162=>x"6000", 163=>x"6100", 164=>x"5f00",
---- 165=>x"6500", 166=>x"6900", 167=>x"6000", 168=>x"6100",
---- 169=>x"6300", 170=>x"6300", 171=>x"6300", 172=>x"6000",
---- 173=>x"6300", 174=>x"6300", 175=>x"6300", 176=>x"5f00",
---- 177=>x"5e00", 178=>x"6200", 179=>x"6600", 180=>x"5f00",
---- 181=>x"5e00", 182=>x"6500", 183=>x"6700", 184=>x"6100",
---- 185=>x"5f00", 186=>x"6200", 187=>x"6300", 188=>x"6700",
---- 189=>x"6200", 190=>x"6100", 191=>x"6100", 192=>x"6400",
---- 193=>x"6600", 194=>x"6100", 195=>x"6300", 196=>x"6300",
---- 197=>x"6300", 198=>x"6300", 199=>x"6500", 200=>x"6000",
---- 201=>x"6600", 202=>x"6300", 203=>x"6400", 204=>x"6200",
---- 205=>x"6200", 206=>x"6200", 207=>x"6100", 208=>x"6100",
---- 209=>x"6000", 210=>x"6000", 211=>x"6600", 212=>x"5f00",
---- 213=>x"6000", 214=>x"6100", 215=>x"6100", 216=>x"6000",
---- 217=>x"6200", 218=>x"6400", 219=>x"6200", 220=>x"5f00",
---- 221=>x"6300", 222=>x"6300", 223=>x"6200", 224=>x"5e00",
---- 225=>x"6100", 226=>x"5d00", 227=>x"6200", 228=>x"5c00",
---- 229=>x"5d00", 230=>x"6100", 231=>x"6300", 232=>x"5c00",
---- 233=>x"5f00", 234=>x"5f00", 235=>x"5f00", 236=>x"5e00",
---- 237=>x"5d00", 238=>x"5f00", 239=>x"6000", 240=>x"5d00",
---- 241=>x"6100", 242=>x"6200", 243=>x"6200", 244=>x"5b00",
---- 245=>x"5e00", 246=>x"6200", 247=>x"6200", 248=>x"5e00",
---- 249=>x"6200", 250=>x"6400", 251=>x"6300", 252=>x"6200",
---- 253=>x"6500", 254=>x"6400", 255=>x"6300", 256=>x"6100",
---- 257=>x"6100", 258=>x"6200", 259=>x"6300", 260=>x"6100",
---- 261=>x"6400", 262=>x"6300", 263=>x"6500", 264=>x"6300",
---- 265=>x"6500", 266=>x"6300", 267=>x"6700", 268=>x"6200",
---- 269=>x"6200", 270=>x"6300", 271=>x"6700", 272=>x"6500",
---- 273=>x"6600", 274=>x"6200", 275=>x"6400", 276=>x"6300",
---- 277=>x"6500", 278=>x"6400", 279=>x"6600", 280=>x"6200",
---- 281=>x"6200", 282=>x"6100", 283=>x"6600", 284=>x"6400",
---- 285=>x"6300", 286=>x"6100", 287=>x"6200", 288=>x"6100",
---- 289=>x"6400", 290=>x"6300", 291=>x"6400", 292=>x"5e00",
---- 293=>x"6300", 294=>x"6400", 295=>x"6500", 296=>x"5d00",
---- 297=>x"5f00", 298=>x"6200", 299=>x"6700", 300=>x"6000",
---- 301=>x"6300", 302=>x"6000", 303=>x"6200", 304=>x"5f00",
---- 305=>x"6300", 306=>x"6300", 307=>x"6300", 308=>x"5f00",
---- 309=>x"6400", 310=>x"6400", 311=>x"6400", 312=>x"5f00",
---- 313=>x"6300", 314=>x"6700", 315=>x"9a00", 316=>x"9d00",
---- 317=>x"6600", 318=>x"6300", 319=>x"6100", 320=>x"6200",
---- 321=>x"6600", 322=>x"6300", 323=>x"6200", 324=>x"6000",
---- 325=>x"6300", 326=>x"6300", 327=>x"6300", 328=>x"6200",
---- 329=>x"6200", 330=>x"6200", 331=>x"6200", 332=>x"6300",
---- 333=>x"6100", 334=>x"6300", 335=>x"6000", 336=>x"5f00",
---- 337=>x"6300", 338=>x"6000", 339=>x"5f00", 340=>x"5c00",
---- 341=>x"6100", 342=>x"6300", 343=>x"6100", 344=>x"6400",
---- 345=>x"6000", 346=>x"6200", 347=>x"6100", 348=>x"6300",
---- 349=>x"6000", 350=>x"6100", 351=>x"6100", 352=>x"6100",
---- 353=>x"6400", 354=>x"6000", 355=>x"6200", 356=>x"5d00",
---- 357=>x"5f00", 358=>x"6000", 359=>x"6400", 360=>x"6200",
---- 361=>x"6000", 362=>x"6200", 363=>x"6300", 364=>x"5e00",
---- 365=>x"6300", 366=>x"6300", 367=>x"6100", 368=>x"6000",
---- 369=>x"6000", 370=>x"6200", 371=>x"6200", 372=>x"5f00",
---- 373=>x"6000", 374=>x"6300", 375=>x"6200", 376=>x"5e00",
---- 377=>x"6100", 378=>x"6500", 379=>x"6200", 380=>x"6000",
---- 381=>x"5f00", 382=>x"6000", 383=>x"5f00", 384=>x"5e00",
---- 385=>x"5e00", 386=>x"5f00", 387=>x"6200", 388=>x"6000",
---- 389=>x"6000", 390=>x"5f00", 391=>x"6400", 392=>x"5f00",
---- 393=>x"6000", 394=>x"5f00", 395=>x"6100", 396=>x"5e00",
---- 397=>x"6000", 398=>x"5f00", 399=>x"6000", 400=>x"5d00",
---- 401=>x"6000", 402=>x"6000", 403=>x"5f00", 404=>x"5e00",
---- 405=>x"5e00", 406=>x"a100", 407=>x"6000", 408=>x"5e00",
---- 409=>x"5e00", 410=>x"6200", 411=>x"6300", 412=>x"5b00",
---- 413=>x"6100", 414=>x"6000", 415=>x"6100", 416=>x"5c00",
---- 417=>x"6200", 418=>x"6100", 419=>x"5f00", 420=>x"5e00",
---- 421=>x"5f00", 422=>x"5d00", 423=>x"5f00", 424=>x"5d00",
---- 425=>x"6000", 426=>x"6000", 427=>x"6100", 428=>x"5c00",
---- 429=>x"6200", 430=>x"6400", 431=>x"6400", 432=>x"5e00",
---- 433=>x"6000", 434=>x"6100", 435=>x"6200", 436=>x"6100",
---- 437=>x"6200", 438=>x"6200", 439=>x"6300", 440=>x"5d00",
---- 441=>x"6100", 442=>x"6300", 443=>x"6400", 444=>x"5f00",
---- 445=>x"6000", 446=>x"9d00", 447=>x"6300", 448=>x"5e00",
---- 449=>x"6300", 450=>x"6300", 451=>x"6300", 452=>x"5f00",
---- 453=>x"6200", 454=>x"6700", 455=>x"6500", 456=>x"6100",
---- 457=>x"6400", 458=>x"6600", 459=>x"6600", 460=>x"6600",
---- 461=>x"6600", 462=>x"6500", 463=>x"6600", 464=>x"6100",
---- 465=>x"6300", 466=>x"6400", 467=>x"6500", 468=>x"6100",
---- 469=>x"6300", 470=>x"6400", 471=>x"6500", 472=>x"6200",
---- 473=>x"6500", 474=>x"6500", 475=>x"6600", 476=>x"9d00",
---- 477=>x"6200", 478=>x"6600", 479=>x"6500", 480=>x"6400",
---- 481=>x"6400", 482=>x"6800", 483=>x"6400", 484=>x"6400",
---- 485=>x"6500", 486=>x"6400", 487=>x"6400", 488=>x"6300",
---- 489=>x"6400", 490=>x"6700", 491=>x"6800", 492=>x"6100",
---- 493=>x"6500", 494=>x"6700", 495=>x"6700", 496=>x"6000",
---- 497=>x"6400", 498=>x"6600", 499=>x"6700", 500=>x"5f00",
---- 501=>x"9c00", 502=>x"6a00", 503=>x"6700", 504=>x"6200",
---- 505=>x"6500", 506=>x"9600", 507=>x"6600", 508=>x"6400",
---- 509=>x"6a00", 510=>x"6700", 511=>x"6300", 512=>x"6200",
---- 513=>x"9c00", 514=>x"6500", 515=>x"6500", 516=>x"6200",
---- 517=>x"6600", 518=>x"6500", 519=>x"6800", 520=>x"6000",
---- 521=>x"6100", 522=>x"6800", 523=>x"6600", 524=>x"5e00",
---- 525=>x"5e00", 526=>x"6200", 527=>x"6400", 528=>x"6100",
---- 529=>x"6200", 530=>x"9f00", 531=>x"6100", 532=>x"6100",
---- 533=>x"6300", 534=>x"6400", 535=>x"6000", 536=>x"6500",
---- 537=>x"6500", 538=>x"6500", 539=>x"6600", 540=>x"6700",
---- 541=>x"6a00", 542=>x"6600", 543=>x"6600", 544=>x"6600",
---- 545=>x"9400", 546=>x"6b00", 547=>x"6800", 548=>x"6b00",
---- 549=>x"6e00", 550=>x"6a00", 551=>x"6d00", 552=>x"6d00",
---- 553=>x"6f00", 554=>x"6f00", 555=>x"6c00", 556=>x"6e00",
---- 557=>x"6f00", 558=>x"6f00", 559=>x"9300", 560=>x"6b00",
---- 561=>x"7000", 562=>x"7000", 563=>x"6c00", 564=>x"6b00",
---- 565=>x"6d00", 566=>x"6b00", 567=>x"6b00", 568=>x"6a00",
---- 569=>x"6e00", 570=>x"6c00", 571=>x"6c00", 572=>x"6c00",
---- 573=>x"6f00", 574=>x"6d00", 575=>x"6e00", 576=>x"6b00",
---- 577=>x"6f00", 578=>x"6d00", 579=>x"6e00", 580=>x"6800",
---- 581=>x"6900", 582=>x"6d00", 583=>x"7500", 584=>x"6800",
---- 585=>x"7900", 586=>x"9200", 587=>x"9800", 588=>x"8400",
---- 589=>x"8600", 590=>x"8400", 591=>x"7b00", 592=>x"7100",
---- 593=>x"6e00", 594=>x"6d00", 595=>x"7300", 596=>x"6800",
---- 597=>x"6d00", 598=>x"7000", 599=>x"7500", 600=>x"6b00",
---- 601=>x"6c00", 602=>x"7000", 603=>x"7200", 604=>x"6800",
---- 605=>x"9400", 606=>x"6e00", 607=>x"6f00", 608=>x"6700",
---- 609=>x"6700", 610=>x"6c00", 611=>x"7f00", 612=>x"6600",
---- 613=>x"7d00", 614=>x"9d00", 615=>x"9c00", 616=>x"9000",
---- 617=>x"a100", 618=>x"8500", 619=>x"7800", 620=>x"8900",
---- 621=>x"7000", 622=>x"6800", 623=>x"7c00", 624=>x"8c00",
---- 625=>x"7500", 626=>x"7700", 627=>x"7d00", 628=>x"7a00",
---- 629=>x"7000", 630=>x"8100", 631=>x"8600", 632=>x"6f00",
---- 633=>x"6800", 634=>x"6f00", 635=>x"7800", 636=>x"6800",
---- 637=>x"6d00", 638=>x"7400", 639=>x"7500", 640=>x"6800",
---- 641=>x"7100", 642=>x"7900", 643=>x"7600", 644=>x"6500",
---- 645=>x"6d00", 646=>x"7a00", 647=>x"7600", 648=>x"6800",
---- 649=>x"6d00", 650=>x"7100", 651=>x"6500", 652=>x"6900",
---- 653=>x"6d00", 654=>x"7500", 655=>x"6600", 656=>x"6900",
---- 657=>x"7700", 658=>x"7900", 659=>x"6600", 660=>x"6b00",
---- 661=>x"7600", 662=>x"7400", 663=>x"7000", 664=>x"6700",
---- 665=>x"6b00", 666=>x"7b00", 667=>x"9300", 668=>x"6800",
---- 669=>x"7600", 670=>x"9500", 671=>x"8e00", 672=>x"6b00",
---- 673=>x"9300", 674=>x"8b00", 675=>x"6d00", 676=>x"8b00",
---- 677=>x"8a00", 678=>x"6e00", 679=>x"7700", 680=>x"8e00",
---- 681=>x"6b00", 682=>x"7600", 683=>x"7800", 684=>x"6d00",
---- 685=>x"6600", 686=>x"7f00", 687=>x"7500", 688=>x"6200",
---- 689=>x"6800", 690=>x"7b00", 691=>x"6700", 692=>x"6000",
---- 693=>x"6600", 694=>x"8000", 695=>x"6900", 696=>x"6200",
---- 697=>x"7400", 698=>x"9000", 699=>x"6500", 700=>x"7100",
---- 701=>x"9300", 702=>x"9600", 703=>x"5d00", 704=>x"7600",
---- 705=>x"9700", 706=>x"8300", 707=>x"5700", 708=>x"9200",
---- 709=>x"7f00", 710=>x"7500", 711=>x"5700", 712=>x"8700",
---- 713=>x"6e00", 714=>x"7100", 715=>x"5d00", 716=>x"7400",
---- 717=>x"6700", 718=>x"6900", 719=>x"5200", 720=>x"6600",
---- 721=>x"6e00", 722=>x"6400", 723=>x"3c00", 724=>x"6300",
---- 725=>x"7600", 726=>x"6300", 727=>x"3a00", 728=>x"6a00",
---- 729=>x"7600", 730=>x"4d00", 731=>x"3500", 732=>x"7100",
---- 733=>x"5f00", 734=>x"3500", 735=>x"3200", 736=>x"6200",
---- 737=>x"4d00", 738=>x"4000", 739=>x"3300", 740=>x"5d00",
---- 741=>x"5700", 742=>x"4200", 743=>x"4700", 744=>x"5b00",
---- 745=>x"4b00", 746=>x"4300", 747=>x"5d00", 748=>x"5d00",
---- 749=>x"4600", 750=>x"4b00", 751=>x"5900", 752=>x"5600",
---- 753=>x"3c00", 754=>x"4b00", 755=>x"3900", 756=>x"4100",
---- 757=>x"3c00", 758=>x"4100", 759=>x"3200", 760=>x"3000",
---- 761=>x"3900", 762=>x"3300", 763=>x"3500", 764=>x"3000",
---- 765=>x"3100", 766=>x"3900", 767=>x"4500", 768=>x"3e00",
---- 769=>x"2800", 770=>x"3f00", 771=>x"5f00", 772=>x"4100",
---- 773=>x"2500", 774=>x"3500", 775=>x"5300", 776=>x"3700",
---- 777=>x"2600", 778=>x"2b00", 779=>x"4d00", 780=>x"3600",
---- 781=>x"3400", 782=>x"2800", 783=>x"4700", 784=>x"2900",
---- 785=>x"2b00", 786=>x"2600", 787=>x"4400", 788=>x"2400",
---- 789=>x"2a00", 790=>x"2400", 791=>x"3d00", 792=>x"2600",
---- 793=>x"2a00", 794=>x"2400", 795=>x"3000", 796=>x"2900",
---- 797=>x"2b00", 798=>x"2700", 799=>x"2900", 800=>x"2800",
---- 801=>x"2700", 802=>x"2600", 803=>x"2d00", 804=>x"2a00",
---- 805=>x"2b00", 806=>x"2b00", 807=>x"2c00", 808=>x"2a00",
---- 809=>x"2a00", 810=>x"2a00", 811=>x"2500", 812=>x"2a00",
---- 813=>x"2400", 814=>x"2600", 815=>x"de00", 816=>x"2a00",
---- 817=>x"2500", 818=>x"2b00", 819=>x"2600", 820=>x"2f00",
---- 821=>x"2f00", 822=>x"2b00", 823=>x"2b00", 824=>x"3900",
---- 825=>x"3c00", 826=>x"3900", 827=>x"3a00", 828=>x"3200",
---- 829=>x"ca00", 830=>x"3100", 831=>x"3500", 832=>x"2a00",
---- 833=>x"3100", 834=>x"2c00", 835=>x"2d00", 836=>x"2700",
---- 837=>x"3100", 838=>x"2a00", 839=>x"3f00", 840=>x"2b00",
---- 841=>x"3300", 842=>x"2a00", 843=>x"5700", 844=>x"2d00",
---- 845=>x"2e00", 846=>x"3b00", 847=>x"5300", 848=>x"3200",
---- 849=>x"3600", 850=>x"4400", 851=>x"3800", 852=>x"2f00",
---- 853=>x"3b00", 854=>x"3a00", 855=>x"3500", 856=>x"3500",
---- 857=>x"3b00", 858=>x"3200", 859=>x"3500", 860=>x"4000",
---- 861=>x"3400", 862=>x"2e00", 863=>x"3400", 864=>x"3b00",
---- 865=>x"cf00", 866=>x"2c00", 867=>x"3200", 868=>x"3000",
---- 869=>x"2c00", 870=>x"2a00", 871=>x"2d00", 872=>x"2d00",
---- 873=>x"2c00", 874=>x"2a00", 875=>x"2e00", 876=>x"2c00",
---- 877=>x"3000", 878=>x"2d00", 879=>x"2d00", 880=>x"3000",
---- 881=>x"2e00", 882=>x"2c00", 883=>x"2f00", 884=>x"2e00",
---- 885=>x"2c00", 886=>x"3200", 887=>x"3100", 888=>x"2b00",
---- 889=>x"2b00", 890=>x"3200", 891=>x"3600", 892=>x"2f00",
---- 893=>x"2e00", 894=>x"3300", 895=>x"3100", 896=>x"2e00",
---- 897=>x"2c00", 898=>x"3100", 899=>x"3100", 900=>x"2b00",
---- 901=>x"2a00", 902=>x"3400", 903=>x"2f00", 904=>x"2600",
---- 905=>x"2d00", 906=>x"3700", 907=>x"2800", 908=>x"2700",
---- 909=>x"2d00", 910=>x"3600", 911=>x"4900", 912=>x"2c00",
---- 913=>x"4600", 914=>x"5400", 915=>x"5000", 916=>x"3300",
---- 917=>x"4000", 918=>x"3b00", 919=>x"3100", 920=>x"2d00",
---- 921=>x"2f00", 922=>x"2e00", 923=>x"3300", 924=>x"3000",
---- 925=>x"3600", 926=>x"3600", 927=>x"3200", 928=>x"3a00",
---- 929=>x"3900", 930=>x"2e00", 931=>x"2d00", 932=>x"3d00",
---- 933=>x"2d00", 934=>x"2c00", 935=>x"2d00", 936=>x"2f00",
---- 937=>x"2a00", 938=>x"2e00", 939=>x"2b00", 940=>x"2900",
---- 941=>x"2e00", 942=>x"2c00", 943=>x"2700", 944=>x"2700",
---- 945=>x"2c00", 946=>x"2b00", 947=>x"2b00", 948=>x"2b00",
---- 949=>x"2f00", 950=>x"3600", 951=>x"3b00", 952=>x"3100",
---- 953=>x"4100", 954=>x"4700", 955=>x"3200", 956=>x"3b00",
---- 957=>x"3b00", 958=>x"3500", 959=>x"2e00", 960=>x"2e00",
---- 961=>x"2f00", 962=>x"3100", 963=>x"2e00", 964=>x"3000",
---- 965=>x"2f00", 966=>x"3100", 967=>x"2d00", 968=>x"2f00",
---- 969=>x"2f00", 970=>x"2d00", 971=>x"3200", 972=>x"3300",
---- 973=>x"3800", 974=>x"2f00", 975=>x"3800", 976=>x"3300",
---- 977=>x"3a00", 978=>x"3000", 979=>x"3b00", 980=>x"3500",
---- 981=>x"3600", 982=>x"2800", 983=>x"3f00", 984=>x"3300",
---- 985=>x"3500", 986=>x"3300", 987=>x"3e00", 988=>x"2e00",
---- 989=>x"3100", 990=>x"3400", 991=>x"4000", 992=>x"2a00",
---- 993=>x"2d00", 994=>x"3800", 995=>x"4300", 996=>x"2e00",
---- 997=>x"3300", 998=>x"3600", 999=>x"3f00", 1000=>x"2f00",
---- 1001=>x"3400", 1002=>x"3900", 1003=>x"3f00", 1004=>x"2e00",
---- 1005=>x"3400", 1006=>x"3800", 1007=>x"3c00", 1008=>x"3500",
---- 1009=>x"3e00", 1010=>x"3d00", 1011=>x"3700", 1012=>x"3800",
---- 1013=>x"3600", 1014=>x"3c00", 1015=>x"3900", 1016=>x"3900",
---- 1017=>x"3d00", 1018=>x"3c00", 1019=>x"3e00", 1020=>x"3800",
---- 1021=>x"3700", 1022=>x"3c00", 1023=>x"4700"),
----
---- 11 => (0=>x"6c00", 1=>x"6a00", 2=>x"6d00", 3=>x"6c00", 4=>x"6c00",
---- 5=>x"6b00", 6=>x"6d00", 7=>x"6b00", 8=>x"6b00",
---- 9=>x"6a00", 10=>x"6d00", 11=>x"6b00", 12=>x"6700",
---- 13=>x"6800", 14=>x"6900", 15=>x"6800", 16=>x"6900",
---- 17=>x"6800", 18=>x"6800", 19=>x"6700", 20=>x"6800",
---- 21=>x"6b00", 22=>x"6700", 23=>x"6600", 24=>x"6c00",
---- 25=>x"6900", 26=>x"6600", 27=>x"6700", 28=>x"6b00",
---- 29=>x"6b00", 30=>x"6600", 31=>x"6800", 32=>x"6700",
---- 33=>x"9700", 34=>x"6700", 35=>x"6a00", 36=>x"6900",
---- 37=>x"6a00", 38=>x"6900", 39=>x"6a00", 40=>x"6800",
---- 41=>x"6800", 42=>x"6600", 43=>x"6500", 44=>x"6700",
---- 45=>x"9500", 46=>x"6500", 47=>x"6600", 48=>x"6400",
---- 49=>x"6a00", 50=>x"6700", 51=>x"6800", 52=>x"6900",
---- 53=>x"6a00", 54=>x"6600", 55=>x"6600", 56=>x"6a00",
---- 57=>x"6900", 58=>x"6800", 59=>x"6700", 60=>x"6900",
---- 61=>x"6a00", 62=>x"6600", 63=>x"6700", 64=>x"6b00",
---- 65=>x"6a00", 66=>x"6400", 67=>x"6600", 68=>x"6900",
---- 69=>x"6700", 70=>x"6700", 71=>x"6700", 72=>x"6700",
---- 73=>x"6700", 74=>x"6700", 75=>x"6400", 76=>x"6600",
---- 77=>x"6800", 78=>x"6600", 79=>x"6600", 80=>x"6600",
---- 81=>x"6500", 82=>x"6500", 83=>x"6700", 84=>x"6600",
---- 85=>x"6a00", 86=>x"6400", 87=>x"9800", 88=>x"6700",
---- 89=>x"6800", 90=>x"6a00", 91=>x"6600", 92=>x"6700",
---- 93=>x"6600", 94=>x"6900", 95=>x"6700", 96=>x"6700",
---- 97=>x"6600", 98=>x"6800", 99=>x"6600", 100=>x"6600",
---- 101=>x"6400", 102=>x"6700", 103=>x"6900", 104=>x"6600",
---- 105=>x"6a00", 106=>x"6700", 107=>x"6600", 108=>x"6800",
---- 109=>x"6900", 110=>x"6600", 111=>x"6700", 112=>x"6600",
---- 113=>x"6600", 114=>x"6700", 115=>x"6500", 116=>x"6500",
---- 117=>x"6300", 118=>x"9b00", 119=>x"6200", 120=>x"6300",
---- 121=>x"6500", 122=>x"6100", 123=>x"6400", 124=>x"6300",
---- 125=>x"6200", 126=>x"6200", 127=>x"6500", 128=>x"6400",
---- 129=>x"6300", 130=>x"6300", 131=>x"6300", 132=>x"6100",
---- 133=>x"6300", 134=>x"6400", 135=>x"6500", 136=>x"6200",
---- 137=>x"6500", 138=>x"6300", 139=>x"6300", 140=>x"6300",
---- 141=>x"6500", 142=>x"6500", 143=>x"6300", 144=>x"6600",
---- 145=>x"6400", 146=>x"6100", 147=>x"9d00", 148=>x"6400",
---- 149=>x"6600", 150=>x"9c00", 151=>x"6300", 152=>x"6200",
---- 153=>x"6400", 154=>x"6300", 155=>x"6500", 156=>x"9b00",
---- 157=>x"6100", 158=>x"6500", 159=>x"6200", 160=>x"6600",
---- 161=>x"6400", 162=>x"6200", 163=>x"6400", 164=>x"6400",
---- 165=>x"6500", 166=>x"6300", 167=>x"6300", 168=>x"6300",
---- 169=>x"6000", 170=>x"6800", 171=>x"6700", 172=>x"6200",
---- 173=>x"6400", 174=>x"6a00", 175=>x"6700", 176=>x"6600",
---- 177=>x"6600", 178=>x"6900", 179=>x"6500", 180=>x"6500",
---- 181=>x"6500", 182=>x"6900", 183=>x"6600", 184=>x"6200",
---- 185=>x"6300", 186=>x"6500", 187=>x"9c00", 188=>x"6300",
---- 189=>x"6200", 190=>x"6600", 191=>x"9e00", 192=>x"6400",
---- 193=>x"6400", 194=>x"6300", 195=>x"6600", 196=>x"6200",
---- 197=>x"6100", 198=>x"6200", 199=>x"6200", 200=>x"6200",
---- 201=>x"6500", 202=>x"6100", 203=>x"6400", 204=>x"6200",
---- 205=>x"6600", 206=>x"6300", 207=>x"6400", 208=>x"6700",
---- 209=>x"6500", 210=>x"6300", 211=>x"6300", 212=>x"6900",
---- 213=>x"6600", 214=>x"6300", 215=>x"6200", 216=>x"6500",
---- 217=>x"6400", 218=>x"6600", 219=>x"6400", 220=>x"6500",
---- 221=>x"6400", 222=>x"6500", 223=>x"6600", 224=>x"6400",
---- 225=>x"6600", 226=>x"6a00", 227=>x"6500", 228=>x"6500",
---- 229=>x"6200", 230=>x"6600", 231=>x"6300", 232=>x"6100",
---- 233=>x"6000", 234=>x"5f00", 235=>x"6000", 236=>x"5f00",
---- 237=>x"6100", 238=>x"6000", 239=>x"5e00", 240=>x"6100",
---- 241=>x"6200", 242=>x"6200", 243=>x"5f00", 244=>x"6200",
---- 245=>x"6500", 246=>x"6300", 247=>x"6300", 248=>x"6100",
---- 249=>x"6500", 250=>x"6400", 251=>x"6300", 252=>x"6300",
---- 253=>x"6600", 254=>x"6600", 255=>x"6300", 256=>x"6300",
---- 257=>x"6600", 258=>x"6600", 259=>x"6300", 260=>x"6400",
---- 261=>x"6500", 262=>x"6500", 263=>x"6500", 264=>x"6600",
---- 265=>x"6400", 266=>x"6800", 267=>x"6a00", 268=>x"6600",
---- 269=>x"6700", 270=>x"6900", 271=>x"6a00", 272=>x"6500",
---- 273=>x"6600", 274=>x"6500", 275=>x"6600", 276=>x"6500",
---- 277=>x"6800", 278=>x"6100", 279=>x"6500", 280=>x"6600",
---- 281=>x"6500", 282=>x"6500", 283=>x"6600", 284=>x"6600",
---- 285=>x"6400", 286=>x"6500", 287=>x"6500", 288=>x"6300",
---- 289=>x"6400", 290=>x"6300", 291=>x"6400", 292=>x"6400",
---- 293=>x"6100", 294=>x"6300", 295=>x"6200", 296=>x"6500",
---- 297=>x"6300", 298=>x"6200", 299=>x"6100", 300=>x"6100",
---- 301=>x"6300", 302=>x"6200", 303=>x"6400", 304=>x"6100",
---- 305=>x"6300", 306=>x"6500", 307=>x"6100", 308=>x"6400",
---- 309=>x"9f00", 310=>x"6400", 311=>x"6300", 312=>x"6400",
---- 313=>x"6000", 314=>x"6200", 315=>x"6400", 316=>x"6300",
---- 317=>x"6200", 318=>x"6300", 319=>x"6300", 320=>x"6200",
---- 321=>x"6400", 322=>x"6200", 323=>x"6200", 324=>x"6300",
---- 325=>x"5f00", 326=>x"5f00", 327=>x"6200", 328=>x"6200",
---- 329=>x"6000", 330=>x"6200", 331=>x"6200", 332=>x"6300",
---- 333=>x"6200", 334=>x"6400", 335=>x"6200", 336=>x"6200",
---- 337=>x"6000", 338=>x"6000", 339=>x"6100", 340=>x"6000",
---- 341=>x"5d00", 342=>x"6100", 343=>x"6300", 344=>x"5e00",
---- 345=>x"5d00", 346=>x"6200", 347=>x"6000", 348=>x"6200",
---- 349=>x"6300", 350=>x"6100", 351=>x"6100", 352=>x"6500",
---- 353=>x"6200", 354=>x"6100", 355=>x"6500", 356=>x"6600",
---- 357=>x"6400", 358=>x"6000", 359=>x"6700", 360=>x"6600",
---- 361=>x"6100", 362=>x"6100", 363=>x"6600", 364=>x"6100",
---- 365=>x"6200", 366=>x"6300", 367=>x"6600", 368=>x"6100",
---- 369=>x"6200", 370=>x"6500", 371=>x"6400", 372=>x"6400",
---- 373=>x"6200", 374=>x"6300", 375=>x"6500", 376=>x"6200",
---- 377=>x"6200", 378=>x"6200", 379=>x"6500", 380=>x"6100",
---- 381=>x"6200", 382=>x"6400", 383=>x"6500", 384=>x"6200",
---- 385=>x"5f00", 386=>x"6300", 387=>x"6300", 388=>x"6200",
---- 389=>x"6300", 390=>x"6200", 391=>x"9d00", 392=>x"6500",
---- 393=>x"6400", 394=>x"6500", 395=>x"6500", 396=>x"6300",
---- 397=>x"6100", 398=>x"6300", 399=>x"6300", 400=>x"6000",
---- 401=>x"5f00", 402=>x"6400", 403=>x"6600", 404=>x"6000",
---- 405=>x"6100", 406=>x"5f00", 407=>x"6000", 408=>x"6100",
---- 409=>x"6300", 410=>x"6000", 411=>x"5f00", 412=>x"6200",
---- 413=>x"6200", 414=>x"6000", 415=>x"6300", 416=>x"6000",
---- 417=>x"5f00", 418=>x"6000", 419=>x"6300", 420=>x"6100",
---- 421=>x"6000", 422=>x"6100", 423=>x"6200", 424=>x"5f00",
---- 425=>x"6000", 426=>x"5f00", 427=>x"5d00", 428=>x"6200",
---- 429=>x"9c00", 430=>x"6400", 431=>x"6100", 432=>x"6300",
---- 433=>x"6300", 434=>x"6400", 435=>x"6200", 436=>x"6400",
---- 437=>x"9a00", 438=>x"6200", 439=>x"6400", 440=>x"6200",
---- 441=>x"6700", 442=>x"6400", 443=>x"6300", 444=>x"6400",
---- 445=>x"6400", 446=>x"6700", 447=>x"6500", 448=>x"6200",
---- 449=>x"6500", 450=>x"6500", 451=>x"6500", 452=>x"6700",
---- 453=>x"6900", 454=>x"6700", 455=>x"6700", 456=>x"6800",
---- 457=>x"6900", 458=>x"6800", 459=>x"6800", 460=>x"6900",
---- 461=>x"6900", 462=>x"6600", 463=>x"6400", 464=>x"6500",
---- 465=>x"6400", 466=>x"6500", 467=>x"6700", 468=>x"6500",
---- 469=>x"6600", 470=>x"6800", 471=>x"6900", 472=>x"6600",
---- 473=>x"6600", 474=>x"6900", 475=>x"6900", 476=>x"6800",
---- 477=>x"6700", 478=>x"6900", 479=>x"6a00", 480=>x"6500",
---- 481=>x"6800", 482=>x"6800", 483=>x"6800", 484=>x"9800",
---- 485=>x"6900", 486=>x"6700", 487=>x"6600", 488=>x"6600",
---- 489=>x"6600", 490=>x"6400", 491=>x"6500", 492=>x"6700",
---- 493=>x"6600", 494=>x"6400", 495=>x"6600", 496=>x"6600",
---- 497=>x"6600", 498=>x"9600", 499=>x"6800", 500=>x"6600",
---- 501=>x"6400", 502=>x"6400", 503=>x"6300", 504=>x"6600",
---- 505=>x"6500", 506=>x"6400", 507=>x"6300", 508=>x"6600",
---- 509=>x"6400", 510=>x"6700", 511=>x"6400", 512=>x"6600",
---- 513=>x"6300", 514=>x"6200", 515=>x"6400", 516=>x"6500",
---- 517=>x"6500", 518=>x"6400", 519=>x"6400", 520=>x"6300",
---- 521=>x"6300", 522=>x"6200", 523=>x"6200", 524=>x"6000",
---- 525=>x"5e00", 526=>x"6200", 527=>x"5e00", 528=>x"6100",
---- 529=>x"6300", 530=>x"6200", 531=>x"6000", 532=>x"6100",
---- 533=>x"6200", 534=>x"6400", 535=>x"6500", 536=>x"6700",
---- 537=>x"6600", 538=>x"6700", 539=>x"6200", 540=>x"6a00",
---- 541=>x"6600", 542=>x"6800", 543=>x"6a00", 544=>x"6900",
---- 545=>x"6600", 546=>x"6900", 547=>x"6300", 548=>x"9200",
---- 549=>x"7900", 550=>x"4b00", 551=>x"3100", 552=>x"7600",
---- 553=>x"8900", 554=>x"2900", 555=>x"2600", 556=>x"7600",
---- 557=>x"8900", 558=>x"3000", 559=>x"3000", 560=>x"6b00",
---- 561=>x"8a00", 562=>x"6d00", 563=>x"7000", 564=>x"6600",
---- 565=>x"8000", 566=>x"9f00", 567=>x"9200", 568=>x"6b00",
---- 569=>x"6e00", 570=>x"8a00", 571=>x"9e00", 572=>x"6c00",
---- 573=>x"7400", 574=>x"7700", 575=>x"8900", 576=>x"6e00",
---- 577=>x"7500", 578=>x"7500", 579=>x"6500", 580=>x"7e00",
---- 581=>x"8a00", 582=>x"8600", 583=>x"8b00", 584=>x"9b00",
---- 585=>x"9700", 586=>x"9200", 587=>x"9c00", 588=>x"8300",
---- 589=>x"7d00", 590=>x"7e00", 591=>x"7600", 592=>x"8300",
---- 593=>x"7800", 594=>x"6b00", 595=>x"6200", 596=>x"8200",
---- 597=>x"6d00", 598=>x"5500", 599=>x"4c00", 600=>x"7900",
---- 601=>x"5b00", 602=>x"4300", 603=>x"6e00", 604=>x"6e00",
---- 605=>x"5900", 606=>x"7c00", 607=>x"9700", 608=>x"8d00",
---- 609=>x"9100", 610=>x"8300", 611=>x"5d00", 612=>x"9500",
---- 613=>x"7200", 614=>x"2e00", 615=>x"2e00", 616=>x"8300",
---- 617=>x"5500", 618=>x"2c00", 619=>x"3c00", 620=>x"7d00",
---- 621=>x"5800", 622=>x"3800", 623=>x"5500", 624=>x"8200",
---- 625=>x"6500", 626=>x"3400", 627=>x"4300", 628=>x"8100",
---- 629=>x"5400", 630=>x"3a00", 631=>x"5200", 632=>x"6900",
---- 633=>x"4000", 634=>x"4a00", 635=>x"5e00", 636=>x"5f00",
---- 637=>x"4900", 638=>x"4200", 639=>x"5300", 640=>x"5a00",
---- 641=>x"4600", 642=>x"3b00", 643=>x"aa00", 644=>x"5700",
---- 645=>x"4a00", 646=>x"3f00", 647=>x"5b00", 648=>x"4a00",
---- 649=>x"5700", 650=>x"4a00", 651=>x"5c00", 652=>x"5400",
---- 653=>x"5e00", 654=>x"4800", 655=>x"5d00", 656=>x"5600",
---- 657=>x"4000", 658=>x"4300", 659=>x"5e00", 660=>x"4500",
---- 661=>x"2500", 662=>x"3700", 663=>x"5c00", 664=>x"5500",
---- 665=>x"2400", 666=>x"3400", 667=>x"5600", 668=>x"5400",
---- 669=>x"2f00", 670=>x"3a00", 671=>x"5a00", 672=>x"5300",
---- 673=>x"3900", 674=>x"3f00", 675=>x"4e00", 676=>x"4c00",
---- 677=>x"3d00", 678=>x"4300", 679=>x"4c00", 680=>x"4300",
---- 681=>x"3b00", 682=>x"4a00", 683=>x"6800", 684=>x"3d00",
---- 685=>x"b700", 686=>x"5d00", 687=>x"6400", 688=>x"4100",
---- 689=>x"5100", 690=>x"3600", 691=>x"5800", 692=>x"3f00",
---- 693=>x"3400", 694=>x"2900", 695=>x"6800", 696=>x"cb00",
---- 697=>x"2800", 698=>x"3f00", 699=>x"4f00", 700=>x"3600",
---- 701=>x"3600", 702=>x"5800", 703=>x"3400", 704=>x"3200",
---- 705=>x"4a00", 706=>x"4500", 707=>x"3300", 708=>x"3e00",
---- 709=>x"4500", 710=>x"3d00", 711=>x"3800", 712=>x"4300",
---- 713=>x"3a00", 714=>x"5700", 715=>x"4c00", 716=>x"4600",
---- 717=>x"3f00", 718=>x"7c00", 719=>x"5900", 720=>x"4000",
---- 721=>x"5700", 722=>x"8800", 723=>x"4700", 724=>x"2e00",
---- 725=>x"6600", 726=>x"8a00", 727=>x"3300", 728=>x"3600",
---- 729=>x"7a00", 730=>x"8700", 731=>x"2a00", 732=>x"4000",
---- 733=>x"7c00", 734=>x"7500", 735=>x"2c00", 736=>x"4300",
---- 737=>x"7800", 738=>x"5100", 739=>x"3000", 740=>x"4a00",
---- 741=>x"5b00", 742=>x"3c00", 743=>x"3400", 744=>x"5b00",
---- 745=>x"5200", 746=>x"3900", 747=>x"3200", 748=>x"5e00",
---- 749=>x"5400", 750=>x"3800", 751=>x"3400", 752=>x"6200",
---- 753=>x"5900", 754=>x"3200", 755=>x"3c00", 756=>x"7400",
---- 757=>x"5700", 758=>x"2d00", 759=>x"3d00", 760=>x"7500",
---- 761=>x"5d00", 762=>x"3000", 763=>x"3900", 764=>x"6400",
---- 765=>x"5600", 766=>x"3500", 767=>x"3800", 768=>x"4f00",
---- 769=>x"4600", 770=>x"3e00", 771=>x"3900", 772=>x"4c00",
---- 773=>x"3a00", 774=>x"4000", 775=>x"3c00", 776=>x"5600",
---- 777=>x"3500", 778=>x"3a00", 779=>x"4300", 780=>x"5900",
---- 781=>x"4200", 782=>x"3e00", 783=>x"4000", 784=>x"6000",
---- 785=>x"4800", 786=>x"3a00", 787=>x"3f00", 788=>x"6000",
---- 789=>x"4c00", 790=>x"3b00", 791=>x"3b00", 792=>x"5600",
---- 793=>x"4f00", 794=>x"2c00", 795=>x"3700", 796=>x"3a00",
---- 797=>x"5400", 798=>x"3f00", 799=>x"4400", 800=>x"2b00",
---- 801=>x"4000", 802=>x"6100", 803=>x"6600", 804=>x"2a00",
---- 805=>x"3100", 806=>x"5c00", 807=>x"7400", 808=>x"4200",
---- 809=>x"6500", 810=>x"6400", 811=>x"6700", 812=>x"d100",
---- 813=>x"6500", 814=>x"8100", 815=>x"8100", 816=>x"2700",
---- 817=>x"3a00", 818=>x"4800", 819=>x"4e00", 820=>x"3600",
---- 821=>x"4b00", 822=>x"3700", 823=>x"1e00", 824=>x"4300",
---- 825=>x"4b00", 826=>x"4100", 827=>x"2a00", 828=>x"4400",
---- 829=>x"4300", 830=>x"4400", 831=>x"3500", 832=>x"4700",
---- 833=>x"3700", 834=>x"3a00", 835=>x"3e00", 836=>x"5000",
---- 837=>x"2d00", 838=>x"3700", 839=>x"3600", 840=>x"4300",
---- 841=>x"2c00", 842=>x"3000", 843=>x"3600", 844=>x"3200",
---- 845=>x"2900", 846=>x"3000", 847=>x"3500", 848=>x"2c00",
---- 849=>x"2d00", 850=>x"3100", 851=>x"3200", 852=>x"2e00",
---- 853=>x"2e00", 854=>x"3000", 855=>x"3100", 856=>x"3300",
---- 857=>x"d100", 858=>x"3000", 859=>x"3200", 860=>x"2c00",
---- 861=>x"2900", 862=>x"3100", 863=>x"3400", 864=>x"2d00",
---- 865=>x"2900", 866=>x"3500", 867=>x"2d00", 868=>x"2a00",
---- 869=>x"2c00", 870=>x"3300", 871=>x"2500", 872=>x"2d00",
---- 873=>x"3100", 874=>x"2900", 875=>x"2500", 876=>x"2d00",
---- 877=>x"2f00", 878=>x"2800", 879=>x"2800", 880=>x"2e00",
---- 881=>x"2d00", 882=>x"3600", 883=>x"4200", 884=>x"2e00",
---- 885=>x"3b00", 886=>x"5d00", 887=>x"4400", 888=>x"2c00",
---- 889=>x"3d00", 890=>x"4c00", 891=>x"2c00", 892=>x"2b00",
---- 893=>x"3100", 894=>x"2f00", 895=>x"3300", 896=>x"2f00",
---- 897=>x"3200", 898=>x"2f00", 899=>x"c200", 900=>x"2c00",
---- 901=>x"3100", 902=>x"4400", 903=>x"4400", 904=>x"3c00",
---- 905=>x"5400", 906=>x"4800", 907=>x"3b00", 908=>x"5b00",
---- 909=>x"4c00", 910=>x"3200", 911=>x"2e00", 912=>x"3c00",
---- 913=>x"2b00", 914=>x"2d00", 915=>x"2c00", 916=>x"3200",
---- 917=>x"3100", 918=>x"2f00", 919=>x"3200", 920=>x"3000",
---- 921=>x"2c00", 922=>x"2e00", 923=>x"3700", 924=>x"3100",
---- 925=>x"2d00", 926=>x"2d00", 927=>x"3100", 928=>x"3100",
---- 929=>x"2f00", 930=>x"2f00", 931=>x"3a00", 932=>x"3000",
---- 933=>x"2f00", 934=>x"2e00", 935=>x"bc00", 936=>x"2c00",
---- 937=>x"2d00", 938=>x"3e00", 939=>x"4600", 940=>x"2b00",
---- 941=>x"4300", 942=>x"4800", 943=>x"3800", 944=>x"3900",
---- 945=>x"4700", 946=>x"3500", 947=>x"3500", 948=>x"3200",
---- 949=>x"2e00", 950=>x"3100", 951=>x"3900", 952=>x"2c00",
---- 953=>x"2d00", 954=>x"2f00", 955=>x"3a00", 956=>x"3200",
---- 957=>x"2d00", 958=>x"3100", 959=>x"3000", 960=>x"2e00",
---- 961=>x"2e00", 962=>x"3200", 963=>x"3700", 964=>x"3000",
---- 965=>x"2e00", 966=>x"3100", 967=>x"3a00", 968=>x"3800",
---- 969=>x"2d00", 970=>x"3000", 971=>x"3700", 972=>x"3a00",
---- 973=>x"2f00", 974=>x"3300", 975=>x"3b00", 976=>x"3c00",
---- 977=>x"d300", 978=>x"2f00", 979=>x"3500", 980=>x"3f00",
---- 981=>x"2f00", 982=>x"3000", 983=>x"2f00", 984=>x"3f00",
---- 985=>x"3100", 986=>x"3400", 987=>x"3000", 988=>x"3a00",
---- 989=>x"3600", 990=>x"3700", 991=>x"3600", 992=>x"4000",
---- 993=>x"3c00", 994=>x"3900", 995=>x"3500", 996=>x"c800",
---- 997=>x"3900", 998=>x"3900", 999=>x"3c00", 1000=>x"3500",
---- 1001=>x"3600", 1002=>x"3a00", 1003=>x"4200", 1004=>x"3600",
---- 1005=>x"3900", 1006=>x"3d00", 1007=>x"4300", 1008=>x"3800",
---- 1009=>x"3b00", 1010=>x"4000", 1011=>x"4200", 1012=>x"3d00",
---- 1013=>x"3f00", 1014=>x"5000", 1015=>x"4c00", 1016=>x"3d00",
---- 1017=>x"4300", 1018=>x"4b00", 1019=>x"4d00", 1020=>x"4000",
---- 1021=>x"4200", 1022=>x"4300", 1023=>x"4100"),
----
---- 12 => (0=>x"6d00", 1=>x"6d00", 2=>x"6800", 3=>x"6a00", 4=>x"6f00",
---- 5=>x"6d00", 6=>x"6900", 7=>x"6a00", 8=>x"6c00",
---- 9=>x"6c00", 10=>x"6900", 11=>x"6800", 12=>x"6a00",
---- 13=>x"6a00", 14=>x"6800", 15=>x"6b00", 16=>x"6700",
---- 17=>x"6a00", 18=>x"6800", 19=>x"6b00", 20=>x"6800",
---- 21=>x"6600", 22=>x"6700", 23=>x"6c00", 24=>x"6700",
---- 25=>x"6700", 26=>x"6500", 27=>x"6700", 28=>x"6900",
---- 29=>x"6500", 30=>x"6600", 31=>x"6800", 32=>x"6700",
---- 33=>x"6800", 34=>x"6500", 35=>x"6700", 36=>x"6500",
---- 37=>x"6700", 38=>x"6600", 39=>x"6900", 40=>x"6900",
---- 41=>x"6800", 42=>x"6600", 43=>x"6500", 44=>x"6600",
---- 45=>x"6700", 46=>x"6700", 47=>x"6900", 48=>x"6600",
---- 49=>x"6600", 50=>x"6800", 51=>x"6b00", 52=>x"6800",
---- 53=>x"6600", 54=>x"6700", 55=>x"6c00", 56=>x"6700",
---- 57=>x"6500", 58=>x"6800", 59=>x"6b00", 60=>x"6900",
---- 61=>x"6600", 62=>x"6600", 63=>x"6b00", 64=>x"6700",
---- 65=>x"6500", 66=>x"6800", 67=>x"6a00", 68=>x"6400",
---- 69=>x"6500", 70=>x"6600", 71=>x"6800", 72=>x"6600",
---- 73=>x"6800", 74=>x"6800", 75=>x"6900", 76=>x"6600",
---- 77=>x"6900", 78=>x"6500", 79=>x"6800", 80=>x"6600",
---- 81=>x"6600", 82=>x"6600", 83=>x"6700", 84=>x"6500",
---- 85=>x"6500", 86=>x"6700", 87=>x"6700", 88=>x"6700",
---- 89=>x"6500", 90=>x"6700", 91=>x"6800", 92=>x"6600",
---- 93=>x"6600", 94=>x"6800", 95=>x"6900", 96=>x"6500",
---- 97=>x"6500", 98=>x"6700", 99=>x"6a00", 100=>x"6700",
---- 101=>x"6500", 102=>x"6700", 103=>x"6a00", 104=>x"6900",
---- 105=>x"6900", 106=>x"6a00", 107=>x"6d00", 108=>x"6a00",
---- 109=>x"6700", 110=>x"6800", 111=>x"6b00", 112=>x"6800",
---- 113=>x"6800", 114=>x"6900", 115=>x"6800", 116=>x"6200",
---- 117=>x"6a00", 118=>x"6c00", 119=>x"9600", 120=>x"6500",
---- 121=>x"6800", 122=>x"6800", 123=>x"6a00", 124=>x"9800",
---- 125=>x"6400", 126=>x"6700", 127=>x"6900", 128=>x"6400",
---- 129=>x"6600", 130=>x"6900", 131=>x"6800", 132=>x"6400",
---- 133=>x"6600", 134=>x"6800", 135=>x"6700", 136=>x"6500",
---- 137=>x"6600", 138=>x"6300", 139=>x"6400", 140=>x"6500",
---- 141=>x"6500", 142=>x"6700", 143=>x"6800", 144=>x"6400",
---- 145=>x"6500", 146=>x"6100", 147=>x"6400", 148=>x"6300",
---- 149=>x"6300", 150=>x"6300", 151=>x"6700", 152=>x"6400",
---- 153=>x"6400", 154=>x"6600", 155=>x"6600", 156=>x"6500",
---- 157=>x"6500", 158=>x"6500", 159=>x"6800", 160=>x"6700",
---- 161=>x"6600", 162=>x"9b00", 163=>x"6700", 164=>x"6400",
---- 165=>x"6500", 166=>x"6600", 167=>x"6800", 168=>x"6300",
---- 169=>x"6500", 170=>x"6500", 171=>x"6700", 172=>x"6600",
---- 173=>x"6400", 174=>x"6400", 175=>x"6600", 176=>x"6600",
---- 177=>x"6300", 178=>x"6500", 179=>x"6600", 180=>x"6400",
---- 181=>x"6400", 182=>x"6300", 183=>x"6500", 184=>x"6200",
---- 185=>x"6200", 186=>x"6600", 187=>x"6700", 188=>x"6600",
---- 189=>x"6300", 190=>x"6300", 191=>x"6a00", 192=>x"6500",
---- 193=>x"6500", 194=>x"6400", 195=>x"6800", 196=>x"6300",
---- 197=>x"6300", 198=>x"6700", 199=>x"6800", 200=>x"6300",
---- 201=>x"6600", 202=>x"6800", 203=>x"6600", 204=>x"6500",
---- 205=>x"6800", 206=>x"6400", 207=>x"6600", 208=>x"6400",
---- 209=>x"6600", 210=>x"6200", 211=>x"6500", 212=>x"6200",
---- 213=>x"6100", 214=>x"6600", 215=>x"6300", 216=>x"6200",
---- 217=>x"6300", 218=>x"6500", 219=>x"6500", 220=>x"9b00",
---- 221=>x"6400", 222=>x"6500", 223=>x"6400", 224=>x"6600",
---- 225=>x"6400", 226=>x"6700", 227=>x"6b00", 228=>x"6000",
---- 229=>x"6500", 230=>x"6800", 231=>x"6d00", 232=>x"6300",
---- 233=>x"6300", 234=>x"6300", 235=>x"6700", 236=>x"6100",
---- 237=>x"6100", 238=>x"6300", 239=>x"6a00", 240=>x"6300",
---- 241=>x"6300", 242=>x"6400", 243=>x"6600", 244=>x"6300",
---- 245=>x"6400", 246=>x"6300", 247=>x"6600", 248=>x"6300",
---- 249=>x"6500", 250=>x"6300", 251=>x"6500", 252=>x"6500",
---- 253=>x"6400", 254=>x"6400", 255=>x"6700", 256=>x"6500",
---- 257=>x"6400", 258=>x"6800", 259=>x"6900", 260=>x"6400",
---- 261=>x"6400", 262=>x"6600", 263=>x"6c00", 264=>x"6700",
---- 265=>x"6500", 266=>x"6600", 267=>x"6900", 268=>x"6600",
---- 269=>x"6300", 270=>x"6300", 271=>x"6600", 272=>x"6700",
---- 273=>x"6200", 274=>x"6000", 275=>x"6600", 276=>x"6700",
---- 277=>x"6200", 278=>x"6300", 279=>x"6600", 280=>x"6500",
---- 281=>x"6400", 282=>x"6300", 283=>x"6400", 284=>x"6100",
---- 285=>x"6500", 286=>x"6400", 287=>x"6400", 288=>x"6000",
---- 289=>x"6200", 290=>x"6500", 291=>x"6600", 292=>x"6000",
---- 293=>x"6300", 294=>x"6300", 295=>x"6200", 296=>x"6200",
---- 297=>x"6200", 298=>x"6300", 299=>x"6300", 300=>x"6300",
---- 301=>x"6000", 302=>x"6200", 303=>x"6500", 304=>x"6100",
---- 305=>x"6400", 306=>x"6100", 307=>x"6300", 308=>x"6100",
---- 309=>x"6300", 310=>x"6200", 311=>x"6200", 312=>x"6200",
---- 313=>x"6200", 314=>x"6200", 315=>x"6400", 316=>x"6200",
---- 317=>x"6200", 318=>x"6200", 319=>x"6600", 320=>x"6400",
---- 321=>x"6100", 322=>x"6100", 323=>x"6300", 324=>x"6200",
---- 325=>x"6200", 326=>x"6100", 327=>x"6300", 328=>x"6200",
---- 329=>x"6200", 330=>x"6800", 331=>x"6600", 332=>x"6100",
---- 333=>x"6000", 334=>x"6300", 335=>x"6200", 336=>x"6200",
---- 337=>x"9e00", 338=>x"6200", 339=>x"6100", 340=>x"6300",
---- 341=>x"6200", 342=>x"6400", 343=>x"6200", 344=>x"6000",
---- 345=>x"6100", 346=>x"6200", 347=>x"6200", 348=>x"9d00",
---- 349=>x"6300", 350=>x"6000", 351=>x"9d00", 352=>x"6300",
---- 353=>x"6400", 354=>x"6200", 355=>x"6300", 356=>x"6300",
---- 357=>x"6400", 358=>x"6400", 359=>x"6100", 360=>x"6200",
---- 361=>x"5f00", 362=>x"6200", 363=>x"6200", 364=>x"6200",
---- 365=>x"6300", 366=>x"6400", 367=>x"6300", 368=>x"6400",
---- 369=>x"6100", 370=>x"6400", 371=>x"6400", 372=>x"6500",
---- 373=>x"6100", 374=>x"6500", 375=>x"6400", 376=>x"6500",
---- 377=>x"5d00", 378=>x"6100", 379=>x"6500", 380=>x"6500",
---- 381=>x"6100", 382=>x"6000", 383=>x"6400", 384=>x"6300",
---- 385=>x"6100", 386=>x"6300", 387=>x"6200", 388=>x"6200",
---- 389=>x"6300", 390=>x"6300", 391=>x"6100", 392=>x"6500",
---- 393=>x"6300", 394=>x"6200", 395=>x"6200", 396=>x"6000",
---- 397=>x"6000", 398=>x"6000", 399=>x"6400", 400=>x"5f00",
---- 401=>x"5d00", 402=>x"5f00", 403=>x"6100", 404=>x"6100",
---- 405=>x"6400", 406=>x"6000", 407=>x"6200", 408=>x"6000",
---- 409=>x"6300", 410=>x"5f00", 411=>x"6100", 412=>x"9b00",
---- 413=>x"6200", 414=>x"a100", 415=>x"6000", 416=>x"6100",
---- 417=>x"6300", 418=>x"6500", 419=>x"6500", 420=>x"6200",
---- 421=>x"6000", 422=>x"6400", 423=>x"6200", 424=>x"6000",
---- 425=>x"6300", 426=>x"6200", 427=>x"6300", 428=>x"6000",
---- 429=>x"6100", 430=>x"6100", 431=>x"6100", 432=>x"6300",
---- 433=>x"6300", 434=>x"6000", 435=>x"6000", 436=>x"6300",
---- 437=>x"6300", 438=>x"6300", 439=>x"6300", 440=>x"6200",
---- 441=>x"6200", 442=>x"6300", 443=>x"6500", 444=>x"6100",
---- 445=>x"6300", 446=>x"6300", 447=>x"6500", 448=>x"6500",
---- 449=>x"6600", 450=>x"6500", 451=>x"6500", 452=>x"6400",
---- 453=>x"6400", 454=>x"6300", 455=>x"6400", 456=>x"6500",
---- 457=>x"6100", 458=>x"6300", 459=>x"6300", 460=>x"6400",
---- 461=>x"6300", 462=>x"6300", 463=>x"6400", 464=>x"6300",
---- 465=>x"6800", 466=>x"6500", 467=>x"6700", 468=>x"6600",
---- 469=>x"6700", 470=>x"6600", 471=>x"6600", 472=>x"6500",
---- 473=>x"6700", 474=>x"6600", 475=>x"6600", 476=>x"6800",
---- 477=>x"6500", 478=>x"6400", 479=>x"6700", 480=>x"6700",
---- 481=>x"6600", 482=>x"6700", 483=>x"6900", 484=>x"6500",
---- 485=>x"6800", 486=>x"6800", 487=>x"6400", 488=>x"6400",
---- 489=>x"9a00", 490=>x"6400", 491=>x"6700", 492=>x"6800",
---- 493=>x"6200", 494=>x"6600", 495=>x"6700", 496=>x"6700",
---- 497=>x"6700", 498=>x"6700", 499=>x"6500", 500=>x"6500",
---- 501=>x"6600", 502=>x"6600", 503=>x"6400", 504=>x"5f00",
---- 505=>x"6300", 506=>x"6500", 507=>x"6600", 508=>x"6100",
---- 509=>x"6500", 510=>x"6400", 511=>x"6500", 512=>x"6400",
---- 513=>x"6500", 514=>x"9f00", 515=>x"6300", 516=>x"6200",
---- 517=>x"6000", 518=>x"6300", 519=>x"6100", 520=>x"6200",
---- 521=>x"6200", 522=>x"6000", 523=>x"5d00", 524=>x"6200",
---- 525=>x"5f00", 526=>x"5b00", 527=>x"5700", 528=>x"5f00",
---- 529=>x"5b00", 530=>x"5900", 531=>x"5900", 532=>x"5f00",
---- 533=>x"5d00", 534=>x"5a00", 535=>x"5b00", 536=>x"6300",
---- 537=>x"6300", 538=>x"6300", 539=>x"5700", 540=>x"7500",
---- 541=>x"6500", 542=>x"4700", 543=>x"4000", 544=>x"6000",
---- 545=>x"3800", 546=>x"3d00", 547=>x"3900", 548=>x"2a00",
---- 549=>x"2d00", 550=>x"5800", 551=>x"7800", 552=>x"3600",
---- 553=>x"4f00", 554=>x"8100", 555=>x"9e00", 556=>x"6600",
---- 557=>x"8500", 558=>x"a200", 559=>x"9b00", 560=>x"8a00",
---- 561=>x"8300", 562=>x"8600", 563=>x"9800", 564=>x"a200",
---- 565=>x"a300", 566=>x"9900", 567=>x"8600", 568=>x"a500",
---- 569=>x"8b00", 570=>x"7900", 571=>x"6c00", 572=>x"7600",
---- 573=>x"9700", 574=>x"6b00", 575=>x"5000", 576=>x"7600",
---- 577=>x"8b00", 578=>x"7200", 579=>x"7100", 580=>x"9e00",
---- 581=>x"ad00", 582=>x"9a00", 583=>x"8a00", 584=>x"9900",
---- 585=>x"7700", 586=>x"4600", 587=>x"3b00", 588=>x"5d00",
---- 589=>x"3d00", 590=>x"3400", 591=>x"4c00", 592=>x"5e00",
---- 593=>x"5900", 594=>x"5400", 595=>x"5a00", 596=>x"4c00",
---- 597=>x"5700", 598=>x"6900", 599=>x"5200", 600=>x"6f00",
---- 601=>x"7c00", 602=>x"a300", 603=>x"4b00", 604=>x"8800",
---- 605=>x"5c00", 606=>x"4200", 607=>x"6700", 608=>x"3b00",
---- 609=>x"4300", 610=>x"7100", 611=>x"8000", 612=>x"3800",
---- 613=>x"6a00", 614=>x"9c00", 615=>x"7200", 616=>x"6200",
---- 617=>x"8700", 618=>x"7700", 619=>x"5e00", 620=>x"8800",
---- 621=>x"7200", 622=>x"4d00", 623=>x"5f00", 624=>x"8a00",
---- 625=>x"5e00", 626=>x"5200", 627=>x"5c00", 628=>x"5b00",
---- 629=>x"4e00", 630=>x"6600", 631=>x"6500", 632=>x"4e00",
---- 633=>x"4900", 634=>x"7e00", 635=>x"6100", 636=>x"5300",
---- 637=>x"6b00", 638=>x"7a00", 639=>x"4e00", 640=>x"6400",
---- 641=>x"7000", 642=>x"6b00", 643=>x"5200", 644=>x"5d00",
---- 645=>x"7000", 646=>x"7900", 647=>x"5600", 648=>x"5700",
---- 649=>x"8700", 650=>x"7800", 651=>x"5200", 652=>x"5000",
---- 653=>x"5f00", 654=>x"5c00", 655=>x"4900", 656=>x"4c00",
---- 657=>x"4a00", 658=>x"4800", 659=>x"2900", 660=>x"5200",
---- 661=>x"4600", 662=>x"3900", 663=>x"2500", 664=>x"4700",
---- 665=>x"4500", 666=>x"3500", 667=>x"5300", 668=>x"4700",
---- 669=>x"4c00", 670=>x"6000", 671=>x"8600", 672=>x"4800",
---- 673=>x"7500", 674=>x"7c00", 675=>x"5a00", 676=>x"7100",
---- 677=>x"8600", 678=>x"3e00", 679=>x"2a00", 680=>x"7e00",
---- 681=>x"6c00", 682=>x"2800", 683=>x"2f00", 684=>x"7700",
---- 685=>x"5600", 686=>x"2e00", 687=>x"3900", 688=>x"6d00",
---- 689=>x"3d00", 690=>x"3500", 691=>x"3500", 692=>x"7a00",
---- 693=>x"4400", 694=>x"3700", 695=>x"3c00", 696=>x"5d00",
---- 697=>x"4d00", 698=>x"3600", 699=>x"3d00", 700=>x"3100",
---- 701=>x"4100", 702=>x"3f00", 703=>x"3f00", 704=>x"2700",
---- 705=>x"ca00", 706=>x"4600", 707=>x"b800", 708=>x"2f00",
---- 709=>x"3600", 710=>x"3400", 711=>x"3100", 712=>x"3a00",
---- 713=>x"2a00", 714=>x"2d00", 715=>x"2700", 716=>x"2d00",
---- 717=>x"2800", 718=>x"2d00", 719=>x"2d00", 720=>x"2e00",
---- 721=>x"3100", 722=>x"2b00", 723=>x"3600", 724=>x"2900",
---- 725=>x"3400", 726=>x"2c00", 727=>x"4900", 728=>x"3000",
---- 729=>x"3000", 730=>x"2400", 731=>x"5c00", 732=>x"2f00",
---- 733=>x"2c00", 734=>x"2f00", 735=>x"5e00", 736=>x"3100",
---- 737=>x"2400", 738=>x"3600", 739=>x"5a00", 740=>x"2e00",
---- 741=>x"2600", 742=>x"3a00", 743=>x"5c00", 744=>x"2900",
---- 745=>x"2600", 746=>x"4300", 747=>x"5c00", 748=>x"d600",
---- 749=>x"2500", 750=>x"4a00", 751=>x"5d00", 752=>x"3200",
---- 753=>x"2500", 754=>x"4600", 755=>x"5a00", 756=>x"3600",
---- 757=>x"2c00", 758=>x"4200", 759=>x"5500", 760=>x"3f00",
---- 761=>x"2f00", 762=>x"3e00", 763=>x"4c00", 764=>x"4400",
---- 765=>x"3c00", 766=>x"4300", 767=>x"4700", 768=>x"3f00",
---- 769=>x"3e00", 770=>x"4700", 771=>x"3f00", 772=>x"3800",
---- 773=>x"4300", 774=>x"3b00", 775=>x"3300", 776=>x"3800",
---- 777=>x"4600", 778=>x"3500", 779=>x"3100", 780=>x"4700",
---- 781=>x"3d00", 782=>x"3200", 783=>x"4200", 784=>x"4b00",
---- 785=>x"3800", 786=>x"3400", 787=>x"5100", 788=>x"3f00",
---- 789=>x"3600", 790=>x"3600", 791=>x"4e00", 792=>x"3e00",
---- 793=>x"3300", 794=>x"3400", 795=>x"4d00", 796=>x"3400",
---- 797=>x"2800", 798=>x"3100", 799=>x"4200", 800=>x"2900",
---- 801=>x"2100", 802=>x"3100", 803=>x"3b00", 804=>x"2500",
---- 805=>x"2100", 806=>x"2900", 807=>x"3200", 808=>x"2900",
---- 809=>x"1c00", 810=>x"2100", 811=>x"4b00", 812=>x"7100",
---- 813=>x"5b00", 814=>x"6700", 815=>x"8800", 816=>x"6400",
---- 817=>x"7500", 818=>x"7c00", 819=>x"6000", 820=>x"3100",
---- 821=>x"4c00", 822=>x"4100", 823=>x"3d00", 824=>x"3d00",
---- 825=>x"5800", 826=>x"4400", 827=>x"3a00", 828=>x"3300",
---- 829=>x"3c00", 830=>x"3300", 831=>x"2d00", 832=>x"2c00",
---- 833=>x"2f00", 834=>x"2b00", 835=>x"2900", 836=>x"3500",
---- 837=>x"2d00", 838=>x"2a00", 839=>x"3000", 840=>x"3800",
---- 841=>x"3100", 842=>x"2a00", 843=>x"3400", 844=>x"3200",
---- 845=>x"3100", 846=>x"2f00", 847=>x"3500", 848=>x"2a00",
---- 849=>x"2d00", 850=>x"2e00", 851=>x"3700", 852=>x"2d00",
---- 853=>x"2d00", 854=>x"2a00", 855=>x"3f00", 856=>x"3300",
---- 857=>x"3100", 858=>x"2b00", 859=>x"5300", 860=>x"3000",
---- 861=>x"d300", 862=>x"2e00", 863=>x"6e00", 864=>x"2600",
---- 865=>x"2600", 866=>x"3d00", 867=>x"7f00", 868=>x"2200",
---- 869=>x"2800", 870=>x"7300", 871=>x"8900", 872=>x"2800",
---- 873=>x"5a00", 874=>x"8500", 875=>x"6100", 876=>x"6000",
---- 877=>x"7800", 878=>x"4100", 879=>x"4b00", 880=>x"5900",
---- 881=>x"3a00", 882=>x"2400", 883=>x"6400", 884=>x"2d00",
---- 885=>x"2a00", 886=>x"3300", 887=>x"5a00", 888=>x"2f00",
---- 889=>x"3400", 890=>x"3200", 891=>x"5000", 892=>x"3b00",
---- 893=>x"3400", 894=>x"2c00", 895=>x"4c00", 896=>x"3900",
---- 897=>x"2d00", 898=>x"3300", 899=>x"4600", 900=>x"3200",
---- 901=>x"3000", 902=>x"3100", 903=>x"3f00", 904=>x"2f00",
---- 905=>x"2d00", 906=>x"2e00", 907=>x"3f00", 908=>x"2a00",
---- 909=>x"2c00", 910=>x"3a00", 911=>x"4200", 912=>x"2b00",
---- 913=>x"2c00", 914=>x"4100", 915=>x"3d00", 916=>x"2d00",
---- 917=>x"3300", 918=>x"3d00", 919=>x"3d00", 920=>x"2c00",
---- 921=>x"3d00", 922=>x"3900", 923=>x"4000", 924=>x"3600",
---- 925=>x"4300", 926=>x"3700", 927=>x"4500", 928=>x"4400",
---- 929=>x"3500", 930=>x"3a00", 931=>x"4100", 932=>x"3f00",
---- 933=>x"2d00", 934=>x"3e00", 935=>x"3d00", 936=>x"3300",
---- 937=>x"d200", 938=>x"4100", 939=>x"3d00", 940=>x"2e00",
---- 941=>x"2c00", 942=>x"4700", 943=>x"3d00", 944=>x"3600",
---- 945=>x"2d00", 946=>x"3f00", 947=>x"3800", 948=>x"3300",
---- 949=>x"2c00", 950=>x"3400", 951=>x"3e00", 952=>x"3300",
---- 953=>x"3100", 954=>x"3100", 955=>x"3d00", 956=>x"3200",
---- 957=>x"3100", 958=>x"3200", 959=>x"3300", 960=>x"3a00",
---- 961=>x"3100", 962=>x"3200", 963=>x"2b00", 964=>x"3c00",
---- 965=>x"3000", 966=>x"3300", 967=>x"3300", 968=>x"3a00",
---- 969=>x"2d00", 970=>x"3100", 971=>x"3000", 972=>x"3c00",
---- 973=>x"3000", 974=>x"2b00", 975=>x"2c00", 976=>x"4800",
---- 977=>x"4000", 978=>x"2b00", 979=>x"2d00", 980=>x"4800",
---- 981=>x"3e00", 982=>x"d400", 983=>x"3400", 984=>x"4f00",
---- 985=>x"3e00", 986=>x"2800", 987=>x"3300", 988=>x"5400",
---- 989=>x"4800", 990=>x"2900", 991=>x"3500", 992=>x"4700",
---- 993=>x"5900", 994=>x"2a00", 995=>x"2f00", 996=>x"3500",
---- 997=>x"5800", 998=>x"3900", 999=>x"2c00", 1000=>x"d000",
---- 1001=>x"4d00", 1002=>x"5300", 1003=>x"2900", 1004=>x"3400",
---- 1005=>x"3700", 1006=>x"5c00", 1007=>x"2f00", 1008=>x"3f00",
---- 1009=>x"2800", 1010=>x"5400", 1011=>x"4800", 1012=>x"4a00",
---- 1013=>x"3400", 1014=>x"3b00", 1015=>x"4e00", 1016=>x"4f00",
---- 1017=>x"3900", 1018=>x"3000", 1019=>x"4300", 1020=>x"4c00",
---- 1021=>x"4400", 1022=>x"3200", 1023=>x"4c00"),
----
---- 13 => (0=>x"9200", 1=>x"7000", 2=>x"7100", 3=>x"7800", 4=>x"6e00",
---- 5=>x"7200", 6=>x"7100", 7=>x"7800", 8=>x"6d00",
---- 9=>x"7200", 10=>x"7200", 11=>x"7700", 12=>x"6b00",
---- 13=>x"6e00", 14=>x"7400", 15=>x"7500", 16=>x"6e00",
---- 17=>x"6e00", 18=>x"7000", 19=>x"7400", 20=>x"6e00",
---- 21=>x"6d00", 22=>x"7200", 23=>x"7400", 24=>x"7000",
---- 25=>x"8f00", 26=>x"7100", 27=>x"7400", 28=>x"6e00",
---- 29=>x"6e00", 30=>x"7000", 31=>x"7400", 32=>x"6b00",
---- 33=>x"6f00", 34=>x"7000", 35=>x"7400", 36=>x"9200",
---- 37=>x"7100", 38=>x"7300", 39=>x"7500", 40=>x"6e00",
---- 41=>x"7100", 42=>x"7300", 43=>x"7100", 44=>x"6d00",
---- 45=>x"6f00", 46=>x"6f00", 47=>x"7300", 48=>x"6b00",
---- 49=>x"6e00", 50=>x"6f00", 51=>x"6f00", 52=>x"6e00",
---- 53=>x"6d00", 54=>x"6f00", 55=>x"7200", 56=>x"6b00",
---- 57=>x"6c00", 58=>x"7100", 59=>x"7300", 60=>x"6c00",
---- 61=>x"6b00", 62=>x"6e00", 63=>x"7300", 64=>x"6b00",
---- 65=>x"6e00", 66=>x"7100", 67=>x"7100", 68=>x"6b00",
---- 69=>x"6f00", 70=>x"6f00", 71=>x"7200", 72=>x"6b00",
---- 73=>x"6e00", 74=>x"7200", 75=>x"7000", 76=>x"6b00",
---- 77=>x"6e00", 78=>x"7000", 79=>x"7300", 80=>x"6900",
---- 81=>x"6f00", 82=>x"7200", 83=>x"7400", 84=>x"6900",
---- 85=>x"6d00", 86=>x"6f00", 87=>x"7100", 88=>x"6d00",
---- 89=>x"6c00", 90=>x"6f00", 91=>x"7400", 92=>x"7000",
---- 93=>x"6c00", 94=>x"7200", 95=>x"7500", 96=>x"6f00",
---- 97=>x"7000", 98=>x"7000", 99=>x"6f00", 100=>x"6e00",
---- 101=>x"7200", 102=>x"7100", 103=>x"7100", 104=>x"6c00",
---- 105=>x"6f00", 106=>x"7100", 107=>x"7400", 108=>x"6d00",
---- 109=>x"7100", 110=>x"7700", 111=>x"7300", 112=>x"6c00",
---- 113=>x"6f00", 114=>x"7700", 115=>x"7300", 116=>x"6a00",
---- 117=>x"6e00", 118=>x"7100", 119=>x"7100", 120=>x"6b00",
---- 121=>x"6e00", 122=>x"7000", 123=>x"7100", 124=>x"6b00",
---- 125=>x"6e00", 126=>x"6e00", 127=>x"7200", 128=>x"6900",
---- 129=>x"6d00", 130=>x"6c00", 131=>x"6f00", 132=>x"6700",
---- 133=>x"6a00", 134=>x"6600", 135=>x"6d00", 136=>x"6900",
---- 137=>x"6a00", 138=>x"6c00", 139=>x"6f00", 140=>x"6b00",
---- 141=>x"6c00", 142=>x"6c00", 143=>x"6f00", 144=>x"6800",
---- 145=>x"6b00", 146=>x"6d00", 147=>x"6d00", 148=>x"6900",
---- 149=>x"6a00", 150=>x"6d00", 151=>x"6d00", 152=>x"6800",
---- 153=>x"6800", 154=>x"6c00", 155=>x"6e00", 156=>x"6700",
---- 157=>x"6a00", 158=>x"6e00", 159=>x"7000", 160=>x"6a00",
---- 161=>x"6c00", 162=>x"6d00", 163=>x"6e00", 164=>x"6900",
---- 165=>x"6b00", 166=>x"6e00", 167=>x"6e00", 168=>x"6600",
---- 169=>x"6900", 170=>x"7000", 171=>x"7000", 172=>x"6700",
---- 173=>x"6a00", 174=>x"6b00", 175=>x"6e00", 176=>x"6900",
---- 177=>x"6d00", 178=>x"9200", 179=>x"6c00", 180=>x"6b00",
---- 181=>x"6e00", 182=>x"6c00", 183=>x"6c00", 184=>x"6a00",
---- 185=>x"6600", 186=>x"6b00", 187=>x"6e00", 188=>x"6900",
---- 189=>x"6700", 190=>x"6b00", 191=>x"6e00", 192=>x"6500",
---- 193=>x"6700", 194=>x"6b00", 195=>x"6f00", 196=>x"9800",
---- 197=>x"6a00", 198=>x"6900", 199=>x"6d00", 200=>x"6700",
---- 201=>x"6a00", 202=>x"6e00", 203=>x"6d00", 204=>x"6600",
---- 205=>x"6a00", 206=>x"6d00", 207=>x"6f00", 208=>x"6700",
---- 209=>x"6900", 210=>x"6d00", 211=>x"6e00", 212=>x"6700",
---- 213=>x"6a00", 214=>x"6b00", 215=>x"6e00", 216=>x"6700",
---- 217=>x"6800", 218=>x"6a00", 219=>x"6e00", 220=>x"6b00",
---- 221=>x"6c00", 222=>x"6d00", 223=>x"6d00", 224=>x"6d00",
---- 225=>x"6a00", 226=>x"6e00", 227=>x"6f00", 228=>x"6c00",
---- 229=>x"6b00", 230=>x"6b00", 231=>x"6c00", 232=>x"6400",
---- 233=>x"6900", 234=>x"6b00", 235=>x"6e00", 236=>x"6700",
---- 237=>x"6800", 238=>x"6900", 239=>x"6a00", 240=>x"6800",
---- 241=>x"9700", 242=>x"6b00", 243=>x"6b00", 244=>x"6800",
---- 245=>x"6800", 246=>x"6900", 247=>x"6900", 248=>x"6800",
---- 249=>x"6800", 250=>x"6a00", 251=>x"6a00", 252=>x"6500",
---- 253=>x"6900", 254=>x"6d00", 255=>x"6f00", 256=>x"6a00",
---- 257=>x"6900", 258=>x"6d00", 259=>x"6d00", 260=>x"6900",
---- 261=>x"6a00", 262=>x"6d00", 263=>x"6c00", 264=>x"6c00",
---- 265=>x"6c00", 266=>x"6e00", 267=>x"6e00", 268=>x"6d00",
---- 269=>x"6f00", 270=>x"6d00", 271=>x"6e00", 272=>x"9300",
---- 273=>x"6900", 274=>x"6c00", 275=>x"6e00", 276=>x"6500",
---- 277=>x"6a00", 278=>x"6c00", 279=>x"6c00", 280=>x"6600",
---- 281=>x"6a00", 282=>x"6a00", 283=>x"6c00", 284=>x"6600",
---- 285=>x"6b00", 286=>x"6c00", 287=>x"6c00", 288=>x"6600",
---- 289=>x"6800", 290=>x"6900", 291=>x"6900", 292=>x"6500",
---- 293=>x"6500", 294=>x"6700", 295=>x"6a00", 296=>x"6300",
---- 297=>x"6500", 298=>x"6a00", 299=>x"6900", 300=>x"6400",
---- 301=>x"6600", 302=>x"6d00", 303=>x"6900", 304=>x"6600",
---- 305=>x"6700", 306=>x"6700", 307=>x"6800", 308=>x"6500",
---- 309=>x"6800", 310=>x"6600", 311=>x"6a00", 312=>x"6300",
---- 313=>x"6600", 314=>x"6500", 315=>x"6700", 316=>x"6300",
---- 317=>x"6500", 318=>x"6800", 319=>x"6600", 320=>x"6500",
---- 321=>x"6500", 322=>x"6700", 323=>x"6600", 324=>x"6600",
---- 325=>x"9b00", 326=>x"6400", 327=>x"6200", 328=>x"6400",
---- 329=>x"6400", 330=>x"6400", 331=>x"6200", 332=>x"6200",
---- 333=>x"6100", 334=>x"6400", 335=>x"6500", 336=>x"6200",
---- 337=>x"6200", 338=>x"6500", 339=>x"6200", 340=>x"6000",
---- 341=>x"6200", 342=>x"6200", 343=>x"5e00", 344=>x"6600",
---- 345=>x"6400", 346=>x"6400", 347=>x"6000", 348=>x"6200",
---- 349=>x"6300", 350=>x"5f00", 351=>x"5f00", 352=>x"6500",
---- 353=>x"6200", 354=>x"6100", 355=>x"5f00", 356=>x"6400",
---- 357=>x"6300", 358=>x"6300", 359=>x"5e00", 360=>x"6400",
---- 361=>x"6400", 362=>x"6100", 363=>x"5f00", 364=>x"6400",
---- 365=>x"6500", 366=>x"6600", 367=>x"6100", 368=>x"6500",
---- 369=>x"6200", 370=>x"6200", 371=>x"6000", 372=>x"6300",
---- 373=>x"6100", 374=>x"6200", 375=>x"6000", 376=>x"6300",
---- 377=>x"6100", 378=>x"5f00", 379=>x"a200", 380=>x"6400",
---- 381=>x"6000", 382=>x"6000", 383=>x"6200", 384=>x"6700",
---- 385=>x"6400", 386=>x"6400", 387=>x"6300", 388=>x"6100",
---- 389=>x"6200", 390=>x"6400", 391=>x"6500", 392=>x"6100",
---- 393=>x"6000", 394=>x"6000", 395=>x"6500", 396=>x"6200",
---- 397=>x"6100", 398=>x"9a00", 399=>x"6600", 400=>x"6000",
---- 401=>x"5f00", 402=>x"6600", 403=>x"6800", 404=>x"6200",
---- 405=>x"6100", 406=>x"6600", 407=>x"6800", 408=>x"6300",
---- 409=>x"6000", 410=>x"6700", 411=>x"6800", 412=>x"6300",
---- 413=>x"6500", 414=>x"6800", 415=>x"6900", 416=>x"6400",
---- 417=>x"6600", 418=>x"6800", 419=>x"6700", 420=>x"6100",
---- 421=>x"6700", 422=>x"6b00", 423=>x"6800", 424=>x"6400",
---- 425=>x"6400", 426=>x"6700", 427=>x"6c00", 428=>x"6600",
---- 429=>x"6400", 430=>x"6900", 431=>x"6700", 432=>x"6300",
---- 433=>x"6400", 434=>x"6900", 435=>x"6800", 436=>x"6200",
---- 437=>x"6700", 438=>x"6900", 439=>x"6a00", 440=>x"6400",
---- 441=>x"6900", 442=>x"6b00", 443=>x"6a00", 444=>x"6800",
---- 445=>x"6700", 446=>x"6800", 447=>x"6e00", 448=>x"6600",
---- 449=>x"6800", 450=>x"6400", 451=>x"9b00", 452=>x"6300",
---- 453=>x"6400", 454=>x"6300", 455=>x"7700", 456=>x"6300",
---- 457=>x"6300", 458=>x"6d00", 459=>x"9600", 460=>x"6800",
---- 461=>x"6700", 462=>x"7200", 463=>x"7700", 464=>x"6800",
---- 465=>x"6800", 466=>x"6d00", 467=>x"7800", 468=>x"6500",
---- 469=>x"6700", 470=>x"6a00", 471=>x"7f00", 472=>x"6800",
---- 473=>x"6b00", 474=>x"6b00", 475=>x"7200", 476=>x"6a00",
---- 477=>x"6b00", 478=>x"6c00", 479=>x"7000", 480=>x"6800",
---- 481=>x"6b00", 482=>x"6d00", 483=>x"6e00", 484=>x"6800",
---- 485=>x"6b00", 486=>x"6f00", 487=>x"7000", 488=>x"6900",
---- 489=>x"6b00", 490=>x"6f00", 491=>x"7200", 492=>x"6900",
---- 493=>x"6900", 494=>x"6d00", 495=>x"7100", 496=>x"6600",
---- 497=>x"6800", 498=>x"6b00", 499=>x"7400", 500=>x"6700",
---- 501=>x"6b00", 502=>x"6d00", 503=>x"7100", 504=>x"6700",
---- 505=>x"6800", 506=>x"6a00", 507=>x"6b00", 508=>x"6500",
---- 509=>x"6500", 510=>x"6b00", 511=>x"6c00", 512=>x"6700",
---- 513=>x"6600", 514=>x"6800", 515=>x"6900", 516=>x"6000",
---- 517=>x"6200", 518=>x"6500", 519=>x"8100", 520=>x"5b00",
---- 521=>x"5c00", 522=>x"7d00", 523=>x"a000", 524=>x"5000",
---- 525=>x"7700", 526=>x"c000", 527=>x"ba00", 528=>x"4f00",
---- 529=>x"8f00", 530=>x"ca00", 531=>x"c000", 532=>x"4c00",
---- 533=>x"6b00", 534=>x"b700", 535=>x"ba00", 536=>x"3200",
---- 537=>x"5100", 538=>x"ad00", 539=>x"6800", 540=>x"2c00",
---- 541=>x"2c00", 542=>x"9100", 543=>x"7a00", 544=>x"3d00",
---- 545=>x"5600", 546=>x"9500", 547=>x"a000", 548=>x"8400",
---- 549=>x"9a00", 550=>x"ac00", 551=>x"bb00", 552=>x"9600",
---- 553=>x"9800", 554=>x"9500", 555=>x"a500", 556=>x"8300",
---- 557=>x"8700", 558=>x"7d00", 559=>x"9700", 560=>x"8600",
---- 561=>x"6800", 562=>x"5100", 563=>x"5700", 564=>x"5f00",
---- 565=>x"4500", 566=>x"4100", 567=>x"4100", 568=>x"4700",
---- 569=>x"3900", 570=>x"4500", 571=>x"6300", 572=>x"4300",
---- 573=>x"4f00", 574=>x"6400", 575=>x"5c00", 576=>x"9100",
---- 577=>x"9100", 578=>x"7200", 579=>x"4200", 580=>x"7f00",
---- 581=>x"6a00", 582=>x"4c00", 583=>x"3d00", 584=>x"4800",
---- 585=>x"4d00", 586=>x"3700", 587=>x"3b00", 588=>x"aa00",
---- 589=>x"3f00", 590=>x"3a00", 591=>x"3e00", 592=>x"4e00",
---- 593=>x"3e00", 594=>x"3f00", 595=>x"3400", 596=>x"5700",
---- 597=>x"5300", 598=>x"3800", 599=>x"3900", 600=>x"7500",
---- 601=>x"5b00", 602=>x"4100", 603=>x"5e00", 604=>x"6a00",
---- 605=>x"4400", 606=>x"6100", 607=>x"7a00", 608=>x"4b00",
---- 609=>x"5f00", 610=>x"7e00", 611=>x"3e00", 612=>x"5900",
---- 613=>x"7600", 614=>x"4200", 615=>x"2f00", 616=>x"6f00",
---- 617=>x"3c00", 618=>x"3a00", 619=>x"3600", 620=>x"5100",
---- 621=>x"5e00", 622=>x"4500", 623=>x"c500", 624=>x"5900",
---- 625=>x"4a00", 626=>x"4000", 627=>x"5d00", 628=>x"5800",
---- 629=>x"4100", 630=>x"5e00", 631=>x"5600", 632=>x"4400",
---- 633=>x"5700", 634=>x"4e00", 635=>x"3b00", 636=>x"5500",
---- 637=>x"4a00", 638=>x"4a00", 639=>x"3300", 640=>x"4a00",
---- 641=>x"3700", 642=>x"3b00", 643=>x"5000", 644=>x"4800",
---- 645=>x"2900", 646=>x"3200", 647=>x"8a00", 648=>x"3d00",
---- 649=>x"1e00", 650=>x"4c00", 651=>x"9200", 652=>x"2b00",
---- 653=>x"3100", 654=>x"8100", 655=>x"7a00", 656=>x"2b00",
---- 657=>x"7000", 658=>x"7e00", 659=>x"4e00", 660=>x"5d00",
---- 661=>x"7b00", 662=>x"4600", 663=>x"3200", 664=>x"8900",
---- 665=>x"4e00", 666=>x"2c00", 667=>x"3100", 668=>x"5c00",
---- 669=>x"3900", 670=>x"3100", 671=>x"3300", 672=>x"3800",
---- 673=>x"3300", 674=>x"2f00", 675=>x"3000", 676=>x"4900",
---- 677=>x"3a00", 678=>x"3800", 679=>x"3200", 680=>x"4500",
---- 681=>x"4c00", 682=>x"4500", 683=>x"3a00", 684=>x"3400",
---- 685=>x"4e00", 686=>x"4500", 687=>x"b800", 688=>x"4400",
---- 689=>x"4300", 690=>x"3a00", 691=>x"4d00", 692=>x"4100",
---- 693=>x"4100", 694=>x"3700", 695=>x"4600", 696=>x"4000",
---- 697=>x"4200", 698=>x"3900", 699=>x"3400", 700=>x"4200",
---- 701=>x"4d00", 702=>x"3b00", 703=>x"3500", 704=>x"4400",
---- 705=>x"4500", 706=>x"3c00", 707=>x"4900", 708=>x"4600",
---- 709=>x"4500", 710=>x"3b00", 711=>x"5700", 712=>x"4900",
---- 713=>x"5100", 714=>x"3400", 715=>x"5a00", 716=>x"5d00",
---- 717=>x"4f00", 718=>x"3600", 719=>x"5400", 720=>x"6400",
---- 721=>x"4400", 722=>x"5100", 723=>x"4900", 724=>x"6700",
---- 725=>x"3300", 726=>x"5100", 727=>x"5500", 728=>x"5b00",
---- 729=>x"3100", 730=>x"3600", 731=>x"5700", 732=>x"4600",
---- 733=>x"3500", 734=>x"2a00", 735=>x"3b00", 736=>x"3f00",
---- 737=>x"3e00", 738=>x"3700", 739=>x"2600", 740=>x"3700",
---- 741=>x"3f00", 742=>x"3d00", 743=>x"3300", 744=>x"2e00",
---- 745=>x"3300", 746=>x"4100", 747=>x"2d00", 748=>x"3000",
---- 749=>x"2e00", 750=>x"3d00", 751=>x"3c00", 752=>x"2e00",
---- 753=>x"3300", 754=>x"3900", 755=>x"4500", 756=>x"3000",
---- 757=>x"3700", 758=>x"3600", 759=>x"3a00", 760=>x"3000",
---- 761=>x"3200", 762=>x"3200", 763=>x"2b00", 764=>x"3300",
---- 765=>x"2d00", 766=>x"3500", 767=>x"2400", 768=>x"3300",
---- 769=>x"2a00", 770=>x"3900", 771=>x"2600", 772=>x"3400",
---- 773=>x"2d00", 774=>x"3300", 775=>x"2900", 776=>x"3000",
---- 777=>x"2e00", 778=>x"3000", 779=>x"2800", 780=>x"3300",
---- 781=>x"2b00", 782=>x"3100", 783=>x"2d00", 784=>x"4100",
---- 785=>x"2f00", 786=>x"3600", 787=>x"2f00", 788=>x"5d00",
---- 789=>x"c700", 790=>x"3800", 791=>x"3200", 792=>x"7000",
---- 793=>x"4600", 794=>x"3d00", 795=>x"3f00", 796=>x"6c00",
---- 797=>x"5400", 798=>x"4400", 799=>x"4100", 800=>x"6a00",
---- 801=>x"6400", 802=>x"4d00", 803=>x"4800", 804=>x"7000",
---- 805=>x"7000", 806=>x"4500", 807=>x"5b00", 808=>x"8c00",
---- 809=>x"6200", 810=>x"4400", 811=>x"6600", 812=>x"6d00",
---- 813=>x"4300", 814=>x"4800", 815=>x"4a00", 816=>x"4200",
---- 817=>x"5200", 818=>x"4300", 819=>x"3b00", 820=>x"3c00",
---- 821=>x"c700", 822=>x"3a00", 823=>x"4900", 824=>x"3b00",
---- 825=>x"3900", 826=>x"c300", 827=>x"3900", 828=>x"4400",
---- 829=>x"aa00", 830=>x"4300", 831=>x"3900", 832=>x"5100",
---- 833=>x"6a00", 834=>x"4300", 835=>x"3b00", 836=>x"6100",
---- 837=>x"6a00", 838=>x"3600", 839=>x"4800", 840=>x"6c00",
---- 841=>x"6b00", 842=>x"2d00", 843=>x"4000", 844=>x"7100",
---- 845=>x"7300", 846=>x"3000", 847=>x"3600", 848=>x"7400",
---- 849=>x"7000", 850=>x"2d00", 851=>x"3700", 852=>x"8500",
---- 853=>x"6c00", 854=>x"2200", 855=>x"3300", 856=>x"9400",
---- 857=>x"6600", 858=>x"2600", 859=>x"2500", 860=>x"9500",
---- 861=>x"5b00", 862=>x"2700", 863=>x"dd00", 864=>x"8800",
---- 865=>x"5400", 866=>x"2a00", 867=>x"2c00", 868=>x"7f00",
---- 869=>x"5800", 870=>x"2b00", 871=>x"2900", 872=>x"7000",
---- 873=>x"3f00", 874=>x"2800", 875=>x"2900", 876=>x"6a00",
---- 877=>x"3c00", 878=>x"3100", 879=>x"2a00", 880=>x"6600",
---- 881=>x"4b00", 882=>x"3600", 883=>x"2d00", 884=>x"5600",
---- 885=>x"5700", 886=>x"3600", 887=>x"3000", 888=>x"5600",
---- 889=>x"5500", 890=>x"3800", 891=>x"2e00", 892=>x"5300",
---- 893=>x"4300", 894=>x"3900", 895=>x"3100", 896=>x"4700",
---- 897=>x"3b00", 898=>x"3100", 899=>x"3500", 900=>x"4300",
---- 901=>x"3d00", 902=>x"3d00", 903=>x"3d00", 904=>x"3c00",
---- 905=>x"3800", 906=>x"4000", 907=>x"3700", 908=>x"3e00",
---- 909=>x"3b00", 910=>x"3100", 911=>x"2d00", 912=>x"4200",
---- 913=>x"3500", 914=>x"3200", 915=>x"3800", 916=>x"4900",
---- 917=>x"3a00", 918=>x"3300", 919=>x"3d00", 920=>x"3b00",
---- 921=>x"3600", 922=>x"3700", 923=>x"4d00", 924=>x"3400",
---- 925=>x"3200", 926=>x"3c00", 927=>x"5100", 928=>x"3200",
---- 929=>x"3200", 930=>x"3c00", 931=>x"3f00", 932=>x"3000",
---- 933=>x"cb00", 934=>x"4000", 935=>x"4100", 936=>x"2e00",
---- 937=>x"2f00", 938=>x"3d00", 939=>x"4300", 940=>x"2e00",
---- 941=>x"3100", 942=>x"3f00", 943=>x"3e00", 944=>x"2a00",
---- 945=>x"3600", 946=>x"4900", 947=>x"3b00", 948=>x"2e00",
---- 949=>x"3700", 950=>x"4500", 951=>x"3d00", 952=>x"3500",
---- 953=>x"3f00", 954=>x"3e00", 955=>x"3800", 956=>x"3800",
---- 957=>x"4600", 958=>x"3400", 959=>x"3b00", 960=>x"3200",
---- 961=>x"3400", 962=>x"2f00", 963=>x"4000", 964=>x"2d00",
---- 965=>x"2800", 966=>x"3400", 967=>x"3f00", 968=>x"2d00",
---- 969=>x"3700", 970=>x"4500", 971=>x"4500", 972=>x"2e00",
---- 973=>x"3900", 974=>x"5100", 975=>x"4e00", 976=>x"2e00",
---- 977=>x"3900", 978=>x"4c00", 979=>x"5100", 980=>x"2e00",
---- 981=>x"3e00", 982=>x"4800", 983=>x"4d00", 984=>x"3000",
---- 985=>x"3c00", 986=>x"3c00", 987=>x"5000", 988=>x"3000",
---- 989=>x"3b00", 990=>x"3f00", 991=>x"5b00", 992=>x"2f00",
---- 993=>x"3700", 994=>x"4e00", 995=>x"5f00", 996=>x"2c00",
---- 997=>x"2e00", 998=>x"4e00", 999=>x"5c00", 1000=>x"2e00",
---- 1001=>x"2b00", 1002=>x"6000", 1003=>x"6800", 1004=>x"2700",
---- 1005=>x"3000", 1006=>x"7600", 1007=>x"6c00", 1008=>x"2800",
---- 1009=>x"3300", 1010=>x"8000", 1011=>x"5b00", 1012=>x"3300",
---- 1013=>x"3e00", 1014=>x"7c00", 1015=>x"4d00", 1016=>x"4100",
---- 1017=>x"5e00", 1018=>x"7f00", 1019=>x"3400", 1020=>x"5600",
---- 1021=>x"7e00", 1022=>x"6d00", 1023=>x"2e00"),
----
---- 14 => (0=>x"7400", 1=>x"8500", 2=>x"7c00", 3=>x"7900", 4=>x"7500",
---- 5=>x"7a00", 6=>x"7a00", 7=>x"7900", 8=>x"7500",
---- 9=>x"7900", 10=>x"7b00", 11=>x"7a00", 12=>x"8900",
---- 13=>x"7900", 14=>x"7d00", 15=>x"7c00", 16=>x"7700",
---- 17=>x"7a00", 18=>x"7a00", 19=>x"7c00", 20=>x"7400",
---- 21=>x"7900", 22=>x"7b00", 23=>x"7c00", 24=>x"7700",
---- 25=>x"7500", 26=>x"7a00", 27=>x"7a00", 28=>x"7600",
---- 29=>x"7600", 30=>x"7a00", 31=>x"7800", 32=>x"7300",
---- 33=>x"7800", 34=>x"7a00", 35=>x"7d00", 36=>x"7700",
---- 37=>x"7700", 38=>x"7800", 39=>x"7a00", 40=>x"7700",
---- 41=>x"7800", 42=>x"7800", 43=>x"7700", 44=>x"7400",
---- 45=>x"7600", 46=>x"7700", 47=>x"7900", 48=>x"7500",
---- 49=>x"7900", 50=>x"7a00", 51=>x"7800", 52=>x"7700",
---- 53=>x"7900", 54=>x"7700", 55=>x"7a00", 56=>x"7500",
---- 57=>x"7a00", 58=>x"7800", 59=>x"7800", 60=>x"7400",
---- 61=>x"7600", 62=>x"7a00", 63=>x"7a00", 64=>x"7500",
---- 65=>x"7700", 66=>x"7a00", 67=>x"7900", 68=>x"7400",
---- 69=>x"7500", 70=>x"7800", 71=>x"7a00", 72=>x"7700",
---- 73=>x"7400", 74=>x"7800", 75=>x"7800", 76=>x"7300",
---- 77=>x"7300", 78=>x"7900", 79=>x"7900", 80=>x"7400",
---- 81=>x"7700", 82=>x"7700", 83=>x"7900", 84=>x"7500",
---- 85=>x"7a00", 86=>x"7800", 87=>x"7700", 88=>x"7500",
---- 89=>x"7800", 90=>x"7800", 91=>x"7800", 92=>x"7500",
---- 93=>x"7800", 94=>x"7800", 95=>x"7900", 96=>x"7200",
---- 97=>x"7700", 98=>x"7900", 99=>x"7a00", 100=>x"7400",
---- 101=>x"7900", 102=>x"7900", 103=>x"7900", 104=>x"7600",
---- 105=>x"7800", 106=>x"7900", 107=>x"7b00", 108=>x"7500",
---- 109=>x"7a00", 110=>x"7900", 111=>x"7a00", 112=>x"7600",
---- 113=>x"7800", 114=>x"7800", 115=>x"7700", 116=>x"7400",
---- 117=>x"7500", 118=>x"7600", 119=>x"7900", 120=>x"7500",
---- 121=>x"7500", 122=>x"7500", 123=>x"7500", 124=>x"7500",
---- 125=>x"7500", 126=>x"7500", 127=>x"7500", 128=>x"7300",
---- 129=>x"7500", 130=>x"7500", 131=>x"7200", 132=>x"7000",
---- 133=>x"7400", 134=>x"7500", 135=>x"7200", 136=>x"7000",
---- 137=>x"7100", 138=>x"7000", 139=>x"8e00", 140=>x"7200",
---- 141=>x"7600", 142=>x"6f00", 143=>x"7100", 144=>x"7100",
---- 145=>x"7200", 146=>x"7200", 147=>x"7400", 148=>x"7100",
---- 149=>x"6f00", 150=>x"7300", 151=>x"8b00", 152=>x"6d00",
---- 153=>x"7100", 154=>x"7200", 155=>x"7600", 156=>x"7200",
---- 157=>x"7500", 158=>x"7400", 159=>x"7300", 160=>x"7000",
---- 161=>x"7200", 162=>x"7700", 163=>x"7100", 164=>x"6e00",
---- 165=>x"7000", 166=>x"7200", 167=>x"7200", 168=>x"7100",
---- 169=>x"7500", 170=>x"7100", 171=>x"7300", 172=>x"7000",
---- 173=>x"7200", 174=>x"7200", 175=>x"7200", 176=>x"6d00",
---- 177=>x"7200", 178=>x"7300", 179=>x"7400", 180=>x"6f00",
---- 181=>x"7200", 182=>x"7400", 183=>x"7300", 184=>x"7000",
---- 185=>x"7000", 186=>x"7400", 187=>x"7600", 188=>x"7400",
---- 189=>x"7200", 190=>x"7300", 191=>x"7400", 192=>x"7000",
---- 193=>x"7000", 194=>x"7700", 195=>x"7800", 196=>x"7000",
---- 197=>x"7300", 198=>x"7900", 199=>x"7500", 200=>x"6d00",
---- 201=>x"7100", 202=>x"7400", 203=>x"7200", 204=>x"7000",
---- 205=>x"7400", 206=>x"7400", 207=>x"7600", 208=>x"6e00",
---- 209=>x"7100", 210=>x"7400", 211=>x"7500", 212=>x"7100",
---- 213=>x"7000", 214=>x"7100", 215=>x"7500", 216=>x"7300",
---- 217=>x"7300", 218=>x"7600", 219=>x"7300", 220=>x"7100",
---- 221=>x"7200", 222=>x"7000", 223=>x"7300", 224=>x"6d00",
---- 225=>x"7200", 226=>x"7300", 227=>x"7200", 228=>x"6e00",
---- 229=>x"7000", 230=>x"7200", 231=>x"8d00", 232=>x"6d00",
---- 233=>x"7100", 234=>x"6f00", 235=>x"6f00", 236=>x"6a00",
---- 237=>x"6d00", 238=>x"6e00", 239=>x"6e00", 240=>x"6c00",
---- 241=>x"6f00", 242=>x"7000", 243=>x"6c00", 244=>x"6d00",
---- 245=>x"7200", 246=>x"7000", 247=>x"6e00", 248=>x"6c00",
---- 249=>x"7100", 250=>x"7200", 251=>x"7500", 252=>x"7000",
---- 253=>x"7000", 254=>x"7300", 255=>x"7300", 256=>x"6e00",
---- 257=>x"7000", 258=>x"7100", 259=>x"6c00", 260=>x"6f00",
---- 261=>x"7100", 262=>x"6f00", 263=>x"6d00", 264=>x"7100",
---- 265=>x"7200", 266=>x"7300", 267=>x"6c00", 268=>x"7000",
---- 269=>x"7200", 270=>x"7200", 271=>x"6d00", 272=>x"6f00",
---- 273=>x"7000", 274=>x"6e00", 275=>x"6800", 276=>x"7000",
---- 277=>x"6d00", 278=>x"6900", 279=>x"6300", 280=>x"6900",
---- 281=>x"6c00", 282=>x"6c00", 283=>x"5e00", 284=>x"6a00",
---- 285=>x"6900", 286=>x"6700", 287=>x"5800", 288=>x"6900",
---- 289=>x"6800", 290=>x"6200", 291=>x"5400", 292=>x"6900",
---- 293=>x"6600", 294=>x"6000", 295=>x"5300", 296=>x"6700",
---- 297=>x"6500", 298=>x"5e00", 299=>x"5b00", 300=>x"6500",
---- 301=>x"6700", 302=>x"5b00", 303=>x"5e00", 304=>x"6700",
---- 305=>x"6600", 306=>x"5b00", 307=>x"6200", 308=>x"6600",
---- 309=>x"6500", 310=>x"5b00", 311=>x"6700", 312=>x"6600",
---- 313=>x"6400", 314=>x"5a00", 315=>x"6300", 316=>x"6500",
---- 317=>x"6500", 318=>x"5900", 319=>x"6600", 320=>x"6100",
---- 321=>x"6200", 322=>x"5500", 323=>x"6b00", 324=>x"6100",
---- 325=>x"5e00", 326=>x"5200", 327=>x"7300", 328=>x"6000",
---- 329=>x"5c00", 330=>x"5000", 331=>x"8100", 332=>x"5e00",
---- 333=>x"5c00", 334=>x"4b00", 335=>x"8c00", 336=>x"5d00",
---- 337=>x"5a00", 338=>x"4b00", 339=>x"9d00", 340=>x"5d00",
---- 341=>x"5600", 342=>x"4900", 343=>x"9800", 344=>x"5c00",
---- 345=>x"5500", 346=>x"4800", 347=>x"9b00", 348=>x"5f00",
---- 349=>x"5700", 350=>x"4600", 351=>x"9500", 352=>x"5b00",
---- 353=>x"5500", 354=>x"4700", 355=>x"9000", 356=>x"5900",
---- 357=>x"5800", 358=>x"4800", 359=>x"8c00", 360=>x"5f00",
---- 361=>x"5b00", 362=>x"4900", 363=>x"7b00", 364=>x"6000",
---- 365=>x"5b00", 366=>x"5000", 367=>x"6600", 368=>x"5f00",
---- 369=>x"5b00", 370=>x"5000", 371=>x"5200", 372=>x"5c00",
---- 373=>x"5a00", 374=>x"5200", 375=>x"4b00", 376=>x"5f00",
---- 377=>x"5f00", 378=>x"5900", 379=>x"4900", 380=>x"6300",
---- 381=>x"5f00", 382=>x"5c00", 383=>x"4900", 384=>x"6400",
---- 385=>x"6000", 386=>x"5b00", 387=>x"5100", 388=>x"6500",
---- 389=>x"6400", 390=>x"5e00", 391=>x"5600", 392=>x"6400",
---- 393=>x"6500", 394=>x"6000", 395=>x"5700", 396=>x"6500",
---- 397=>x"6400", 398=>x"6200", 399=>x"5d00", 400=>x"9300",
---- 401=>x"6700", 402=>x"6500", 403=>x"6100", 404=>x"6700",
---- 405=>x"6a00", 406=>x"9800", 407=>x"6500", 408=>x"6800",
---- 409=>x"6b00", 410=>x"6700", 411=>x"6500", 412=>x"6b00",
---- 413=>x"6800", 414=>x"6a00", 415=>x"6900", 416=>x"6c00",
---- 417=>x"6a00", 418=>x"6c00", 419=>x"6d00", 420=>x"6c00",
---- 421=>x"6f00", 422=>x"7000", 423=>x"6c00", 424=>x"6b00",
---- 425=>x"6d00", 426=>x"7200", 427=>x"7100", 428=>x"6b00",
---- 429=>x"7200", 430=>x"7100", 431=>x"6e00", 432=>x"6c00",
---- 433=>x"7000", 434=>x"7100", 435=>x"7000", 436=>x"6f00",
---- 437=>x"7200", 438=>x"7400", 439=>x"7300", 440=>x"6f00",
---- 441=>x"7100", 442=>x"7100", 443=>x"7100", 444=>x"6b00",
---- 445=>x"6b00", 446=>x"7200", 447=>x"7500", 448=>x"7600",
---- 449=>x"7b00", 450=>x"6e00", 451=>x"7600", 452=>x"a500",
---- 453=>x"7a00", 454=>x"6d00", 455=>x"7500", 456=>x"8200",
---- 457=>x"6d00", 458=>x"7400", 459=>x"7300", 460=>x"6c00",
---- 461=>x"7300", 462=>x"7300", 463=>x"7400", 464=>x"7300",
---- 465=>x"7100", 466=>x"7100", 467=>x"7900", 468=>x"7500",
---- 469=>x"7300", 470=>x"7300", 471=>x"7900", 472=>x"7400",
---- 473=>x"7300", 474=>x"7300", 475=>x"7400", 476=>x"8a00",
---- 477=>x"7600", 478=>x"7200", 479=>x"7000", 480=>x"8c00",
---- 481=>x"7600", 482=>x"7800", 483=>x"7800", 484=>x"8e00",
---- 485=>x"7300", 486=>x"7300", 487=>x"7700", 488=>x"7100",
---- 489=>x"7600", 490=>x"7500", 491=>x"7700", 492=>x"7500",
---- 493=>x"7700", 494=>x"7600", 495=>x"7700", 496=>x"7700",
---- 497=>x"7500", 498=>x"7700", 499=>x"8600", 500=>x"7200",
---- 501=>x"7200", 502=>x"7600", 503=>x"7400", 504=>x"6d00",
---- 505=>x"7400", 506=>x"7200", 507=>x"7900", 508=>x"6b00",
---- 509=>x"9300", 510=>x"7000", 511=>x"8c00", 512=>x"6f00",
---- 513=>x"7900", 514=>x"8700", 515=>x"8e00", 516=>x"6f00",
---- 517=>x"9f00", 518=>x"9200", 519=>x"9100", 520=>x"c300",
---- 521=>x"b200", 522=>x"8100", 523=>x"9500", 524=>x"d400",
---- 525=>x"9200", 526=>x"8200", 527=>x"9100", 528=>x"b300",
---- 529=>x"7800", 530=>x"8800", 531=>x"9100", 532=>x"b900",
---- 533=>x"9800", 534=>x"8a00", 535=>x"9200", 536=>x"7500",
---- 537=>x"b600", 538=>x"b700", 539=>x"9b00", 540=>x"7900",
---- 541=>x"b000", 542=>x"cf00", 543=>x"cf00", 544=>x"a900",
---- 545=>x"be00", 546=>x"e100", 547=>x"f900", 548=>x"a000",
---- 549=>x"d200", 550=>x"d700", 551=>x"8800", 552=>x"b700",
---- 553=>x"ae00", 554=>x"4e00", 555=>x"2a00", 556=>x"9300",
---- 557=>x"4b00", 558=>x"3a00", 559=>x"4300", 560=>x"5600",
---- 561=>x"5000", 562=>x"3e00", 563=>x"3000", 564=>x"6000",
---- 565=>x"4d00", 566=>x"2c00", 567=>x"2700", 568=>x"5300",
---- 569=>x"3c00", 570=>x"2b00", 571=>x"2600", 572=>x"3300",
---- 573=>x"3700", 574=>x"2c00", 575=>x"2f00", 576=>x"3600",
---- 577=>x"c900", 578=>x"cd00", 579=>x"3900", 580=>x"3b00",
---- 581=>x"4500", 582=>x"4000", 583=>x"4400", 584=>x"3e00",
---- 585=>x"4200", 586=>x"3c00", 587=>x"5100", 588=>x"3f00",
---- 589=>x"3900", 590=>x"4b00", 591=>x"5c00", 592=>x"3c00",
---- 593=>x"5000", 594=>x"6f00", 595=>x"4900", 596=>x"5700",
---- 597=>x"7500", 598=>x"5a00", 599=>x"3300", 600=>x"7400",
---- 601=>x"5500", 602=>x"3000", 603=>x"3400", 604=>x"4e00",
---- 605=>x"3200", 606=>x"3d00", 607=>x"3d00", 608=>x"2d00",
---- 609=>x"4c00", 610=>x"5100", 611=>x"4800", 612=>x"2e00",
---- 613=>x"6800", 614=>x"5700", 615=>x"4900", 616=>x"4500",
---- 617=>x"6600", 618=>x"6300", 619=>x"6200", 620=>x"6400",
---- 621=>x"5100", 622=>x"7500", 623=>x"5200", 624=>x"5100",
---- 625=>x"6500", 626=>x"7900", 627=>x"4d00", 628=>x"3f00",
---- 629=>x"7900", 630=>x"5800", 631=>x"3f00", 632=>x"5400",
---- 633=>x"8400", 634=>x"3700", 635=>x"3400", 636=>x"6f00",
---- 637=>x"6e00", 638=>x"2e00", 639=>x"3500", 640=>x"7e00",
---- 641=>x"5300", 642=>x"3300", 643=>x"2c00", 644=>x"7a00",
---- 645=>x"4800", 646=>x"4300", 647=>x"2b00", 648=>x"5100",
---- 649=>x"3d00", 650=>x"5c00", 651=>x"3500", 652=>x"4100",
---- 653=>x"4a00", 654=>x"6b00", 655=>x"3500", 656=>x"4f00",
---- 657=>x"5400", 658=>x"5500", 659=>x"3d00", 660=>x"5000",
---- 661=>x"5300", 662=>x"4500", 663=>x"5900", 664=>x"4b00",
---- 665=>x"4d00", 666=>x"4400", 667=>x"6300", 668=>x"4400",
---- 669=>x"4d00", 670=>x"4400", 671=>x"4d00", 672=>x"4100",
---- 673=>x"4600", 674=>x"4800", 675=>x"4300", 676=>x"4400",
---- 677=>x"4300", 678=>x"4d00", 679=>x"3e00", 680=>x"4700",
---- 681=>x"3800", 682=>x"5200", 683=>x"4600", 684=>x"4600",
---- 685=>x"3b00", 686=>x"4a00", 687=>x"5400", 688=>x"3f00",
---- 689=>x"5400", 690=>x"5300", 691=>x"5300", 692=>x"4300",
---- 693=>x"4d00", 694=>x"6a00", 695=>x"5600", 696=>x"3900",
---- 697=>x"4600", 698=>x"7800", 699=>x"5f00", 700=>x"3300",
---- 701=>x"4e00", 702=>x"8800", 703=>x"7700", 704=>x"3500",
---- 705=>x"4d00", 706=>x"8800", 707=>x"7f00", 708=>x"3400",
---- 709=>x"4a00", 710=>x"6300", 711=>x"8600", 712=>x"3700",
---- 713=>x"4b00", 714=>x"aa00", 715=>x"8400", 716=>x"4500",
---- 717=>x"5000", 718=>x"ac00", 719=>x"8500", 720=>x"5400",
---- 721=>x"6b00", 722=>x"a700", 723=>x"7900", 724=>x"4e00",
---- 725=>x"8800", 726=>x"6800", 727=>x"5e00", 728=>x"5200",
---- 729=>x"9b00", 730=>x"9900", 731=>x"5500", 732=>x"6200",
---- 733=>x"ad00", 734=>x"9a00", 735=>x"6700", 736=>x"7000",
---- 737=>x"ad00", 738=>x"8500", 739=>x"8d00", 740=>x"6d00",
---- 741=>x"ab00", 742=>x"8200", 743=>x"7100", 744=>x"5200",
---- 745=>x"9700", 746=>x"6c00", 747=>x"6500", 748=>x"5300",
---- 749=>x"8f00", 750=>x"6000", 751=>x"5e00", 752=>x"5b00",
---- 753=>x"7e00", 754=>x"6700", 755=>x"4e00", 756=>x"6600",
---- 757=>x"8300", 758=>x"6300", 759=>x"4900", 760=>x"6600",
---- 761=>x"8a00", 762=>x"7e00", 763=>x"5c00", 764=>x"5300",
---- 765=>x"9200", 766=>x"8100", 767=>x"7100", 768=>x"4000",
---- 769=>x"9900", 770=>x"8400", 771=>x"7d00", 772=>x"3700",
---- 773=>x"9000", 774=>x"9000", 775=>x"9000", 776=>x"3400",
---- 777=>x"8500", 778=>x"8300", 779=>x"9200", 780=>x"4000",
---- 781=>x"8500", 782=>x"7800", 783=>x"7b00", 784=>x"4200",
---- 785=>x"7e00", 786=>x"8200", 787=>x"6f00", 788=>x"3800",
---- 789=>x"5600", 790=>x"7b00", 791=>x"8300", 792=>x"3a00",
---- 793=>x"3500", 794=>x"4a00", 795=>x"8700", 796=>x"4a00",
---- 797=>x"3200", 798=>x"2100", 799=>x"6b00", 800=>x"5d00",
---- 801=>x"2d00", 802=>x"1f00", 803=>x"3800", 804=>x"6a00",
---- 805=>x"2e00", 806=>x"2900", 807=>x"2500", 808=>x"4900",
---- 809=>x"3300", 810=>x"2c00", 811=>x"2e00", 812=>x"4c00",
---- 813=>x"3200", 814=>x"2a00", 815=>x"6000", 816=>x"4800",
---- 817=>x"4300", 818=>x"6700", 819=>x"8000", 820=>x"a500",
---- 821=>x"6700", 822=>x"6600", 823=>x"4c00", 824=>x"3a00",
---- 825=>x"3100", 826=>x"2f00", 827=>x"3500", 828=>x"2d00",
---- 829=>x"2800", 830=>x"2a00", 831=>x"4000", 832=>x"3500",
---- 833=>x"2800", 834=>x"2800", 835=>x"4500", 836=>x"4800",
---- 837=>x"2900", 838=>x"2700", 839=>x"3700", 840=>x"4900",
---- 841=>x"2a00", 842=>x"2500", 843=>x"2700", 844=>x"4600",
---- 845=>x"3200", 846=>x"2600", 847=>x"2300", 848=>x"5200",
---- 849=>x"3a00", 850=>x"2400", 851=>x"2600", 852=>x"5200",
---- 853=>x"3800", 854=>x"2400", 855=>x"2700", 856=>x"4b00",
---- 857=>x"4700", 858=>x"2600", 859=>x"2e00", 860=>x"3e00",
---- 861=>x"4d00", 862=>x"2800", 863=>x"3500", 864=>x"3000",
---- 865=>x"3f00", 866=>x"2900", 867=>x"3e00", 868=>x"2b00",
---- 869=>x"3700", 870=>x"3000", 871=>x"4100", 872=>x"2900",
---- 873=>x"2e00", 874=>x"3a00", 875=>x"4500", 876=>x"2e00",
---- 877=>x"3200", 878=>x"4500", 879=>x"4a00", 880=>x"2d00",
---- 881=>x"3300", 882=>x"4f00", 883=>x"4300", 884=>x"2800",
---- 885=>x"3600", 886=>x"4600", 887=>x"3a00", 888=>x"3400",
---- 889=>x"3e00", 890=>x"2f00", 891=>x"3700", 892=>x"3c00",
---- 893=>x"3d00", 894=>x"2c00", 895=>x"3500", 896=>x"3a00",
---- 897=>x"3000", 898=>x"2f00", 899=>x"3c00", 900=>x"2b00",
---- 901=>x"2d00", 902=>x"2e00", 903=>x"3500", 904=>x"3000",
---- 905=>x"3200", 906=>x"3300", 907=>x"2f00", 908=>x"c600",
---- 909=>x"3800", 910=>x"3800", 911=>x"2f00", 912=>x"3f00",
---- 913=>x"4500", 914=>x"4100", 915=>x"3300", 916=>x"3f00",
---- 917=>x"3a00", 918=>x"3d00", 919=>x"3b00", 920=>x"4500",
---- 921=>x"3000", 922=>x"3100", 923=>x"3200", 924=>x"4900",
---- 925=>x"2f00", 926=>x"2a00", 927=>x"2b00", 928=>x"4900",
---- 929=>x"3500", 930=>x"3000", 931=>x"2c00", 932=>x"4300",
---- 933=>x"3700", 934=>x"3400", 935=>x"2f00", 936=>x"4200",
---- 937=>x"3900", 938=>x"3d00", 939=>x"3900", 940=>x"4300",
---- 941=>x"4000", 942=>x"4100", 943=>x"3a00", 944=>x"3b00",
---- 945=>x"3b00", 946=>x"3900", 947=>x"3600", 948=>x"3b00",
---- 949=>x"3a00", 950=>x"3a00", 951=>x"3800", 952=>x"4200",
---- 953=>x"3600", 954=>x"3f00", 955=>x"3d00", 956=>x"4700",
---- 957=>x"3c00", 958=>x"4000", 959=>x"3e00", 960=>x"4800",
---- 961=>x"3b00", 962=>x"3a00", 963=>x"3a00", 964=>x"4200",
---- 965=>x"3500", 966=>x"3000", 967=>x"3f00", 968=>x"4500",
---- 969=>x"3100", 970=>x"3000", 971=>x"4b00", 972=>x"5400",
---- 973=>x"3000", 974=>x"3800", 975=>x"4b00", 976=>x"6300",
---- 977=>x"2f00", 978=>x"c900", 979=>x"5100", 980=>x"6200",
---- 981=>x"2900", 982=>x"3500", 983=>x"5000", 984=>x"5600",
---- 985=>x"2800", 986=>x"3500", 987=>x"5600", 988=>x"4c00",
---- 989=>x"2700", 990=>x"2e00", 991=>x"5100", 992=>x"3a00",
---- 993=>x"2a00", 994=>x"2900", 995=>x"4800", 996=>x"2a00",
---- 997=>x"2c00", 998=>x"2700", 999=>x"4400", 1000=>x"2f00",
---- 1001=>x"2c00", 1002=>x"2b00", 1003=>x"4200", 1004=>x"2d00",
---- 1005=>x"3000", 1006=>x"2f00", 1007=>x"4700", 1008=>x"3100",
---- 1009=>x"2f00", 1010=>x"2c00", 1011=>x"5000", 1012=>x"3a00",
---- 1013=>x"2e00", 1014=>x"3700", 1015=>x"5300", 1016=>x"3d00",
---- 1017=>x"3400", 1018=>x"3c00", 1019=>x"4f00", 1020=>x"4500",
---- 1021=>x"3200", 1022=>x"3600", 1023=>x"4e00"),
----
---- 15 => (0=>x"7d00", 1=>x"8000", 2=>x"7a00", 3=>x"8300", 4=>x"7f00",
---- 5=>x"8000", 6=>x"7b00", 7=>x"8300", 8=>x"7e00",
---- 9=>x"8000", 10=>x"7b00", 11=>x"8100", 12=>x"7d00",
---- 13=>x"7b00", 14=>x"7c00", 15=>x"7c00", 16=>x"7d00",
---- 17=>x"7d00", 18=>x"7b00", 19=>x"7c00", 20=>x"7b00",
---- 21=>x"7c00", 22=>x"7d00", 23=>x"8000", 24=>x"7a00",
---- 25=>x"7d00", 26=>x"7f00", 27=>x"7d00", 28=>x"7d00",
---- 29=>x"7c00", 30=>x"7d00", 31=>x"8000", 32=>x"7c00",
---- 33=>x"7e00", 34=>x"7f00", 35=>x"8000", 36=>x"7b00",
---- 37=>x"7d00", 38=>x"7a00", 39=>x"7f00", 40=>x"7c00",
---- 41=>x"7c00", 42=>x"7a00", 43=>x"7d00", 44=>x"7b00",
---- 45=>x"7d00", 46=>x"7d00", 47=>x"7b00", 48=>x"7800",
---- 49=>x"7800", 50=>x"7f00", 51=>x"7f00", 52=>x"7a00",
---- 53=>x"7c00", 54=>x"7b00", 55=>x"7d00", 56=>x"7c00",
---- 57=>x"7d00", 58=>x"7c00", 59=>x"7f00", 60=>x"7a00",
---- 61=>x"7c00", 62=>x"7d00", 63=>x"7b00", 64=>x"7c00",
---- 65=>x"7800", 66=>x"7a00", 67=>x"8200", 68=>x"7c00",
---- 69=>x"7c00", 70=>x"7b00", 71=>x"7e00", 72=>x"7600",
---- 73=>x"7800", 74=>x"7d00", 75=>x"7b00", 76=>x"7600",
---- 77=>x"7700", 78=>x"7a00", 79=>x"7c00", 80=>x"7900",
---- 81=>x"7a00", 82=>x"7700", 83=>x"7800", 84=>x"7600",
---- 85=>x"8500", 86=>x"8300", 87=>x"7a00", 88=>x"7700",
---- 89=>x"7a00", 90=>x"7d00", 91=>x"7b00", 92=>x"7a00",
---- 93=>x"7c00", 94=>x"7a00", 95=>x"7b00", 96=>x"8700",
---- 97=>x"7c00", 98=>x"7c00", 99=>x"7c00", 100=>x"7800",
---- 101=>x"8500", 102=>x"7e00", 103=>x"7c00", 104=>x"7800",
---- 105=>x"7800", 106=>x"7a00", 107=>x"7c00", 108=>x"7c00",
---- 109=>x"7a00", 110=>x"7b00", 111=>x"7e00", 112=>x"7a00",
---- 113=>x"7a00", 114=>x"7e00", 115=>x"7b00", 116=>x"7a00",
---- 117=>x"7900", 118=>x"7b00", 119=>x"7a00", 120=>x"7800",
---- 121=>x"7b00", 122=>x"7900", 123=>x"7900", 124=>x"7700",
---- 125=>x"7a00", 126=>x"7900", 127=>x"7700", 128=>x"7800",
---- 129=>x"7700", 130=>x"7900", 131=>x"7600", 132=>x"7700",
---- 133=>x"7400", 134=>x"7300", 135=>x"7500", 136=>x"7200",
---- 137=>x"8900", 138=>x"7500", 139=>x"7600", 140=>x"7400",
---- 141=>x"7500", 142=>x"7600", 143=>x"7700", 144=>x"7300",
---- 145=>x"7500", 146=>x"7300", 147=>x"7600", 148=>x"7100",
---- 149=>x"7200", 150=>x"7400", 151=>x"7600", 152=>x"8d00",
---- 153=>x"7300", 154=>x"7500", 155=>x"7a00", 156=>x"7200",
---- 157=>x"7100", 158=>x"7200", 159=>x"7400", 160=>x"7400",
---- 161=>x"7400", 162=>x"7800", 163=>x"7700", 164=>x"7100",
---- 165=>x"7400", 166=>x"7500", 167=>x"7900", 168=>x"7500",
---- 169=>x"7500", 170=>x"7600", 171=>x"7600", 172=>x"7400",
---- 173=>x"7500", 174=>x"7500", 175=>x"7600", 176=>x"7500",
---- 177=>x"7300", 178=>x"7600", 179=>x"7800", 180=>x"7400",
---- 181=>x"7500", 182=>x"7800", 183=>x"7b00", 184=>x"7400",
---- 185=>x"7600", 186=>x"7800", 187=>x"7800", 188=>x"7400",
---- 189=>x"7600", 190=>x"7700", 191=>x"7600", 192=>x"7300",
---- 193=>x"7400", 194=>x"7500", 195=>x"7500", 196=>x"7400",
---- 197=>x"7200", 198=>x"7600", 199=>x"7800", 200=>x"7200",
---- 201=>x"7700", 202=>x"7700", 203=>x"7500", 204=>x"7600",
---- 205=>x"7600", 206=>x"7600", 207=>x"7600", 208=>x"7700",
---- 209=>x"7a00", 210=>x"7800", 211=>x"7300", 212=>x"7600",
---- 213=>x"7400", 214=>x"7500", 215=>x"7200", 216=>x"7000",
---- 217=>x"7300", 218=>x"7200", 219=>x"7100", 220=>x"7500",
---- 221=>x"7400", 222=>x"6e00", 223=>x"6b00", 224=>x"6f00",
---- 225=>x"6e00", 226=>x"6d00", 227=>x"6700", 228=>x"6f00",
---- 229=>x"6f00", 230=>x"6b00", 231=>x"6b00", 232=>x"6c00",
---- 233=>x"6b00", 234=>x"6100", 235=>x"8300", 236=>x"6b00",
---- 237=>x"6500", 238=>x"6100", 239=>x"a700", 240=>x"6e00",
---- 241=>x"6500", 242=>x"6f00", 243=>x"c700", 244=>x"6c00",
---- 245=>x"6200", 246=>x"8000", 247=>x"d100", 248=>x"6d00",
---- 249=>x"5f00", 250=>x"9e00", 251=>x"dc00", 252=>x"6e00",
---- 253=>x"6500", 254=>x"b000", 255=>x"d600", 256=>x"6400",
---- 257=>x"6900", 258=>x"c400", 259=>x"d100", 260=>x"6400",
---- 261=>x"7300", 262=>x"cf00", 263=>x"cf00", 264=>x"5f00",
---- 265=>x"8700", 266=>x"d800", 267=>x"cc00", 268=>x"6000",
---- 269=>x"9a00", 270=>x"2400", 271=>x"ca00", 272=>x"5b00",
---- 273=>x"ab00", 274=>x"df00", 275=>x"bf00", 276=>x"5d00",
---- 277=>x"b700", 278=>x"db00", 279=>x"ac00", 280=>x"6a00",
---- 281=>x"cb00", 282=>x"d400", 283=>x"a400", 284=>x"7900",
---- 285=>x"d800", 286=>x"cb00", 287=>x"ad00", 288=>x"8d00",
---- 289=>x"de00", 290=>x"c900", 291=>x"aa00", 292=>x"a500",
---- 293=>x"de00", 294=>x"c300", 295=>x"af00", 296=>x"bb00",
---- 297=>x"dd00", 298=>x"c200", 299=>x"b000", 300=>x"c000",
---- 301=>x"db00", 302=>x"bb00", 303=>x"b700", 304=>x"c800",
---- 305=>x"d500", 306=>x"be00", 307=>x"af00", 308=>x"2f00",
---- 309=>x"d500", 310=>x"bb00", 311=>x"b200", 312=>x"cc00",
---- 313=>x"d000", 314=>x"b900", 315=>x"ad00", 316=>x"d200",
---- 317=>x"cc00", 318=>x"ba00", 319=>x"b100", 320=>x"d100",
---- 321=>x"c300", 322=>x"bb00", 323=>x"ad00", 324=>x"d700",
---- 325=>x"c500", 326=>x"b200", 327=>x"b100", 328=>x"db00",
---- 329=>x"ba00", 330=>x"b900", 331=>x"ad00", 332=>x"d500",
---- 333=>x"c300", 334=>x"b600", 335=>x"bd00", 336=>x"db00",
---- 337=>x"c100", 338=>x"c500", 339=>x"b400", 340=>x"da00",
---- 341=>x"cc00", 342=>x"be00", 343=>x"c100", 344=>x"e000",
---- 345=>x"c500", 346=>x"c800", 347=>x"bd00", 348=>x"dc00",
---- 349=>x"3100", 350=>x"c400", 351=>x"c400", 352=>x"1d00",
---- 353=>x"c700", 354=>x"c400", 355=>x"c700", 356=>x"db00",
---- 357=>x"ce00", 358=>x"c800", 359=>x"c000", 360=>x"dd00",
---- 361=>x"ce00", 362=>x"c400", 363=>x"c800", 364=>x"ce00",
---- 365=>x"2e00", 366=>x"c900", 367=>x"c100", 368=>x"bb00",
---- 369=>x"d900", 370=>x"c600", 371=>x"ce00", 372=>x"ab00",
---- 373=>x"da00", 374=>x"cf00", 375=>x"c700", 376=>x"8a00",
---- 377=>x"e000", 378=>x"c200", 379=>x"d000", 380=>x"6c00",
---- 381=>x"d200", 382=>x"d200", 383=>x"c500", 384=>x"4f00",
---- 385=>x"ba00", 386=>x"d900", 387=>x"ca00", 388=>x"4900",
---- 389=>x"8d00", 390=>x"dd00", 391=>x"c500", 392=>x"4a00",
---- 393=>x"7300", 394=>x"da00", 395=>x"ce00", 396=>x"5200",
---- 397=>x"5c00", 398=>x"c300", 399=>x"d300", 400=>x"5b00",
---- 401=>x"5100", 402=>x"8100", 403=>x"dd00", 404=>x"6000",
---- 405=>x"5500", 406=>x"5a00", 407=>x"bb00", 408=>x"6400",
---- 409=>x"5f00", 410=>x"5100", 411=>x"7500", 412=>x"6600",
---- 413=>x"5f00", 414=>x"5b00", 415=>x"5000", 416=>x"6a00",
---- 417=>x"6600", 418=>x"5f00", 419=>x"5100", 420=>x"6b00",
---- 421=>x"6900", 422=>x"6200", 423=>x"5c00", 424=>x"6c00",
---- 425=>x"6900", 426=>x"6500", 427=>x"5f00", 428=>x"6d00",
---- 429=>x"9200", 430=>x"6900", 431=>x"5f00", 432=>x"6e00",
---- 433=>x"6b00", 434=>x"6800", 435=>x"6200", 436=>x"6f00",
---- 437=>x"6d00", 438=>x"6a00", 439=>x"6500", 440=>x"7100",
---- 441=>x"6f00", 442=>x"6d00", 443=>x"6600", 444=>x"7100",
---- 445=>x"6d00", 446=>x"7000", 447=>x"6800", 448=>x"7100",
---- 449=>x"7200", 450=>x"7000", 451=>x"6d00", 452=>x"7100",
---- 453=>x"7100", 454=>x"6f00", 455=>x"6c00", 456=>x"7300",
---- 457=>x"7200", 458=>x"7300", 459=>x"7400", 460=>x"7500",
---- 461=>x"7500", 462=>x"7300", 463=>x"7300", 464=>x"7700",
---- 465=>x"7700", 466=>x"7500", 467=>x"7500", 468=>x"7800",
---- 469=>x"7800", 470=>x"7900", 471=>x"7900", 472=>x"7700",
---- 473=>x"7400", 474=>x"7500", 475=>x"7500", 476=>x"6f00",
---- 477=>x"6e00", 478=>x"6d00", 479=>x"6b00", 480=>x"7500",
---- 481=>x"7900", 482=>x"7600", 483=>x"7600", 484=>x"7700",
---- 485=>x"7900", 486=>x"7800", 487=>x"7600", 488=>x"7800",
---- 489=>x"7700", 490=>x"7500", 491=>x"8300", 492=>x"7700",
---- 493=>x"7900", 494=>x"7200", 495=>x"b500", 496=>x"8300",
---- 497=>x"7a00", 498=>x"7900", 499=>x"b300", 500=>x"7b00",
---- 501=>x"8400", 502=>x"8700", 503=>x"8d00", 504=>x"8e00",
---- 505=>x"9a00", 506=>x"9100", 507=>x"8700", 508=>x"9b00",
---- 509=>x"9d00", 510=>x"9600", 511=>x"9000", 512=>x"9800",
---- 513=>x"9d00", 514=>x"9a00", 515=>x"9700", 516=>x"9700",
---- 517=>x"9b00", 518=>x"9a00", 519=>x"9800", 520=>x"9300",
---- 521=>x"6800", 522=>x"9900", 523=>x"9b00", 524=>x"9300",
---- 525=>x"9800", 526=>x"9e00", 527=>x"9000", 528=>x"9600",
---- 529=>x"9b00", 530=>x"9800", 531=>x"6900", 532=>x"9500",
---- 533=>x"9700", 534=>x"9200", 535=>x"7200", 536=>x"9400",
---- 537=>x"9a00", 538=>x"8600", 539=>x"6100", 540=>x"c000",
---- 541=>x"9400", 542=>x"4300", 543=>x"2700", 544=>x"bf00",
---- 545=>x"4f00", 546=>x"3f00", 547=>x"2a00", 548=>x"3d00",
---- 549=>x"2d00", 550=>x"5c00", 551=>x"3400", 552=>x"2e00",
---- 553=>x"2a00", 554=>x"5200", 555=>x"6400", 556=>x"3500",
---- 557=>x"3200", 558=>x"3a00", 559=>x"7300", 560=>x"2800",
---- 561=>x"3000", 562=>x"2500", 563=>x"4200", 564=>x"3000",
---- 565=>x"3400", 566=>x"2c00", 567=>x"3300", 568=>x"4400",
---- 569=>x"4000", 570=>x"3800", 571=>x"4400", 572=>x"af00",
---- 573=>x"4700", 574=>x"4f00", 575=>x"6c00", 576=>x"6400",
---- 577=>x"5100", 578=>x"6700", 579=>x"7600", 580=>x"6c00",
---- 581=>x"4c00", 582=>x"6900", 583=>x"7600", 584=>x"6500",
---- 585=>x"4c00", 586=>x"6e00", 587=>x"5a00", 588=>x"4f00",
---- 589=>x"6100", 590=>x"7000", 591=>x"7100", 592=>x"4200",
---- 593=>x"7200", 594=>x"8200", 595=>x"8700", 596=>x"4b00",
---- 597=>x"8800", 598=>x"7900", 599=>x"6500", 600=>x"4700",
---- 601=>x"7500", 602=>x"7f00", 603=>x"6000", 604=>x"3000",
---- 605=>x"4a00", 606=>x"8700", 607=>x"6200", 608=>x"3800",
---- 609=>x"4d00", 610=>x"8800", 611=>x"6d00", 612=>x"3900",
---- 613=>x"8100", 614=>x"7300", 615=>x"7700", 616=>x"4b00",
---- 617=>x"8b00", 618=>x"7000", 619=>x"7e00", 620=>x"5a00",
---- 621=>x"8000", 622=>x"6800", 623=>x"8f00", 624=>x"5f00",
---- 625=>x"6a00", 626=>x"6800", 627=>x"9b00", 628=>x"6000",
---- 629=>x"5900", 630=>x"6200", 631=>x"9c00", 632=>x"7200",
---- 633=>x"5900", 634=>x"5a00", 635=>x"9800", 636=>x"8500",
---- 637=>x"6500", 638=>x"4b00", 639=>x"9500", 640=>x"6a00",
---- 641=>x"6c00", 642=>x"3f00", 643=>x"8100", 644=>x"5a00",
---- 645=>x"8c00", 646=>x"5100", 647=>x"7300", 648=>x"5500",
---- 649=>x"6d00", 650=>x"5900", 651=>x"6f00", 652=>x"4d00",
---- 653=>x"7900", 654=>x"5c00", 655=>x"6c00", 656=>x"4900",
---- 657=>x"7e00", 658=>x"5300", 659=>x"6300", 660=>x"5100",
---- 661=>x"7200", 662=>x"5500", 663=>x"7400", 664=>x"6b00",
---- 665=>x"7000", 666=>x"6800", 667=>x"7900", 668=>x"6700",
---- 669=>x"6100", 670=>x"6700", 671=>x"7a00", 672=>x"5900",
---- 673=>x"4800", 674=>x"5b00", 675=>x"6f00", 676=>x"5100",
---- 677=>x"4800", 678=>x"5900", 679=>x"7000", 680=>x"4500",
---- 681=>x"4a00", 682=>x"4500", 683=>x"7000", 684=>x"4100",
---- 685=>x"4500", 686=>x"4100", 687=>x"5d00", 688=>x"4a00",
---- 689=>x"4000", 690=>x"4a00", 691=>x"b100", 692=>x"6000",
---- 693=>x"5400", 694=>x"4f00", 695=>x"4f00", 696=>x"6400",
---- 697=>x"6600", 698=>x"5700", 699=>x"4b00", 700=>x"6700",
---- 701=>x"6300", 702=>x"6900", 703=>x"5a00", 704=>x"6700",
---- 705=>x"5e00", 706=>x"6600", 707=>x"6500", 708=>x"5500",
---- 709=>x"5b00", 710=>x"6200", 711=>x"5f00", 712=>x"4a00",
---- 713=>x"3d00", 714=>x"5c00", 715=>x"6d00", 716=>x"4f00",
---- 717=>x"3200", 718=>x"5100", 719=>x"5a00", 720=>x"8800",
---- 721=>x"3c00", 722=>x"4800", 723=>x"5800", 724=>x"8100",
---- 725=>x"9a00", 726=>x"4c00", 727=>x"7000", 728=>x"5b00",
---- 729=>x"8600", 730=>x"6600", 731=>x"7d00", 732=>x"3e00",
---- 733=>x"8800", 734=>x"7900", 735=>x"7b00", 736=>x"5400",
---- 737=>x"6700", 738=>x"9000", 739=>x"8000", 740=>x"7b00",
---- 741=>x"5e00", 742=>x"9300", 743=>x"8b00", 744=>x"7500",
---- 745=>x"6d00", 746=>x"7600", 747=>x"9500", 748=>x"6d00",
---- 749=>x"7700", 750=>x"6e00", 751=>x"8400", 752=>x"3e00",
---- 753=>x"5200", 754=>x"7300", 755=>x"7b00", 756=>x"3200",
---- 757=>x"3600", 758=>x"4600", 759=>x"6e00", 760=>x"2f00",
---- 761=>x"4200", 762=>x"4300", 763=>x"a400", 764=>x"3600",
---- 765=>x"4800", 766=>x"5000", 767=>x"5a00", 768=>x"4000",
---- 769=>x"4300", 770=>x"5200", 771=>x"4400", 772=>x"5f00",
---- 773=>x"5600", 774=>x"5f00", 775=>x"3f00", 776=>x"8900",
---- 777=>x"5800", 778=>x"5700", 779=>x"4300", 780=>x"9300",
---- 781=>x"5f00", 782=>x"4c00", 783=>x"4e00", 784=>x"8100",
---- 785=>x"9400", 786=>x"5f00", 787=>x"3f00", 788=>x"6c00",
---- 789=>x"7f00", 790=>x"8b00", 791=>x"5100", 792=>x"7b00",
---- 793=>x"ab00", 794=>x"7e00", 795=>x"8400", 796=>x"8e00",
---- 797=>x"6e00", 798=>x"5500", 799=>x"4500", 800=>x"7400",
---- 801=>x"8b00", 802=>x"7800", 803=>x"5000", 804=>x"4000",
---- 805=>x"7600", 806=>x"8300", 807=>x"8a00", 808=>x"5b00",
---- 809=>x"5300", 810=>x"3c00", 811=>x"6000", 812=>x"6f00",
---- 813=>x"4200", 814=>x"3800", 815=>x"5200", 816=>x"4500",
---- 817=>x"2c00", 818=>x"3a00", 819=>x"7a00", 820=>x"2900",
---- 821=>x"2000", 822=>x"5400", 823=>x"9200", 824=>x"2e00",
---- 825=>x"2b00", 826=>x"9e00", 827=>x"8b00", 828=>x"4000",
---- 829=>x"2900", 830=>x"3900", 831=>x"5700", 832=>x"5b00",
---- 833=>x"2700", 834=>x"2700", 835=>x"3e00", 836=>x"6a00",
---- 837=>x"3800", 838=>x"2700", 839=>x"3800", 840=>x"5f00",
---- 841=>x"5800", 842=>x"2700", 843=>x"2d00", 844=>x"3600",
---- 845=>x"5c00", 846=>x"4b00", 847=>x"2600", 848=>x"2700",
---- 849=>x"3100", 850=>x"6000", 851=>x"5100", 852=>x"3300",
---- 853=>x"2900", 854=>x"3e00", 855=>x"5800", 856=>x"3b00",
---- 857=>x"2b00", 858=>x"3800", 859=>x"3600", 860=>x"4200",
---- 861=>x"2d00", 862=>x"3f00", 863=>x"3a00", 864=>x"4400",
---- 865=>x"3000", 866=>x"3600", 867=>x"3b00", 868=>x"3b00",
---- 869=>x"3600", 870=>x"2e00", 871=>x"3200", 872=>x"2f00",
---- 873=>x"3500", 874=>x"2700", 875=>x"2700", 876=>x"2a00",
---- 877=>x"3500", 878=>x"2d00", 879=>x"2600", 880=>x"2d00",
---- 881=>x"2d00", 882=>x"3000", 883=>x"2700", 884=>x"3500",
---- 885=>x"2900", 886=>x"2e00", 887=>x"2a00", 888=>x"3800",
---- 889=>x"2e00", 890=>x"3300", 891=>x"3100", 892=>x"3d00",
---- 893=>x"3000", 894=>x"3200", 895=>x"2c00", 896=>x"4500",
---- 897=>x"2e00", 898=>x"2a00", 899=>x"2600", 900=>x"4c00",
---- 901=>x"3700", 902=>x"2500", 903=>x"2b00", 904=>x"4100",
---- 905=>x"3d00", 906=>x"2500", 907=>x"2b00", 908=>x"3500",
---- 909=>x"5100", 910=>x"2a00", 911=>x"3200", 912=>x"2900",
---- 913=>x"4200", 914=>x"3c00", 915=>x"3c00", 916=>x"3500",
---- 917=>x"4000", 918=>x"3e00", 919=>x"2e00", 920=>x"3c00",
---- 921=>x"3700", 922=>x"2c00", 923=>x"2700", 924=>x"3100",
---- 925=>x"3400", 926=>x"2f00", 927=>x"2900", 928=>x"2e00",
---- 929=>x"2b00", 930=>x"3100", 931=>x"2800", 932=>x"2b00",
---- 933=>x"2b00", 934=>x"3200", 935=>x"3300", 936=>x"2a00",
---- 937=>x"2b00", 938=>x"3100", 939=>x"3500", 940=>x"3200",
---- 941=>x"2800", 942=>x"3500", 943=>x"3200", 944=>x"3a00",
---- 945=>x"3700", 946=>x"3400", 947=>x"2e00", 948=>x"3400",
---- 949=>x"3c00", 950=>x"2d00", 951=>x"2a00", 952=>x"3100",
---- 953=>x"2f00", 954=>x"2a00", 955=>x"2c00", 956=>x"2d00",
---- 957=>x"2f00", 958=>x"2f00", 959=>x"2a00", 960=>x"3b00",
---- 961=>x"2e00", 962=>x"2c00", 963=>x"2c00", 964=>x"5400",
---- 965=>x"3700", 966=>x"3100", 967=>x"3100", 968=>x"5b00",
---- 969=>x"3900", 970=>x"2a00", 971=>x"3400", 972=>x"5b00",
---- 973=>x"4d00", 974=>x"2a00", 975=>x"2e00", 976=>x"5f00",
---- 977=>x"5800", 978=>x"3d00", 979=>x"2600", 980=>x"6500",
---- 981=>x"6100", 982=>x"5b00", 983=>x"3200", 984=>x"6c00",
---- 985=>x"7300", 986=>x"6b00", 987=>x"4a00", 988=>x"6900",
---- 989=>x"7000", 990=>x"6c00", 991=>x"5200", 992=>x"6500",
---- 993=>x"5d00", 994=>x"7f00", 995=>x"9e00", 996=>x"7000",
---- 997=>x"4700", 998=>x"7000", 999=>x"8000", 1000=>x"7700",
---- 1001=>x"4600", 1002=>x"5100", 1003=>x"8e00", 1004=>x"7900",
---- 1005=>x"5000", 1006=>x"4200", 1007=>x"8800", 1008=>x"7e00",
---- 1009=>x"4c00", 1010=>x"4600", 1011=>x"6700", 1012=>x"7700",
---- 1013=>x"3d00", 1014=>x"4c00", 1015=>x"4a00", 1016=>x"7d00",
---- 1017=>x"3800", 1018=>x"4300", 1019=>x"5300", 1020=>x"7a00",
---- 1021=>x"3b00", 1022=>x"3300", 1023=>x"5300"),
----
---- 16 => (0=>x"7c00", 1=>x"8300", 2=>x"8000", 3=>x"8100", 4=>x"8300",
---- 5=>x"8300", 6=>x"8100", 7=>x"8100", 8=>x"8200",
---- 9=>x"8300", 10=>x"8200", 11=>x"8100", 12=>x"7c00",
---- 13=>x"8100", 14=>x"8400", 15=>x"8000", 16=>x"7e00",
---- 17=>x"8000", 18=>x"8000", 19=>x"8200", 20=>x"7f00",
---- 21=>x"8300", 22=>x"7f00", 23=>x"8000", 24=>x"7e00",
---- 25=>x"7e00", 26=>x"7f00", 27=>x"8300", 28=>x"7e00",
---- 29=>x"7d00", 30=>x"8000", 31=>x"8000", 32=>x"7f00",
---- 33=>x"8100", 34=>x"7f00", 35=>x"8300", 36=>x"8000",
---- 37=>x"8000", 38=>x"8000", 39=>x"8200", 40=>x"7d00",
---- 41=>x"7f00", 42=>x"8000", 43=>x"8100", 44=>x"7c00",
---- 45=>x"8000", 46=>x"8000", 47=>x"8200", 48=>x"8000",
---- 49=>x"8300", 50=>x"7f00", 51=>x"7e00", 52=>x"7f00",
---- 53=>x"8100", 54=>x"8000", 55=>x"7d00", 56=>x"8000",
---- 57=>x"7e00", 58=>x"7d00", 59=>x"7e00", 60=>x"7e00",
---- 61=>x"7e00", 62=>x"8000", 63=>x"7f00", 64=>x"7e00",
---- 65=>x"7e00", 66=>x"8100", 67=>x"7d00", 68=>x"7d00",
---- 69=>x"7d00", 70=>x"7f00", 71=>x"8100", 72=>x"7a00",
---- 73=>x"7c00", 74=>x"7f00", 75=>x"8000", 76=>x"7c00",
---- 77=>x"7d00", 78=>x"7e00", 79=>x"7e00", 80=>x"7c00",
---- 81=>x"7a00", 82=>x"7900", 83=>x"7e00", 84=>x"7c00",
---- 85=>x"7d00", 86=>x"7800", 87=>x"7c00", 88=>x"7d00",
---- 89=>x"7d00", 90=>x"7c00", 91=>x"7b00", 92=>x"7b00",
---- 93=>x"7c00", 94=>x"7b00", 95=>x"7e00", 96=>x"7b00",
---- 97=>x"7d00", 98=>x"7c00", 99=>x"7f00", 100=>x"7f00",
---- 101=>x"7c00", 102=>x"8400", 103=>x"7e00", 104=>x"7f00",
---- 105=>x"8000", 106=>x"7d00", 107=>x"7d00", 108=>x"8200",
---- 109=>x"7e00", 110=>x"7f00", 111=>x"7c00", 112=>x"7f00",
---- 113=>x"7c00", 114=>x"7c00", 115=>x"7d00", 116=>x"7c00",
---- 117=>x"7900", 118=>x"7a00", 119=>x"7b00", 120=>x"7800",
---- 121=>x"7a00", 122=>x"7d00", 123=>x"7a00", 124=>x"7a00",
---- 125=>x"7a00", 126=>x"7d00", 127=>x"7b00", 128=>x"7b00",
---- 129=>x"7900", 130=>x"7b00", 131=>x"7b00", 132=>x"7c00",
---- 133=>x"7c00", 134=>x"7a00", 135=>x"7c00", 136=>x"7900",
---- 137=>x"7c00", 138=>x"7800", 139=>x"7900", 140=>x"7600",
---- 141=>x"7700", 142=>x"7700", 143=>x"7700", 144=>x"7700",
---- 145=>x"7700", 146=>x"7500", 147=>x"7800", 148=>x"7900",
---- 149=>x"7900", 150=>x"7700", 151=>x"7700", 152=>x"8800",
---- 153=>x"7500", 154=>x"7700", 155=>x"7600", 156=>x"7800",
---- 157=>x"7900", 158=>x"7800", 159=>x"7800", 160=>x"7b00",
---- 161=>x"7900", 162=>x"7d00", 163=>x"7900", 164=>x"7900",
---- 165=>x"7600", 166=>x"7a00", 167=>x"7a00", 168=>x"7900",
---- 169=>x"7900", 170=>x"7900", 171=>x"7800", 172=>x"7800",
---- 173=>x"7800", 174=>x"7800", 175=>x"7800", 176=>x"7900",
---- 177=>x"7700", 178=>x"7900", 179=>x"7900", 180=>x"7a00",
---- 181=>x"7a00", 182=>x"7800", 183=>x"7c00", 184=>x"7900",
---- 185=>x"7c00", 186=>x"7800", 187=>x"7800", 188=>x"7600",
---- 189=>x"7800", 190=>x"7b00", 191=>x"7c00", 192=>x"7700",
---- 193=>x"7700", 194=>x"7800", 195=>x"7a00", 196=>x"8500",
---- 197=>x"7900", 198=>x"7800", 199=>x"7a00", 200=>x"7b00",
---- 201=>x"7700", 202=>x"7800", 203=>x"8500", 204=>x"7900",
---- 205=>x"7600", 206=>x"7a00", 207=>x"8900", 208=>x"7300",
---- 209=>x"7400", 210=>x"9400", 211=>x"8500", 212=>x"6f00",
---- 213=>x"8700", 214=>x"b600", 215=>x"7b00", 216=>x"6c00",
---- 217=>x"9f00", 218=>x"b300", 219=>x"7400", 220=>x"7400",
---- 221=>x"c000", 222=>x"a900", 223=>x"6900", 224=>x"9800",
---- 225=>x"cf00", 226=>x"9400", 227=>x"6400", 228=>x"be00",
---- 229=>x"c700", 230=>x"8a00", 231=>x"6100", 232=>x"d600",
---- 233=>x"b600", 234=>x"7a00", 235=>x"6000", 236=>x"d900",
---- 237=>x"a000", 238=>x"7b00", 239=>x"6600", 240=>x"c800",
---- 241=>x"a700", 242=>x"8400", 243=>x"6700", 244=>x"c300",
---- 245=>x"a200", 246=>x"7a00", 247=>x"6600", 248=>x"be00",
---- 249=>x"9600", 250=>x"7300", 251=>x"6000", 252=>x"b800",
---- 253=>x"9600", 254=>x"6e00", 255=>x"5c00", 256=>x"b100",
---- 257=>x"5e00", 258=>x"7200", 259=>x"5b00", 260=>x"b100",
---- 261=>x"8d00", 262=>x"7100", 263=>x"6200", 264=>x"a800",
---- 265=>x"8300", 266=>x"6f00", 267=>x"6200", 268=>x"9b00",
---- 269=>x"7b00", 270=>x"7000", 271=>x"6400", 272=>x"9300",
---- 273=>x"7400", 274=>x"7500", 275=>x"6a00", 276=>x"8900",
---- 277=>x"8300", 278=>x"7800", 279=>x"6c00", 280=>x"9200",
---- 281=>x"8200", 282=>x"7c00", 283=>x"6c00", 284=>x"9200",
---- 285=>x"8200", 286=>x"7e00", 287=>x"6b00", 288=>x"9e00",
---- 289=>x"8600", 290=>x"7f00", 291=>x"7100", 292=>x"9d00",
---- 293=>x"8b00", 294=>x"8000", 295=>x"7400", 296=>x"9d00",
---- 297=>x"9100", 298=>x"7a00", 299=>x"7700", 300=>x"9f00",
---- 301=>x"9400", 302=>x"8a00", 303=>x"8200", 304=>x"9900",
---- 305=>x"9000", 306=>x"8b00", 307=>x"8800", 308=>x"a000",
---- 309=>x"9d00", 310=>x"8800", 311=>x"9000", 312=>x"aa00",
---- 313=>x"a400", 314=>x"9a00", 315=>x"8b00", 316=>x"9c00",
---- 317=>x"a000", 318=>x"9500", 319=>x"8f00", 320=>x"a900",
---- 321=>x"9c00", 322=>x"ad00", 323=>x"9200", 324=>x"a200",
---- 325=>x"a000", 326=>x"9600", 327=>x"9400", 328=>x"b000",
---- 329=>x"9700", 330=>x"9800", 331=>x"9600", 332=>x"ae00",
---- 333=>x"a300", 334=>x"9400", 335=>x"9e00", 336=>x"b500",
---- 337=>x"a800", 338=>x"a200", 339=>x"9d00", 340=>x"b700",
---- 341=>x"a900", 342=>x"aa00", 343=>x"5d00", 344=>x"b300",
---- 345=>x"ac00", 346=>x"a100", 347=>x"a900", 348=>x"bc00",
---- 349=>x"a400", 350=>x"a800", 351=>x"9f00", 352=>x"ba00",
---- 353=>x"b600", 354=>x"a600", 355=>x"a600", 356=>x"c500",
---- 357=>x"b600", 358=>x"b600", 359=>x"a300", 360=>x"bd00",
---- 361=>x"c600", 362=>x"b100", 363=>x"a900", 364=>x"d000",
---- 365=>x"c200", 366=>x"b900", 367=>x"9e00", 368=>x"c400",
---- 369=>x"ca00", 370=>x"4600", 371=>x"ac00", 372=>x"ca00",
---- 373=>x"c600", 374=>x"bf00", 375=>x"a200", 376=>x"c500",
---- 377=>x"d100", 378=>x"c000", 379=>x"a200", 380=>x"c700",
---- 381=>x"c300", 382=>x"c400", 383=>x"a200", 384=>x"c000",
---- 385=>x"c500", 386=>x"be00", 387=>x"b700", 388=>x"c800",
---- 389=>x"bd00", 390=>x"ca00", 391=>x"b700", 392=>x"c100",
---- 393=>x"c900", 394=>x"c100", 395=>x"c600", 396=>x"cd00",
---- 397=>x"c500", 398=>x"c600", 399=>x"c500", 400=>x"cf00",
---- 401=>x"cd00", 402=>x"cc00", 403=>x"b400", 404=>x"de00",
---- 405=>x"d100", 406=>x"c900", 407=>x"c100", 408=>x"d100",
---- 409=>x"d200", 410=>x"d400", 411=>x"c300", 412=>x"9900",
---- 413=>x"e100", 414=>x"cf00", 415=>x"bf00", 416=>x"6600",
---- 417=>x"ca00", 418=>x"d200", 419=>x"c200", 420=>x"5100",
---- 421=>x"9f00", 422=>x"e100", 423=>x"cc00", 424=>x"5200",
---- 425=>x"8d00", 426=>x"df00", 427=>x"d900", 428=>x"5100",
---- 429=>x"8a00", 430=>x"dd00", 431=>x"d500", 432=>x"5300",
---- 433=>x"8800", 434=>x"e000", 435=>x"d500", 436=>x"5200",
---- 437=>x"8800", 438=>x"db00", 439=>x"d800", 440=>x"5900",
---- 441=>x"7900", 442=>x"d900", 443=>x"da00", 444=>x"6100",
---- 445=>x"6600", 446=>x"c600", 447=>x"dd00", 448=>x"6500",
---- 449=>x"5b00", 450=>x"a600", 451=>x"e100", 452=>x"6b00",
---- 453=>x"6100", 454=>x"8500", 455=>x"dd00", 456=>x"7000",
---- 457=>x"6b00", 458=>x"6c00", 459=>x"b900", 460=>x"7300",
---- 461=>x"6f00", 462=>x"6600", 463=>x"8800", 464=>x"7500",
---- 465=>x"7300", 466=>x"6e00", 467=>x"6f00", 468=>x"7900",
---- 469=>x"7400", 470=>x"7400", 471=>x"7000", 472=>x"7600",
---- 473=>x"7400", 474=>x"7700", 475=>x"8000", 476=>x"6800",
---- 477=>x"6a00", 478=>x"8400", 479=>x"8800", 480=>x"7700",
---- 481=>x"7a00", 482=>x"8d00", 483=>x"5f00", 484=>x"7400",
---- 485=>x"7500", 486=>x"a200", 487=>x"8a00", 488=>x"ac00",
---- 489=>x"9e00", 490=>x"9500", 491=>x"5000", 492=>x"c900",
---- 493=>x"7a00", 494=>x"5500", 495=>x"2100", 496=>x"b100",
---- 497=>x"5600", 498=>x"3200", 499=>x"3400", 500=>x"6100",
---- 501=>x"8600", 502=>x"4400", 503=>x"3100", 504=>x"9500",
---- 505=>x"8200", 506=>x"3100", 507=>x"3d00", 508=>x"9800",
---- 509=>x"af00", 510=>x"7100", 511=>x"7600", 512=>x"9700",
---- 513=>x"b500", 514=>x"ad00", 515=>x"a400", 516=>x"9a00",
---- 517=>x"9a00", 518=>x"7b00", 519=>x"7d00", 520=>x"9d00",
---- 521=>x"9100", 522=>x"6c00", 523=>x"4000", 524=>x"8800",
---- 525=>x"8300", 526=>x"5800", 527=>x"3b00", 528=>x"7800",
---- 529=>x"8500", 530=>x"5300", 531=>x"4c00", 532=>x"9900",
---- 533=>x"7d00", 534=>x"3700", 535=>x"3e00", 536=>x"6a00",
---- 537=>x"4200", 538=>x"2400", 539=>x"2800", 540=>x"2800",
---- 541=>x"2b00", 542=>x"2700", 543=>x"2a00", 544=>x"2b00",
---- 545=>x"2500", 546=>x"2200", 547=>x"3600", 548=>x"2500",
---- 549=>x"3200", 550=>x"4c00", 551=>x"7700", 552=>x"5200",
---- 553=>x"6a00", 554=>x"7600", 555=>x"5a00", 556=>x"7e00",
---- 557=>x"4800", 558=>x"3000", 559=>x"4800", 560=>x"8f00",
---- 561=>x"7a00", 562=>x"5600", 563=>x"8300", 564=>x"4600",
---- 565=>x"8d00", 566=>x"8f00", 567=>x"8600", 568=>x"4a00",
---- 569=>x"6800", 570=>x"6a00", 571=>x"6300", 572=>x"7300",
---- 573=>x"6900", 574=>x"3400", 575=>x"3a00", 576=>x"6f00",
---- 577=>x"5b00", 578=>x"3c00", 579=>x"6800", 580=>x"5e00",
---- 581=>x"6100", 582=>x"6d00", 583=>x"7600", 584=>x"6300",
---- 585=>x"7f00", 586=>x"7600", 587=>x"4f00", 588=>x"8a00",
---- 589=>x"8500", 590=>x"4900", 591=>x"2f00", 592=>x"5700",
---- 593=>x"4d00", 594=>x"4d00", 595=>x"2e00", 596=>x"4600",
---- 597=>x"4000", 598=>x"5800", 599=>x"3400", 600=>x"5d00",
---- 601=>x"4000", 602=>x"4600", 603=>x"3500", 604=>x"6400",
---- 605=>x"3800", 606=>x"3a00", 607=>x"3c00", 608=>x"7600",
---- 609=>x"5000", 610=>x"3100", 611=>x"3d00", 612=>x"6800",
---- 613=>x"6e00", 614=>x"3000", 615=>x"3500", 616=>x"5600",
---- 617=>x"8100", 618=>x"4200", 619=>x"c600", 620=>x"5d00",
---- 621=>x"7c00", 622=>x"5700", 623=>x"2e00", 624=>x"6200",
---- 625=>x"5000", 626=>x"5600", 627=>x"1f00", 628=>x"6c00",
---- 629=>x"3e00", 630=>x"6b00", 631=>x"2500", 632=>x"7e00",
---- 633=>x"3500", 634=>x"6f00", 635=>x"3f00", 636=>x"8700",
---- 637=>x"3000", 638=>x"5a00", 639=>x"5700", 640=>x"6400",
---- 641=>x"3a00", 642=>x"4d00", 643=>x"7f00", 644=>x"b100",
---- 645=>x"5d00", 646=>x"3d00", 647=>x"9200", 648=>x"a600",
---- 649=>x"8300", 650=>x"3000", 651=>x"8400", 652=>x"8900",
---- 653=>x"9600", 654=>x"3b00", 655=>x"8200", 656=>x"7800",
---- 657=>x"9c00", 658=>x"6200", 659=>x"7700", 660=>x"6800",
---- 661=>x"8100", 662=>x"8200", 663=>x"7900", 664=>x"5100",
---- 665=>x"6400", 666=>x"8c00", 667=>x"7c00", 668=>x"5f00",
---- 669=>x"a600", 670=>x"9200", 671=>x"6900", 672=>x"6900",
---- 673=>x"4d00", 674=>x"7600", 675=>x"6a00", 676=>x"5100",
---- 677=>x"4a00", 678=>x"6800", 679=>x"7c00", 680=>x"4800",
---- 681=>x"4100", 682=>x"6e00", 683=>x"8600", 684=>x"6000",
---- 685=>x"3700", 686=>x"3c00", 687=>x"7000", 688=>x"5e00",
---- 689=>x"5900", 690=>x"2e00", 691=>x"3f00", 692=>x"4300",
---- 693=>x"6900", 694=>x"5800", 695=>x"3200", 696=>x"4400",
---- 697=>x"4700", 698=>x"7000", 699=>x"5300", 700=>x"b200",
---- 701=>x"3e00", 702=>x"4900", 703=>x"6e00", 704=>x"6a00",
---- 705=>x"5900", 706=>x"4a00", 707=>x"5800", 708=>x"6600",
---- 709=>x"6a00", 710=>x"6300", 711=>x"5f00", 712=>x"6f00",
---- 713=>x"5f00", 714=>x"5100", 715=>x"5e00", 716=>x"6600",
---- 717=>x"7700", 718=>x"6300", 719=>x"5800", 720=>x"4000",
---- 721=>x"5c00", 722=>x"8200", 723=>x"6500", 724=>x"5200",
---- 725=>x"3b00", 726=>x"5d00", 727=>x"8200", 728=>x"6300",
---- 729=>x"4100", 730=>x"3900", 731=>x"5d00", 732=>x"6a00",
---- 733=>x"4900", 734=>x"4700", 735=>x"5000", 736=>x"7000",
---- 737=>x"5f00", 738=>x"7300", 739=>x"7200", 740=>x"6b00",
---- 741=>x"6d00", 742=>x"7f00", 743=>x"5000", 744=>x"7000",
---- 745=>x"7300", 746=>x"6400", 747=>x"5100", 748=>x"7c00",
---- 749=>x"7500", 750=>x"7200", 751=>x"6800", 752=>x"8200",
---- 753=>x"8500", 754=>x"7d00", 755=>x"7a00", 756=>x"8700",
---- 757=>x"8e00", 758=>x"7200", 759=>x"7b00", 760=>x"6a00",
---- 761=>x"7a00", 762=>x"7700", 763=>x"8400", 764=>x"6700",
---- 765=>x"6700", 766=>x"7400", 767=>x"7b00", 768=>x"5800",
---- 769=>x"7100", 770=>x"7500", 771=>x"5f00", 772=>x"4400",
---- 773=>x"7400", 774=>x"7a00", 775=>x"6c00", 776=>x"3800",
---- 777=>x"5b00", 778=>x"8c00", 779=>x"6f00", 780=>x"3500",
---- 781=>x"3a00", 782=>x"5a00", 783=>x"5b00", 784=>x"2d00",
---- 785=>x"2e00", 786=>x"5700", 787=>x"7500", 788=>x"2e00",
---- 789=>x"4000", 790=>x"5f00", 791=>x"7f00", 792=>x"7700",
---- 793=>x"7b00", 794=>x"7b00", 795=>x"9100", 796=>x"6100",
---- 797=>x"7300", 798=>x"7d00", 799=>x"9f00", 800=>x"4a00",
---- 801=>x"5000", 802=>x"5300", 803=>x"8c00", 804=>x"6e00",
---- 805=>x"5a00", 806=>x"7a00", 807=>x"8100", 808=>x"7000",
---- 809=>x"8000", 810=>x"8200", 811=>x"4e00", 812=>x"8100",
---- 813=>x"6c00", 814=>x"4b00", 815=>x"3900", 816=>x"6700",
---- 817=>x"3700", 818=>x"4200", 819=>x"4000", 820=>x"3f00",
---- 821=>x"3300", 822=>x"4200", 823=>x"4a00", 824=>x"5100",
---- 825=>x"2b00", 826=>x"3d00", 827=>x"5000", 828=>x"6d00",
---- 829=>x"3c00", 830=>x"3000", 831=>x"4600", 832=>x"6800",
---- 833=>x"6400", 834=>x"3500", 835=>x"3300", 836=>x"5a00",
---- 837=>x"5400", 838=>x"5a00", 839=>x"3700", 840=>x"a300",
---- 841=>x"4200", 842=>x"5200", 843=>x"5d00", 844=>x"5400",
---- 845=>x"4700", 846=>x"3900", 847=>x"6300", 848=>x"4a00",
---- 849=>x"5000", 850=>x"3100", 851=>x"4b00", 852=>x"6100",
---- 853=>x"5c00", 854=>x"3400", 855=>x"4200", 856=>x"3a00",
---- 857=>x"4600", 858=>x"cf00", 859=>x"4b00", 860=>x"2100",
---- 861=>x"3200", 862=>x"cc00", 863=>x"c000", 864=>x"2e00",
---- 865=>x"2f00", 866=>x"3100", 867=>x"3200", 868=>x"3000",
---- 869=>x"3400", 870=>x"3300", 871=>x"2c00", 872=>x"2b00",
---- 873=>x"3a00", 874=>x"3d00", 875=>x"2b00", 876=>x"2c00",
---- 877=>x"c500", 878=>x"4100", 879=>x"2600", 880=>x"2a00",
---- 881=>x"3a00", 882=>x"4500", 883=>x"2500", 884=>x"2e00",
---- 885=>x"4100", 886=>x"3a00", 887=>x"2b00", 888=>x"2f00",
---- 889=>x"3c00", 890=>x"4000", 891=>x"2d00", 892=>x"2700",
---- 893=>x"3800", 894=>x"3f00", 895=>x"2900", 896=>x"2700",
---- 897=>x"3f00", 898=>x"3300", 899=>x"2a00", 900=>x"2f00",
---- 901=>x"4000", 902=>x"2500", 903=>x"3800", 904=>x"3300",
---- 905=>x"4000", 906=>x"2500", 907=>x"4f00", 908=>x"3400",
---- 909=>x"3900", 910=>x"3900", 911=>x"4c00", 912=>x"2c00",
---- 913=>x"3400", 914=>x"6200", 915=>x"4300", 916=>x"2400",
---- 917=>x"3d00", 918=>x"6700", 919=>x"3c00", 920=>x"2300",
---- 921=>x"4a00", 922=>x"4f00", 923=>x"3000", 924=>x"2800",
---- 925=>x"4d00", 926=>x"3600", 927=>x"2e00", 928=>x"2b00",
---- 929=>x"3c00", 930=>x"3000", 931=>x"3500", 932=>x"3100",
---- 933=>x"2b00", 934=>x"3400", 935=>x"5c00", 936=>x"3400",
---- 937=>x"2e00", 938=>x"3800", 939=>x"4600", 940=>x"3800",
---- 941=>x"3800", 942=>x"3000", 943=>x"2500", 944=>x"2b00",
---- 945=>x"3900", 946=>x"3b00", 947=>x"2e00", 948=>x"2700",
---- 949=>x"2800", 950=>x"4100", 951=>x"3a00", 952=>x"3000",
---- 953=>x"2800", 954=>x"2e00", 955=>x"3900", 956=>x"3200",
---- 957=>x"3500", 958=>x"2200", 959=>x"3400", 960=>x"2d00",
---- 961=>x"3e00", 962=>x"3700", 963=>x"2700", 964=>x"2500",
---- 965=>x"3a00", 966=>x"4f00", 967=>x"3900", 968=>x"2500",
---- 969=>x"3300", 970=>x"5a00", 971=>x"5b00", 972=>x"2b00",
---- 973=>x"3100", 974=>x"5400", 975=>x"4f00", 976=>x"3300",
---- 977=>x"2c00", 978=>x"5500", 979=>x"4800", 980=>x"3100",
---- 981=>x"2b00", 982=>x"3d00", 983=>x"6400", 984=>x"3300",
---- 985=>x"3500", 986=>x"2d00", 987=>x"6000", 988=>x"2900",
---- 989=>x"2900", 990=>x"4500", 991=>x"5700", 992=>x"2900",
---- 993=>x"2400", 994=>x"3900", 995=>x"5e00", 996=>x"3c00",
---- 997=>x"2100", 998=>x"2700", 999=>x"5600", 1000=>x"6200",
---- 1001=>x"3400", 1002=>x"2a00", 1003=>x"4900", 1004=>x"8600",
---- 1005=>x"4400", 1006=>x"2800", 1007=>x"2d00", 1008=>x"9100",
---- 1009=>x"5800", 1010=>x"2600", 1011=>x"2800", 1012=>x"7d00",
---- 1013=>x"8500", 1014=>x"3600", 1015=>x"2700", 1016=>x"5200",
---- 1017=>x"7f00", 1018=>x"6400", 1019=>x"2b00", 1020=>x"4300",
---- 1021=>x"5300", 1022=>x"8400", 1023=>x"5500"),
----
---- 17 => (0=>x"8500", 1=>x"8600", 2=>x"8300", 3=>x"8000", 4=>x"8500",
---- 5=>x"8600", 6=>x"8400", 7=>x"8100", 8=>x"8400",
---- 9=>x"8500", 10=>x"8400", 11=>x"8200", 12=>x"8100",
---- 13=>x"8200", 14=>x"8400", 15=>x"8100", 16=>x"8300",
---- 17=>x"8200", 18=>x"8200", 19=>x"8200", 20=>x"8100",
---- 21=>x"8100", 22=>x"8000", 23=>x"8300", 24=>x"7e00",
---- 25=>x"8200", 26=>x"8100", 27=>x"8400", 28=>x"7d00",
---- 29=>x"8300", 30=>x"8300", 31=>x"8300", 32=>x"7f00",
---- 33=>x"8200", 34=>x"8200", 35=>x"8200", 36=>x"8100",
---- 37=>x"8100", 38=>x"8500", 39=>x"8400", 40=>x"8100",
---- 41=>x"8100", 42=>x"8300", 43=>x"8100", 44=>x"8200",
---- 45=>x"8000", 46=>x"8300", 47=>x"8100", 48=>x"8000",
---- 49=>x"8300", 50=>x"8100", 51=>x"8200", 52=>x"7f00",
---- 53=>x"8100", 54=>x"8100", 55=>x"8200", 56=>x"8100",
---- 57=>x"7e00", 58=>x"7e00", 59=>x"8100", 60=>x"7f00",
---- 61=>x"8000", 62=>x"7f00", 63=>x"7e00", 64=>x"7e00",
---- 65=>x"8100", 66=>x"8000", 67=>x"7f00", 68=>x"8000",
---- 69=>x"7f00", 70=>x"8000", 71=>x"8200", 72=>x"7f00",
---- 73=>x"7d00", 74=>x"8200", 75=>x"8100", 76=>x"7b00",
---- 77=>x"7b00", 78=>x"8100", 79=>x"8100", 80=>x"7e00",
---- 81=>x"7d00", 82=>x"7d00", 83=>x"7e00", 84=>x"7c00",
---- 85=>x"8000", 86=>x"7e00", 87=>x"7a00", 88=>x"8200",
---- 89=>x"7e00", 90=>x"7d00", 91=>x"7c00", 92=>x"7e00",
---- 93=>x"7f00", 94=>x"7d00", 95=>x"7b00", 96=>x"7f00",
---- 97=>x"7f00", 98=>x"8000", 99=>x"7f00", 100=>x"7d00",
---- 101=>x"7e00", 102=>x"7d00", 103=>x"7f00", 104=>x"7b00",
---- 105=>x"7d00", 106=>x"7d00", 107=>x"7d00", 108=>x"7c00",
---- 109=>x"7c00", 110=>x"8000", 111=>x"8100", 112=>x"7e00",
---- 113=>x"7d00", 114=>x"8000", 115=>x"8000", 116=>x"7700",
---- 117=>x"7e00", 118=>x"7e00", 119=>x"7b00", 120=>x"7b00",
---- 121=>x"7900", 122=>x"7e00", 123=>x"7e00", 124=>x"8300",
---- 125=>x"7c00", 126=>x"7c00", 127=>x"7d00", 128=>x"7800",
---- 129=>x"7a00", 130=>x"7c00", 131=>x"7e00", 132=>x"7b00",
---- 133=>x"7b00", 134=>x"7c00", 135=>x"7c00", 136=>x"7a00",
---- 137=>x"7d00", 138=>x"7a00", 139=>x"7b00", 140=>x"7b00",
---- 141=>x"7b00", 142=>x"7a00", 143=>x"7e00", 144=>x"7900",
---- 145=>x"7600", 146=>x"7b00", 147=>x"7b00", 148=>x"7900",
---- 149=>x"8500", 150=>x"7a00", 151=>x"7c00", 152=>x"7800",
---- 153=>x"7b00", 154=>x"7800", 155=>x"7900", 156=>x"7c00",
---- 157=>x"7a00", 158=>x"7900", 159=>x"7900", 160=>x"7b00",
---- 161=>x"7d00", 162=>x"7600", 163=>x"7700", 164=>x"7a00",
---- 165=>x"7700", 166=>x"7900", 167=>x"7b00", 168=>x"7c00",
---- 169=>x"7900", 170=>x"7d00", 171=>x"7b00", 172=>x"7b00",
---- 173=>x"7a00", 174=>x"7e00", 175=>x"7b00", 176=>x"7a00",
---- 177=>x"7b00", 178=>x"7b00", 179=>x"8100", 180=>x"7800",
---- 181=>x"7700", 182=>x"8100", 183=>x"8100", 184=>x"8400",
---- 185=>x"7b00", 186=>x"7f00", 187=>x"7200", 188=>x"7b00",
---- 189=>x"7f00", 190=>x"7900", 191=>x"7000", 192=>x"7f00",
---- 193=>x"7e00", 194=>x"7400", 195=>x"7500", 196=>x"8900",
---- 197=>x"7800", 198=>x"6f00", 199=>x"7100", 200=>x"8900",
---- 201=>x"6f00", 202=>x"6b00", 203=>x"6c00", 204=>x"7b00",
---- 205=>x"6d00", 206=>x"6e00", 207=>x"6900", 208=>x"6d00",
---- 209=>x"6900", 210=>x"6700", 211=>x"6500", 212=>x"6400",
---- 213=>x"6500", 214=>x"6800", 215=>x"6700", 216=>x"5f00",
---- 217=>x"6700", 218=>x"6b00", 219=>x"6c00", 220=>x"6200",
---- 221=>x"6700", 222=>x"6d00", 223=>x"6900", 224=>x"6600",
---- 225=>x"6900", 226=>x"6700", 227=>x"6900", 228=>x"6600",
---- 229=>x"6b00", 230=>x"6700", 231=>x"6700", 232=>x"6700",
---- 233=>x"6800", 234=>x"6600", 235=>x"6a00", 236=>x"6300",
---- 237=>x"6700", 238=>x"6700", 239=>x"6a00", 240=>x"6100",
---- 241=>x"6800", 242=>x"6800", 243=>x"6a00", 244=>x"9a00",
---- 245=>x"6200", 246=>x"6400", 247=>x"6a00", 248=>x"6100",
---- 249=>x"6600", 250=>x"6900", 251=>x"6800", 252=>x"6000",
---- 253=>x"6700", 254=>x"6600", 255=>x"6800", 256=>x"6400",
---- 257=>x"6700", 258=>x"6600", 259=>x"6d00", 260=>x"6800",
---- 261=>x"6700", 262=>x"6700", 263=>x"6b00", 264=>x"6100",
---- 265=>x"6200", 266=>x"6500", 267=>x"6700", 268=>x"5d00",
---- 269=>x"6100", 270=>x"6400", 271=>x"9a00", 272=>x"5f00",
---- 273=>x"6000", 274=>x"6400", 275=>x"6b00", 276=>x"6400",
---- 277=>x"6400", 278=>x"6800", 279=>x"6c00", 280=>x"6900",
---- 281=>x"6800", 282=>x"6900", 283=>x"6700", 284=>x"6600",
---- 285=>x"6d00", 286=>x"6800", 287=>x"6900", 288=>x"9800",
---- 289=>x"6800", 290=>x"6200", 291=>x"6b00", 292=>x"6a00",
---- 293=>x"6300", 294=>x"6c00", 295=>x"6d00", 296=>x"7000",
---- 297=>x"7000", 298=>x"6f00", 299=>x"6900", 300=>x"7b00",
---- 301=>x"7e00", 302=>x"6f00", 303=>x"6e00", 304=>x"7a00",
---- 305=>x"8000", 306=>x"7700", 307=>x"7300", 308=>x"8100",
---- 309=>x"8300", 310=>x"8100", 311=>x"6c00", 312=>x"9300",
---- 313=>x"8200", 314=>x"7e00", 315=>x"6f00", 316=>x"8d00",
---- 317=>x"8800", 318=>x"8400", 319=>x"7f00", 320=>x"8e00",
---- 321=>x"8700", 322=>x"8e00", 323=>x"8200", 324=>x"8e00",
---- 325=>x"8900", 326=>x"8c00", 327=>x"8400", 328=>x"9000",
---- 329=>x"7d00", 330=>x"8b00", 331=>x"8400", 332=>x"9400",
---- 333=>x"8b00", 334=>x"8d00", 335=>x"8e00", 336=>x"9a00",
---- 337=>x"8f00", 338=>x"8c00", 339=>x"9100", 340=>x"9b00",
---- 341=>x"8c00", 342=>x"9100", 343=>x"9800", 344=>x"9800",
---- 345=>x"a500", 346=>x"9200", 347=>x"9c00", 348=>x"a000",
---- 349=>x"9200", 350=>x"9f00", 351=>x"9400", 352=>x"9100",
---- 353=>x"9b00", 354=>x"8e00", 355=>x"a000", 356=>x"9800",
---- 357=>x"8400", 358=>x"6f00", 359=>x"9200", 360=>x"8c00",
---- 361=>x"7900", 362=>x"7b00", 363=>x"8f00", 364=>x"9200",
---- 365=>x"7c00", 366=>x"7a00", 367=>x"8900", 368=>x"8700",
---- 369=>x"7400", 370=>x"6f00", 371=>x"7b00", 372=>x"9300",
---- 373=>x"8800", 374=>x"6c00", 375=>x"9c00", 376=>x"8800",
---- 377=>x"7c00", 378=>x"8a00", 379=>x"9400", 380=>x"9400",
---- 381=>x"8400", 382=>x"8700", 383=>x"8a00", 384=>x"9b00",
---- 385=>x"8600", 386=>x"7400", 387=>x"9700", 388=>x"a800",
---- 389=>x"a000", 390=>x"8700", 391=>x"8600", 392=>x"ba00",
---- 393=>x"9c00", 394=>x"a900", 395=>x"8e00", 396=>x"a300",
---- 397=>x"ac00", 398=>x"aa00", 399=>x"a400", 400=>x"9f00",
---- 401=>x"af00", 402=>x"b400", 403=>x"a400", 404=>x"9d00",
---- 405=>x"a500", 406=>x"b400", 407=>x"b300", 408=>x"b400",
---- 409=>x"a800", 410=>x"b100", 411=>x"bf00", 412=>x"c400",
---- 413=>x"bb00", 414=>x"ba00", 415=>x"af00", 416=>x"c100",
---- 417=>x"bf00", 418=>x"c700", 419=>x"9600", 420=>x"c200",
---- 421=>x"bf00", 422=>x"ca00", 423=>x"9a00", 424=>x"c900",
---- 425=>x"c700", 426=>x"c600", 427=>x"b000", 428=>x"d300",
---- 429=>x"c800", 430=>x"c600", 431=>x"b100", 432=>x"2800",
---- 433=>x"d200", 434=>x"c500", 435=>x"8f00", 436=>x"d200",
---- 437=>x"d900", 438=>x"b100", 439=>x"6f00", 440=>x"d500",
---- 441=>x"d400", 442=>x"9400", 443=>x"6200", 444=>x"da00",
---- 445=>x"c500", 446=>x"7300", 447=>x"6900", 448=>x"dd00",
---- 449=>x"b700", 450=>x"6d00", 451=>x"6e00", 452=>x"e300",
---- 453=>x"a400", 454=>x"6f00", 455=>x"6f00", 456=>x"e900",
---- 457=>x"a800", 458=>x"6c00", 459=>x"7400", 460=>x"e300",
---- 461=>x"c000", 462=>x"7400", 463=>x"7500", 464=>x"c100",
---- 465=>x"d100", 466=>x"8100", 467=>x"7700", 468=>x"9000",
---- 469=>x"c700", 470=>x"8600", 471=>x"7900", 472=>x"7f00",
---- 473=>x"9400", 474=>x"7a00", 475=>x"7500", 476=>x"5c00",
---- 477=>x"6400", 478=>x"7500", 479=>x"6800", 480=>x"6000",
---- 481=>x"8300", 482=>x"9500", 483=>x"7300", 484=>x"7b00",
---- 485=>x"9400", 486=>x"bc00", 487=>x"9700", 488=>x"3d00",
---- 489=>x"4a00", 490=>x"5a00", 491=>x"7700", 492=>x"2000",
---- 493=>x"2200", 494=>x"2800", 495=>x"7400", 496=>x"2a00",
---- 497=>x"2a00", 498=>x"5200", 499=>x"7000", 500=>x"2400",
---- 501=>x"2700", 502=>x"5300", 503=>x"8f00", 504=>x"3e00",
---- 505=>x"1d00", 506=>x"4e00", 507=>x"8600", 508=>x"8d00",
---- 509=>x"4e00", 510=>x"6800", 511=>x"8100", 512=>x"ab00",
---- 513=>x"8900", 514=>x"6600", 515=>x"5200", 516=>x"9900",
---- 517=>x"6f00", 518=>x"3000", 519=>x"2b00", 520=>x"5600",
---- 521=>x"5d00", 522=>x"2c00", 523=>x"2400", 524=>x"4300",
---- 525=>x"3200", 526=>x"2600", 527=>x"1c00", 528=>x"2d00",
---- 529=>x"2700", 530=>x"2a00", 531=>x"3500", 532=>x"2500",
---- 533=>x"2c00", 534=>x"4b00", 535=>x"6400", 536=>x"2500",
---- 537=>x"4700", 538=>x"7300", 539=>x"4800", 540=>x"4100",
---- 541=>x"5f00", 542=>x"4500", 543=>x"3600", 544=>x"6000",
---- 545=>x"5400", 546=>x"4900", 547=>x"4b00", 548=>x"7a00",
---- 549=>x"6500", 550=>x"3900", 551=>x"2a00", 552=>x"5a00",
---- 553=>x"4e00", 554=>x"2000", 555=>x"2500", 556=>x"6b00",
---- 557=>x"2c00", 558=>x"2300", 559=>x"2c00", 560=>x"6e00",
---- 561=>x"af00", 562=>x"4300", 563=>x"3100", 564=>x"7a00",
---- 565=>x"7600", 566=>x"4b00", 567=>x"3200", 568=>x"6700",
---- 569=>x"5300", 570=>x"3200", 571=>x"2b00", 572=>x"6600",
---- 573=>x"5000", 574=>x"2800", 575=>x"2600", 576=>x"7100",
---- 577=>x"3200", 578=>x"2100", 579=>x"2a00", 580=>x"4400",
---- 581=>x"2400", 582=>x"2700", 583=>x"2700", 584=>x"2d00",
---- 585=>x"2d00", 586=>x"2e00", 587=>x"2700", 588=>x"3500",
---- 589=>x"3400", 590=>x"2e00", 591=>x"2f00", 592=>x"3700",
---- 593=>x"2e00", 594=>x"2e00", 595=>x"2e00", 596=>x"2f00",
---- 597=>x"2b00", 598=>x"2d00", 599=>x"3500", 600=>x"2900",
---- 601=>x"2e00", 602=>x"3700", 603=>x"3300", 604=>x"3300",
---- 605=>x"3300", 606=>x"3b00", 607=>x"3000", 608=>x"3a00",
---- 609=>x"3600", 610=>x"3e00", 611=>x"3400", 612=>x"3e00",
---- 613=>x"3e00", 614=>x"3b00", 615=>x"3100", 616=>x"4000",
---- 617=>x"3a00", 618=>x"3700", 619=>x"3100", 620=>x"3100",
---- 621=>x"c600", 622=>x"3800", 623=>x"3000", 624=>x"2b00",
---- 625=>x"2e00", 626=>x"3500", 627=>x"3200", 628=>x"2a00",
---- 629=>x"3200", 630=>x"2b00", 631=>x"3000", 632=>x"2200",
---- 633=>x"3000", 634=>x"2f00", 635=>x"4400", 636=>x"2800",
---- 637=>x"3b00", 638=>x"4500", 639=>x"3600", 640=>x"2f00",
---- 641=>x"3a00", 642=>x"3600", 643=>x"2900", 644=>x"4100",
---- 645=>x"2700", 646=>x"3000", 647=>x"3f00", 648=>x"4d00",
---- 649=>x"2600", 650=>x"3000", 651=>x"4900", 652=>x"6300",
---- 653=>x"1900", 654=>x"2600", 655=>x"2f00", 656=>x"7400",
---- 657=>x"1c00", 658=>x"2100", 659=>x"3400", 660=>x"8400",
---- 661=>x"3500", 662=>x"2000", 663=>x"3600", 664=>x"9200",
---- 665=>x"5800", 666=>x"2600", 667=>x"3300", 668=>x"8e00",
---- 669=>x"7500", 670=>x"4500", 671=>x"3d00", 672=>x"8900",
---- 673=>x"8000", 674=>x"5600", 675=>x"4600", 676=>x"8400",
---- 677=>x"8b00", 678=>x"9e00", 679=>x"3500", 680=>x"7600",
---- 681=>x"7b00", 682=>x"7a00", 683=>x"4900", 684=>x"8600",
---- 685=>x"6e00", 686=>x"7b00", 687=>x"8600", 688=>x"8100",
---- 689=>x"8300", 690=>x"7a00", 691=>x"9a00", 692=>x"4600",
---- 693=>x"5d00", 694=>x"7000", 695=>x"8800", 696=>x"3b00",
---- 697=>x"5d00", 698=>x"6400", 699=>x"7c00", 700=>x"6f00",
---- 701=>x"6e00", 702=>x"4200", 703=>x"6200", 704=>x"8e00",
---- 705=>x"7700", 706=>x"3800", 707=>x"4900", 708=>x"5b00",
---- 709=>x"5e00", 710=>x"5c00", 711=>x"4300", 712=>x"3b00",
---- 713=>x"3b00", 714=>x"6d00", 715=>x"6000", 716=>x"4500",
---- 717=>x"4200", 718=>x"5200", 719=>x"6300", 720=>x"6a00",
---- 721=>x"5600", 722=>x"6000", 723=>x"6000", 724=>x"7000",
---- 725=>x"7200", 726=>x"8a00", 727=>x"6e00", 728=>x"8200",
---- 729=>x"8600", 730=>x"6d00", 731=>x"7f00", 732=>x"8800",
---- 733=>x"8a00", 734=>x"7200", 735=>x"6f00", 736=>x"5b00",
---- 737=>x"7400", 738=>x"8400", 739=>x"6b00", 740=>x"4e00",
---- 741=>x"7000", 742=>x"8300", 743=>x"7500", 744=>x"ac00",
---- 745=>x"5500", 746=>x"7c00", 747=>x"7c00", 748=>x"5200",
---- 749=>x"4600", 750=>x"7c00", 751=>x"7e00", 752=>x"6800",
---- 753=>x"4700", 754=>x"7800", 755=>x"8a00", 756=>x"8200",
---- 757=>x"6700", 758=>x"7300", 759=>x"9100", 760=>x"8c00",
---- 761=>x"7300", 762=>x"6c00", 763=>x"7a00", 764=>x"8f00",
---- 765=>x"8a00", 766=>x"8800", 767=>x"7500", 768=>x"6d00",
---- 769=>x"9600", 770=>x"7800", 771=>x"7800", 772=>x"4f00",
---- 773=>x"7600", 774=>x"5e00", 775=>x"7b00", 776=>x"3e00",
---- 777=>x"6b00", 778=>x"8100", 779=>x"a300", 780=>x"5300",
---- 781=>x"8c00", 782=>x"6600", 783=>x"5800", 784=>x"7400",
---- 785=>x"9e00", 786=>x"7600", 787=>x"5800", 788=>x"9200",
---- 789=>x"9500", 790=>x"4e00", 791=>x"5a00", 792=>x"a300",
---- 793=>x"6000", 794=>x"4a00", 795=>x"4f00", 796=>x"7a00",
---- 797=>x"4300", 798=>x"5400", 799=>x"6500", 800=>x"4600",
---- 801=>x"5900", 802=>x"6c00", 803=>x"6100", 804=>x"4100",
---- 805=>x"4400", 806=>x"8d00", 807=>x"7200", 808=>x"4400",
---- 809=>x"4b00", 810=>x"4700", 811=>x"7600", 812=>x"4500",
---- 813=>x"5300", 814=>x"4c00", 815=>x"5100", 816=>x"3700",
---- 817=>x"4f00", 818=>x"6500", 819=>x"4e00", 820=>x"3d00",
---- 821=>x"3e00", 822=>x"5f00", 823=>x"9900", 824=>x"4d00",
---- 825=>x"4400", 826=>x"4700", 827=>x"9300", 828=>x"4200",
---- 829=>x"4c00", 830=>x"4b00", 831=>x"5300", 832=>x"4600",
---- 833=>x"4a00", 834=>x"4700", 835=>x"4500", 836=>x"4100",
---- 837=>x"5000", 838=>x"4c00", 839=>x"b700", 840=>x"3900",
---- 841=>x"5800", 842=>x"6100", 843=>x"4c00", 844=>x"5800",
---- 845=>x"4f00", 846=>x"6900", 847=>x"6500", 848=>x"5b00",
---- 849=>x"5400", 850=>x"5d00", 851=>x"7400", 852=>x"4400",
---- 853=>x"5d00", 854=>x"5700", 855=>x"7200", 856=>x"4500",
---- 857=>x"5400", 858=>x"5f00", 859=>x"6400", 860=>x"5200",
---- 861=>x"4500", 862=>x"6700", 863=>x"6000", 864=>x"4c00",
---- 865=>x"4300", 866=>x"5900", 867=>x"5c00", 868=>x"4100",
---- 869=>x"4400", 870=>x"4d00", 871=>x"4f00", 872=>x"3b00",
---- 873=>x"4400", 874=>x"3b00", 875=>x"3700", 876=>x"3600",
---- 877=>x"4b00", 878=>x"3700", 879=>x"4300", 880=>x"2f00",
---- 881=>x"5c00", 882=>x"3900", 883=>x"3700", 884=>x"3500",
---- 885=>x"5c00", 886=>x"4300", 887=>x"2d00", 888=>x"4d00",
---- 889=>x"5d00", 890=>x"3b00", 891=>x"3500", 892=>x"5800",
---- 893=>x"6300", 894=>x"2700", 895=>x"4000", 896=>x"5900",
---- 897=>x"6100", 898=>x"2500", 899=>x"3200", 900=>x"5700",
---- 901=>x"4a00", 902=>x"5300", 903=>x"2800", 904=>x"5600",
---- 905=>x"3400", 906=>x"6000", 907=>x"5300", 908=>x"4300",
---- 909=>x"3b00", 910=>x"4c00", 911=>x"6900", 912=>x"2d00",
---- 913=>x"3700", 914=>x"3600", 915=>x"6400", 916=>x"2600",
---- 917=>x"2e00", 918=>x"3b00", 919=>x"6400", 920=>x"2f00",
---- 921=>x"2b00", 922=>x"4c00", 923=>x"7800", 924=>x"4200",
---- 925=>x"3100", 926=>x"3b00", 927=>x"7000", 928=>x"4800",
---- 929=>x"6100", 930=>x"5800", 931=>x"6100", 932=>x"2700",
---- 933=>x"5300", 934=>x"7a00", 935=>x"5d00", 936=>x"1e00",
---- 937=>x"2900", 938=>x"5e00", 939=>x"5100", 940=>x"2b00",
---- 941=>x"2e00", 942=>x"2f00", 943=>x"5800", 944=>x"3400",
---- 945=>x"cc00", 946=>x"2300", 947=>x"3300", 948=>x"2b00",
---- 949=>x"3a00", 950=>x"2e00", 951=>x"2b00", 952=>x"3100",
---- 953=>x"4a00", 954=>x"3c00", 955=>x"3100", 956=>x"4600",
---- 957=>x"3f00", 958=>x"4000", 959=>x"3000", 960=>x"3d00",
---- 961=>x"4400", 962=>x"4000", 963=>x"3700", 964=>x"2800",
---- 965=>x"3c00", 966=>x"4c00", 967=>x"3400", 968=>x"cb00",
---- 969=>x"3000", 970=>x"5300", 971=>x"3e00", 972=>x"4600",
---- 973=>x"3800", 974=>x"4100", 975=>x"5500", 976=>x"2d00",
---- 977=>x"3400", 978=>x"2f00", 979=>x"6f00", 980=>x"2b00",
---- 981=>x"2c00", 982=>x"3a00", 983=>x"5500", 984=>x"4700",
---- 985=>x"2a00", 986=>x"3300", 987=>x"3600", 988=>x"7100",
---- 989=>x"2a00", 990=>x"1e00", 991=>x"3d00", 992=>x"7a00",
---- 993=>x"5200", 994=>x"1c00", 995=>x"3100", 996=>x"7800",
---- 997=>x"7000", 998=>x"2e00", 999=>x"1c00", 1000=>x"7100",
---- 1001=>x"6e00", 1002=>x"4800", 1003=>x"2800", 1004=>x"5300",
---- 1005=>x"6d00", 1006=>x"4200", 1007=>x"3f00", 1008=>x"3500",
---- 1009=>x"6c00", 1010=>x"4b00", 1011=>x"3800", 1012=>x"3b00",
---- 1013=>x"6e00", 1014=>x"6d00", 1015=>x"3400", 1016=>x"3900",
---- 1017=>x"7400", 1018=>x"7800", 1019=>x"4000", 1020=>x"2e00",
---- 1021=>x"7700", 1022=>x"7000", 1023=>x"3100"),
----
---- 18 => (0=>x"8300", 1=>x"7f00", 2=>x"8400", 3=>x"8200", 4=>x"8200",
---- 5=>x"7f00", 6=>x"8300", 7=>x"8200", 8=>x"8300",
---- 9=>x"7e00", 10=>x"8300", 11=>x"8200", 12=>x"8100",
---- 13=>x"8300", 14=>x"7b00", 15=>x"8200", 16=>x"8300",
---- 17=>x"8200", 18=>x"8300", 19=>x"8200", 20=>x"8300",
---- 21=>x"8300", 22=>x"8300", 23=>x"8000", 24=>x"8400",
---- 25=>x"8400", 26=>x"8200", 27=>x"8100", 28=>x"8200",
---- 29=>x"7c00", 30=>x"8200", 31=>x"8100", 32=>x"8300",
---- 33=>x"8300", 34=>x"8200", 35=>x"8300", 36=>x"8100",
---- 37=>x"8300", 38=>x"8500", 39=>x"8400", 40=>x"8000",
---- 41=>x"8500", 42=>x"8200", 43=>x"8300", 44=>x"8100",
---- 45=>x"8200", 46=>x"8200", 47=>x"8000", 48=>x"8200",
---- 49=>x"8100", 50=>x"8200", 51=>x"8400", 52=>x"8000",
---- 53=>x"8000", 54=>x"7f00", 55=>x"8100", 56=>x"7f00",
---- 57=>x"7f00", 58=>x"8200", 59=>x"8000", 60=>x"7f00",
---- 61=>x"7d00", 62=>x"8000", 63=>x"8000", 64=>x"7e00",
---- 65=>x"7c00", 66=>x"7f00", 67=>x"8100", 68=>x"7f00",
---- 69=>x"8100", 70=>x"7f00", 71=>x"7f00", 72=>x"7f00",
---- 73=>x"8000", 74=>x"7c00", 75=>x"7e00", 76=>x"7d00",
---- 77=>x"7d00", 78=>x"7a00", 79=>x"7e00", 80=>x"8000",
---- 81=>x"7c00", 82=>x"7b00", 83=>x"7c00", 84=>x"7c00",
---- 85=>x"7d00", 86=>x"7e00", 87=>x"7e00", 88=>x"7c00",
---- 89=>x"7d00", 90=>x"7d00", 91=>x"8000", 92=>x"7e00",
---- 93=>x"8000", 94=>x"7f00", 95=>x"8300", 96=>x"7d00",
---- 97=>x"7e00", 98=>x"7f00", 99=>x"8100", 100=>x"7e00",
---- 101=>x"8100", 102=>x"8200", 103=>x"8000", 104=>x"7e00",
---- 105=>x"8400", 106=>x"8100", 107=>x"8000", 108=>x"8300",
---- 109=>x"8200", 110=>x"7e00", 111=>x"7e00", 112=>x"7f00",
---- 113=>x"7d00", 114=>x"8100", 115=>x"7e00", 116=>x"7d00",
---- 117=>x"7f00", 118=>x"7d00", 119=>x"7e00", 120=>x"7c00",
---- 121=>x"8000", 122=>x"7e00", 123=>x"8000", 124=>x"7f00",
---- 125=>x"7e00", 126=>x"7e00", 127=>x"7d00", 128=>x"7d00",
---- 129=>x"7a00", 130=>x"7d00", 131=>x"7c00", 132=>x"7d00",
---- 133=>x"8300", 134=>x"7d00", 135=>x"7a00", 136=>x"7c00",
---- 137=>x"7c00", 138=>x"7c00", 139=>x"7c00", 140=>x"7f00",
---- 141=>x"7a00", 142=>x"7e00", 143=>x"7f00", 144=>x"7d00",
---- 145=>x"7900", 146=>x"7a00", 147=>x"7700", 148=>x"7c00",
---- 149=>x"7b00", 150=>x"7a00", 151=>x"7900", 152=>x"7d00",
---- 153=>x"7d00", 154=>x"7600", 155=>x"8a00", 156=>x"7c00",
---- 157=>x"7c00", 158=>x"7900", 159=>x"9500", 160=>x"7c00",
---- 161=>x"7e00", 162=>x"8300", 163=>x"8500", 164=>x"7c00",
---- 165=>x"7d00", 166=>x"8200", 167=>x"7b00", 168=>x"7c00",
---- 169=>x"8400", 170=>x"7c00", 171=>x"6d00", 172=>x"7e00",
---- 173=>x"8000", 174=>x"7000", 175=>x"6800", 176=>x"7c00",
---- 177=>x"7200", 178=>x"6e00", 179=>x"6c00", 180=>x"7000",
---- 181=>x"6c00", 182=>x"6a00", 183=>x"6b00", 184=>x"6a00",
---- 185=>x"6e00", 186=>x"6b00", 187=>x"6e00", 188=>x"6d00",
---- 189=>x"6900", 190=>x"6f00", 191=>x"7500", 192=>x"6f00",
---- 193=>x"7000", 194=>x"6e00", 195=>x"7100", 196=>x"7200",
---- 197=>x"7500", 198=>x"6e00", 199=>x"9200", 200=>x"6d00",
---- 201=>x"7400", 202=>x"7400", 203=>x"6d00", 204=>x"6b00",
---- 205=>x"7100", 206=>x"7400", 207=>x"7100", 208=>x"6700",
---- 209=>x"6c00", 210=>x"7600", 211=>x"7400", 212=>x"6900",
---- 213=>x"6c00", 214=>x"7000", 215=>x"7100", 216=>x"6800",
---- 217=>x"7200", 218=>x"6f00", 219=>x"7000", 220=>x"6c00",
---- 221=>x"6d00", 222=>x"6d00", 223=>x"7100", 224=>x"6c00",
---- 225=>x"6d00", 226=>x"6b00", 227=>x"6f00", 228=>x"6900",
---- 229=>x"7000", 230=>x"6f00", 231=>x"6d00", 232=>x"6b00",
---- 233=>x"6c00", 234=>x"7400", 235=>x"7700", 236=>x"6e00",
---- 237=>x"6d00", 238=>x"7000", 239=>x"7400", 240=>x"7000",
---- 241=>x"6c00", 242=>x"6900", 243=>x"7400", 244=>x"6e00",
---- 245=>x"6700", 246=>x"6f00", 247=>x"7b00", 248=>x"6900",
---- 249=>x"6d00", 250=>x"7200", 251=>x"8600", 252=>x"6a00",
---- 253=>x"7200", 254=>x"7400", 255=>x"6b00", 256=>x"6d00",
---- 257=>x"9500", 258=>x"6600", 259=>x"5e00", 260=>x"6a00",
---- 261=>x"5e00", 262=>x"5b00", 263=>x"7300", 264=>x"6300",
---- 265=>x"6400", 266=>x"7000", 267=>x"7b00", 268=>x"6a00",
---- 269=>x"7200", 270=>x"6f00", 271=>x"6f00", 272=>x"6e00",
---- 273=>x"8e00", 274=>x"6500", 275=>x"6d00", 276=>x"6a00",
---- 277=>x"6400", 278=>x"6700", 279=>x"6000", 280=>x"6100",
---- 281=>x"6500", 282=>x"6000", 283=>x"6800", 284=>x"6f00",
---- 285=>x"6700", 286=>x"6600", 287=>x"6a00", 288=>x"6b00",
---- 289=>x"6e00", 290=>x"6900", 291=>x"6c00", 292=>x"6a00",
---- 293=>x"6300", 294=>x"6900", 295=>x"7000", 296=>x"6600",
---- 297=>x"6600", 298=>x"6a00", 299=>x"6e00", 300=>x"6d00",
---- 301=>x"6900", 302=>x"6900", 303=>x"6900", 304=>x"6900",
---- 305=>x"6a00", 306=>x"6800", 307=>x"6d00", 308=>x"6800",
---- 309=>x"6800", 310=>x"6a00", 311=>x"6b00", 312=>x"7300",
---- 313=>x"7000", 314=>x"5e00", 315=>x"5a00", 316=>x"7800",
---- 317=>x"6700", 318=>x"5c00", 319=>x"6300", 320=>x"7000",
---- 321=>x"6600", 322=>x"6700", 323=>x"5b00", 324=>x"6a00",
---- 325=>x"6b00", 326=>x"6200", 327=>x"6600", 328=>x"7400",
---- 329=>x"7200", 330=>x"6b00", 331=>x"6900", 332=>x"7900",
---- 333=>x"7b00", 334=>x"7200", 335=>x"6a00", 336=>x"8100",
---- 337=>x"7700", 338=>x"6a00", 339=>x"9600", 340=>x"8e00",
---- 341=>x"7c00", 342=>x"7100", 343=>x"a600", 344=>x"9200",
---- 345=>x"8700", 346=>x"6c00", 347=>x"6200", 348=>x"9d00",
---- 349=>x"8600", 350=>x"7100", 351=>x"7a00", 352=>x"9300",
---- 353=>x"8800", 354=>x"7b00", 355=>x"7500", 356=>x"9f00",
---- 357=>x"9600", 358=>x"7300", 359=>x"6d00", 360=>x"9c00",
---- 361=>x"7800", 362=>x"6900", 363=>x"6c00", 364=>x"7f00",
---- 365=>x"7400", 366=>x"7100", 367=>x"7000", 368=>x"8800",
---- 369=>x"8100", 370=>x"7300", 371=>x"8800", 372=>x"8f00",
---- 373=>x"9300", 374=>x"7e00", 375=>x"7900", 376=>x"9500",
---- 377=>x"8200", 378=>x"8f00", 379=>x"7f00", 380=>x"9200",
---- 381=>x"9600", 382=>x"8900", 383=>x"8400", 384=>x"8c00",
---- 385=>x"9800", 386=>x"8e00", 387=>x"6c00", 388=>x"9a00",
---- 389=>x"7d00", 390=>x"7700", 391=>x"6b00", 392=>x"a100",
---- 393=>x"8c00", 394=>x"6400", 395=>x"6900", 396=>x"9100",
---- 397=>x"8e00", 398=>x"5e00", 399=>x"7100", 400=>x"8c00",
---- 401=>x"6000", 402=>x"6300", 403=>x"7e00", 404=>x"9300",
---- 405=>x"5c00", 406=>x"7100", 407=>x"8c00", 408=>x"9000",
---- 409=>x"6e00", 410=>x"8400", 411=>x"8400", 412=>x"6d00",
---- 413=>x"8200", 414=>x"8c00", 415=>x"7400", 416=>x"6b00",
---- 417=>x"9400", 418=>x"7f00", 419=>x"7100", 420=>x"8800",
---- 421=>x"8c00", 422=>x"7700", 423=>x"7300", 424=>x"9400",
---- 425=>x"7800", 426=>x"8300", 427=>x"7d00", 428=>x"8600",
---- 429=>x"7800", 430=>x"7c00", 431=>x"7e00", 432=>x"6900",
---- 433=>x"7400", 434=>x"7e00", 435=>x"7800", 436=>x"6300",
---- 437=>x"7600", 438=>x"7b00", 439=>x"7400", 440=>x"6600",
---- 441=>x"6e00", 442=>x"7300", 443=>x"7000", 444=>x"6c00",
---- 445=>x"6900", 446=>x"6b00", 447=>x"7400", 448=>x"7200",
---- 449=>x"7300", 450=>x"6e00", 451=>x"7300", 452=>x"7700",
---- 453=>x"7a00", 454=>x"7400", 455=>x"6800", 456=>x"7300",
---- 457=>x"7700", 458=>x"7600", 459=>x"6900", 460=>x"7000",
---- 461=>x"6b00", 462=>x"7300", 463=>x"7f00", 464=>x"7300",
---- 465=>x"6900", 466=>x"7b00", 467=>x"8300", 468=>x"6a00",
---- 469=>x"7300", 470=>x"7800", 471=>x"8500", 472=>x"7100",
---- 473=>x"8300", 474=>x"8900", 475=>x"8700", 476=>x"8100",
---- 477=>x"7f00", 478=>x"8600", 479=>x"7400", 480=>x"7800",
---- 481=>x"7f00", 482=>x"7f00", 483=>x"8100", 484=>x"7100",
---- 485=>x"7b00", 486=>x"7f00", 487=>x"8500", 488=>x"8200",
---- 489=>x"7800", 490=>x"8100", 491=>x"7f00", 492=>x"9d00",
---- 493=>x"ac00", 494=>x"8400", 495=>x"6e00", 496=>x"b300",
---- 497=>x"c100", 498=>x"8800", 499=>x"5800", 500=>x"8c00",
---- 501=>x"6000", 502=>x"6a00", 503=>x"4800", 504=>x"7e00",
---- 505=>x"5500", 506=>x"ac00", 507=>x"5c00", 508=>x"9000",
---- 509=>x"7000", 510=>x"4100", 511=>x"4900", 512=>x"5800",
---- 513=>x"4100", 514=>x"3900", 515=>x"3800", 516=>x"2100",
---- 517=>x"2200", 518=>x"bf00", 519=>x"5200", 520=>x"1f00",
---- 521=>x"4100", 522=>x"7100", 523=>x"5b00", 524=>x"4400",
---- 525=>x"7f00", 526=>x"5c00", 527=>x"3100", 528=>x"7600",
---- 529=>x"5f00", 530=>x"2300", 531=>x"4400", 532=>x"4600",
---- 533=>x"2600", 534=>x"c700", 535=>x"5a00", 536=>x"2500",
---- 537=>x"3900", 538=>x"5000", 539=>x"3800", 540=>x"3400",
---- 541=>x"4900", 542=>x"4600", 543=>x"3700", 544=>x"3600",
---- 545=>x"3f00", 546=>x"5200", 547=>x"4a00", 548=>x"2100",
---- 549=>x"4500", 550=>x"4700", 551=>x"5400", 552=>x"2700",
---- 553=>x"5f00", 554=>x"3f00", 555=>x"4f00", 556=>x"3000",
---- 557=>x"5e00", 558=>x"4900", 559=>x"4e00", 560=>x"2700",
---- 561=>x"4d00", 562=>x"4e00", 563=>x"4300", 564=>x"2700",
---- 565=>x"3900", 566=>x"5600", 567=>x"3d00", 568=>x"2600",
---- 569=>x"3700", 570=>x"4900", 571=>x"4200", 572=>x"3000",
---- 573=>x"3400", 574=>x"4900", 575=>x"5a00", 576=>x"2e00",
---- 577=>x"3700", 578=>x"5f00", 579=>x"7900", 580=>x"3000",
---- 581=>x"3000", 582=>x"3a00", 583=>x"6000", 584=>x"2c00",
---- 585=>x"d300", 586=>x"2a00", 587=>x"3d00", 588=>x"2e00",
---- 589=>x"2e00", 590=>x"2e00", 591=>x"3000", 592=>x"d200",
---- 593=>x"2d00", 594=>x"3300", 595=>x"3300", 596=>x"3200",
---- 597=>x"2e00", 598=>x"cb00", 599=>x"3300", 600=>x"3500",
---- 601=>x"3200", 602=>x"3100", 603=>x"3200", 604=>x"2e00",
---- 605=>x"3300", 606=>x"2e00", 607=>x"2f00", 608=>x"2e00",
---- 609=>x"2d00", 610=>x"2a00", 611=>x"2f00", 612=>x"d800",
---- 613=>x"2800", 614=>x"2800", 615=>x"2c00", 616=>x"2500",
---- 617=>x"2700", 618=>x"2200", 619=>x"2600", 620=>x"2400",
---- 621=>x"2900", 622=>x"2400", 623=>x"3400", 624=>x"2900",
---- 625=>x"2a00", 626=>x"2800", 627=>x"3000", 628=>x"3500",
---- 629=>x"3300", 630=>x"2f00", 631=>x"2a00", 632=>x"3e00",
---- 633=>x"2800", 634=>x"2200", 635=>x"2900", 636=>x"2c00",
---- 637=>x"3500", 638=>x"2800", 639=>x"2800", 640=>x"3000",
---- 641=>x"4d00", 642=>x"2c00", 643=>x"2100", 644=>x"3900",
---- 645=>x"5000", 646=>x"2d00", 647=>x"2200", 648=>x"4d00",
---- 649=>x"3c00", 650=>x"2f00", 651=>x"2200", 652=>x"3100",
---- 653=>x"5200", 654=>x"7100", 655=>x"3800", 656=>x"2600",
---- 657=>x"6b00", 658=>x"a900", 659=>x"6000", 660=>x"2a00",
---- 661=>x"6000", 662=>x"a500", 663=>x"9c00", 664=>x"3100",
---- 665=>x"4f00", 666=>x"8900", 667=>x"7a00", 668=>x"4700",
---- 669=>x"4c00", 670=>x"6f00", 671=>x"5e00", 672=>x"5e00",
---- 673=>x"5800", 674=>x"5900", 675=>x"5a00", 676=>x"7000",
---- 677=>x"6c00", 678=>x"4000", 679=>x"4000", 680=>x"9600",
---- 681=>x"5f00", 682=>x"2d00", 683=>x"2a00", 684=>x"9400",
---- 685=>x"3600", 686=>x"2700", 687=>x"2c00", 688=>x"5e00",
---- 689=>x"1b00", 690=>x"2200", 691=>x"3200", 692=>x"7b00",
---- 693=>x"3a00", 694=>x"1b00", 695=>x"5200", 696=>x"7300",
---- 697=>x"6d00", 698=>x"5a00", 699=>x"9000", 700=>x"5900",
---- 701=>x"4600", 702=>x"8300", 703=>x"9900", 704=>x"3900",
---- 705=>x"4400", 706=>x"7100", 707=>x"8100", 708=>x"5500",
---- 709=>x"6b00", 710=>x"9200", 711=>x"9500", 712=>x"7400",
---- 713=>x"7e00", 714=>x"9200", 715=>x"9600", 716=>x"8100",
---- 717=>x"8200", 718=>x"8f00", 719=>x"9600", 720=>x"8600",
---- 721=>x"9800", 722=>x"8d00", 723=>x"9900", 724=>x"9100",
---- 725=>x"a700", 726=>x"9f00", 727=>x"8f00", 728=>x"6300",
---- 729=>x"8000", 730=>x"9300", 731=>x"8700", 732=>x"5f00",
---- 733=>x"6800", 734=>x"7600", 735=>x"7400", 736=>x"4500",
---- 737=>x"7200", 738=>x"7f00", 739=>x"6d00", 740=>x"3200",
---- 741=>x"6400", 742=>x"7b00", 743=>x"7300", 744=>x"5f00",
---- 745=>x"7900", 746=>x"6100", 747=>x"6000", 748=>x"6f00",
---- 749=>x"8c00", 750=>x"5e00", 751=>x"4f00", 752=>x"6100",
---- 753=>x"9600", 754=>x"6f00", 755=>x"3a00", 756=>x"7600",
---- 757=>x"9300", 758=>x"7d00", 759=>x"5700", 760=>x"8800",
---- 761=>x"9500", 762=>x"6a00", 763=>x"5f00", 764=>x"7e00",
---- 765=>x"9300", 766=>x"9f00", 767=>x"5600", 768=>x"7f00",
---- 769=>x"9600", 770=>x"a800", 771=>x"7c00", 772=>x"8f00",
---- 773=>x"9d00", 774=>x"9000", 775=>x"8700", 776=>x"8200",
---- 777=>x"9e00", 778=>x"9100", 779=>x"7200", 780=>x"5800",
---- 781=>x"9400", 782=>x"a100", 783=>x"8800", 784=>x"5b00",
---- 785=>x"7c00", 786=>x"9400", 787=>x"7e00", 788=>x"6000",
---- 789=>x"5c00", 790=>x"7200", 791=>x"7e00", 792=>x"6900",
---- 793=>x"5f00", 794=>x"5c00", 795=>x"8200", 796=>x"5300",
---- 797=>x"6d00", 798=>x"7000", 799=>x"6900", 800=>x"6300",
---- 801=>x"6400", 802=>x"7600", 803=>x"7600", 804=>x"6900",
---- 805=>x"6f00", 806=>x"5300", 807=>x"8a00", 808=>x"7700",
---- 809=>x"7700", 810=>x"5b00", 811=>x"7300", 812=>x"7700",
---- 813=>x"7a00", 814=>x"7500", 815=>x"8500", 816=>x"6000",
---- 817=>x"7900", 818=>x"7d00", 819=>x"8a00", 820=>x"5600",
---- 821=>x"5c00", 822=>x"7000", 823=>x"8100", 824=>x"6200",
---- 825=>x"5200", 826=>x"5a00", 827=>x"7e00", 828=>x"7400",
---- 829=>x"6000", 830=>x"5100", 831=>x"7400", 832=>x"6700",
---- 833=>x"7200", 834=>x"5400", 835=>x"6f00", 836=>x"4b00",
---- 837=>x"6d00", 838=>x"5d00", 839=>x"7100", 840=>x"3d00",
---- 841=>x"5000", 842=>x"5f00", 843=>x"7500", 844=>x"5c00",
---- 845=>x"4300", 846=>x"4d00", 847=>x"7200", 848=>x"7600",
---- 849=>x"6500", 850=>x"4300", 851=>x"5e00", 852=>x"6a00",
---- 853=>x"6600", 854=>x"4f00", 855=>x"5500", 856=>x"6500",
---- 857=>x"5700", 858=>x"4e00", 859=>x"5800", 860=>x"6f00",
---- 861=>x"5d00", 862=>x"5700", 863=>x"4c00", 864=>x"7700",
---- 865=>x"6500", 866=>x"5200", 867=>x"4f00", 868=>x"8100",
---- 869=>x"7200", 870=>x"3f00", 871=>x"3b00", 872=>x"6b00",
---- 873=>x"8500", 874=>x"4700", 875=>x"3600", 876=>x"7200",
---- 877=>x"7600", 878=>x"6900", 879=>x"5800", 880=>x"4e00",
---- 881=>x"5400", 882=>x"7000", 883=>x"7e00", 884=>x"2c00",
---- 885=>x"3500", 886=>x"4a00", 887=>x"7500", 888=>x"2200",
---- 889=>x"2c00", 890=>x"3f00", 891=>x"6e00", 892=>x"2700",
---- 893=>x"2d00", 894=>x"4400", 895=>x"6700", 896=>x"5100",
---- 897=>x"3d00", 898=>x"5000", 899=>x"6100", 900=>x"5500",
---- 901=>x"5b00", 902=>x"4e00", 903=>x"6200", 904=>x"2a00",
---- 905=>x"5e00", 906=>x"6900", 907=>x"5000", 908=>x"2e00",
---- 909=>x"2800", 910=>x"7400", 911=>x"9a00", 912=>x"5600",
---- 913=>x"2100", 914=>x"3200", 915=>x"6d00", 916=>x"6100",
---- 917=>x"4300", 918=>x"3100", 919=>x"2700", 920=>x"7800",
---- 921=>x"4d00", 922=>x"4700", 923=>x"3800", 924=>x"8000",
---- 925=>x"7600", 926=>x"3a00", 927=>x"4400", 928=>x"7c00",
---- 929=>x"9100", 930=>x"5a00", 931=>x"2a00", 932=>x"8a00",
---- 933=>x"8000", 934=>x"9600", 935=>x"5400", 936=>x"6600",
---- 937=>x"7600", 938=>x"8900", 939=>x"9600", 940=>x"9c00",
---- 941=>x"7400", 942=>x"7900", 943=>x"8500", 944=>x"5e00",
---- 945=>x"6c00", 946=>x"8600", 947=>x"8f00", 948=>x"3000",
---- 949=>x"5200", 950=>x"7000", 951=>x"9d00", 952=>x"2c00",
---- 953=>x"2700", 954=>x"4d00", 955=>x"7d00", 956=>x"2e00",
---- 957=>x"2b00", 958=>x"3900", 959=>x"5200", 960=>x"3600",
---- 961=>x"4100", 962=>x"3c00", 963=>x"4300", 964=>x"3000",
---- 965=>x"4c00", 966=>x"5600", 967=>x"3500", 968=>x"3200",
---- 969=>x"4000", 970=>x"6700", 971=>x"3f00", 972=>x"3300",
---- 973=>x"4300", 974=>x"3e00", 975=>x"5200", 976=>x"4800",
---- 977=>x"3800", 978=>x"3b00", 979=>x"4b00", 980=>x"7b00",
---- 981=>x"3500", 982=>x"3700", 983=>x"3a00", 984=>x"6e00",
---- 985=>x"5d00", 986=>x"4000", 987=>x"3800", 988=>x"4600",
---- 989=>x"6a00", 990=>x"4c00", 991=>x"4200", 992=>x"4800",
---- 993=>x"5200", 994=>x"6600", 995=>x"3c00", 996=>x"d200",
---- 997=>x"5200", 998=>x"7200", 999=>x"4a00", 1000=>x"2000",
---- 1001=>x"4400", 1002=>x"5b00", 1003=>x"7c00", 1004=>x"1e00",
---- 1005=>x"3800", 1006=>x"4900", 1007=>x"6900", 1008=>x"3d00",
---- 1009=>x"2a00", 1010=>x"4e00", 1011=>x"4600", 1012=>x"4000",
---- 1013=>x"3a00", 1014=>x"4500", 1015=>x"5600", 1016=>x"2500",
---- 1017=>x"3000", 1018=>x"3f00", 1019=>x"5800", 1020=>x"2d00",
---- 1021=>x"2e00", 1022=>x"3000", 1023=>x"4200"),
----
---- 19 => (0=>x"8300", 1=>x"8100", 2=>x"8500", 3=>x"8700", 4=>x"8200",
---- 5=>x"8000", 6=>x"8600", 7=>x"8700", 8=>x"8100",
---- 9=>x"8100", 10=>x"8600", 11=>x"8700", 12=>x"8000",
---- 13=>x"8400", 14=>x"8300", 15=>x"8300", 16=>x"8200",
---- 17=>x"8200", 18=>x"8200", 19=>x"8300", 20=>x"8200",
---- 21=>x"8200", 22=>x"8000", 23=>x"8300", 24=>x"8300",
---- 25=>x"7d00", 26=>x"8100", 27=>x"8600", 28=>x"8200",
---- 29=>x"8100", 30=>x"8300", 31=>x"8300", 32=>x"8300",
---- 33=>x"8300", 34=>x"8000", 35=>x"8200", 36=>x"8500",
---- 37=>x"8300", 38=>x"8100", 39=>x"8200", 40=>x"8400",
---- 41=>x"8300", 42=>x"8200", 43=>x"8300", 44=>x"8100",
---- 45=>x"8000", 46=>x"8200", 47=>x"8200", 48=>x"8000",
---- 49=>x"8000", 50=>x"8100", 51=>x"8100", 52=>x"8000",
---- 53=>x"8200", 54=>x"8400", 55=>x"8000", 56=>x"8300",
---- 57=>x"8200", 58=>x"8100", 59=>x"8300", 60=>x"8000",
---- 61=>x"8200", 62=>x"8100", 63=>x"8000", 64=>x"7f00",
---- 65=>x"8300", 66=>x"8100", 67=>x"8100", 68=>x"7e00",
---- 69=>x"7f00", 70=>x"8100", 71=>x"8300", 72=>x"7b00",
---- 73=>x"7d00", 74=>x"8100", 75=>x"8100", 76=>x"7e00",
---- 77=>x"7f00", 78=>x"7f00", 79=>x"8000", 80=>x"7d00",
---- 81=>x"7d00", 82=>x"8100", 83=>x"7f00", 84=>x"7f00",
---- 85=>x"7f00", 86=>x"8100", 87=>x"7f00", 88=>x"8000",
---- 89=>x"8200", 90=>x"8300", 91=>x"8000", 92=>x"8000",
---- 93=>x"7f00", 94=>x"8300", 95=>x"8100", 96=>x"7f00",
---- 97=>x"8200", 98=>x"8000", 99=>x"7e00", 100=>x"8100",
---- 101=>x"8200", 102=>x"8200", 103=>x"7c00", 104=>x"8000",
---- 105=>x"8100", 106=>x"8100", 107=>x"7d00", 108=>x"7e00",
---- 109=>x"8000", 110=>x"8300", 111=>x"8100", 112=>x"8000",
---- 113=>x"8100", 114=>x"8000", 115=>x"8000", 116=>x"7f00",
---- 117=>x"8000", 118=>x"8000", 119=>x"8000", 120=>x"7f00",
---- 121=>x"7f00", 122=>x"7b00", 123=>x"7b00", 124=>x"7d00",
---- 125=>x"7f00", 126=>x"7800", 127=>x"8500", 128=>x"7b00",
---- 129=>x"7b00", 130=>x"7b00", 131=>x"a900", 132=>x"7900",
---- 133=>x"7600", 134=>x"9b00", 135=>x"a800", 136=>x"7d00",
---- 137=>x"7500", 138=>x"6400", 139=>x"8e00", 140=>x"7d00",
---- 141=>x"8600", 142=>x"7400", 143=>x"6a00", 144=>x"8100",
---- 145=>x"9100", 146=>x"7000", 147=>x"6f00", 148=>x"ac00",
---- 149=>x"8900", 150=>x"6a00", 151=>x"7300", 152=>x"a500",
---- 153=>x"7400", 154=>x"7200", 155=>x"7300", 156=>x"8400",
---- 157=>x"7000", 158=>x"7300", 159=>x"6b00", 160=>x"7700",
---- 161=>x"7000", 162=>x"6c00", 163=>x"6d00", 164=>x"6d00",
---- 165=>x"6d00", 166=>x"6c00", 167=>x"6e00", 168=>x"6d00",
---- 169=>x"6a00", 170=>x"6f00", 171=>x"6d00", 172=>x"6a00",
---- 173=>x"6c00", 174=>x"6f00", 175=>x"7000", 176=>x"6a00",
---- 177=>x"6b00", 178=>x"6f00", 179=>x"7300", 180=>x"6d00",
---- 181=>x"6d00", 182=>x"6f00", 183=>x"7300", 184=>x"7300",
---- 185=>x"7100", 186=>x"7100", 187=>x"6f00", 188=>x"6f00",
---- 189=>x"6f00", 190=>x"7400", 191=>x"7000", 192=>x"7200",
---- 193=>x"7000", 194=>x"7000", 195=>x"7400", 196=>x"6e00",
---- 197=>x"7000", 198=>x"7100", 199=>x"7400", 200=>x"6d00",
---- 201=>x"6e00", 202=>x"7100", 203=>x"7100", 204=>x"7200",
---- 205=>x"7000", 206=>x"7000", 207=>x"6f00", 208=>x"7300",
---- 209=>x"7100", 210=>x"7100", 211=>x"7500", 212=>x"7300",
---- 213=>x"7000", 214=>x"6e00", 215=>x"6f00", 216=>x"6f00",
---- 217=>x"7100", 218=>x"7100", 219=>x"7200", 220=>x"6c00",
---- 221=>x"7000", 222=>x"7300", 223=>x"7100", 224=>x"6e00",
---- 225=>x"8e00", 226=>x"7200", 227=>x"7200", 228=>x"7300",
---- 229=>x"7100", 230=>x"6c00", 231=>x"6b00", 232=>x"6f00",
---- 233=>x"6e00", 234=>x"7400", 235=>x"6c00", 236=>x"7000",
---- 237=>x"7100", 238=>x"7500", 239=>x"7500", 240=>x"7300",
---- 241=>x"7400", 242=>x"7300", 243=>x"7800", 244=>x"6e00",
---- 245=>x"7000", 246=>x"7400", 247=>x"7300", 248=>x"7000",
---- 249=>x"6800", 250=>x"7900", 251=>x"7200", 252=>x"6000",
---- 253=>x"6f00", 254=>x"7500", 255=>x"6f00", 256=>x"6d00",
---- 257=>x"7700", 258=>x"7700", 259=>x"7800", 260=>x"7500",
---- 261=>x"7200", 262=>x"7500", 263=>x"8200", 264=>x"7200",
---- 265=>x"7800", 266=>x"7500", 267=>x"7500", 268=>x"7300",
---- 269=>x"6f00", 270=>x"6800", 271=>x"7600", 272=>x"6c00",
---- 273=>x"6200", 274=>x"7200", 275=>x"7800", 276=>x"6600",
---- 277=>x"7400", 278=>x"7700", 279=>x"7700", 280=>x"6900",
---- 281=>x"6b00", 282=>x"7200", 283=>x"6700", 284=>x"6800",
---- 285=>x"7000", 286=>x"6a00", 287=>x"6c00", 288=>x"6a00",
---- 289=>x"6b00", 290=>x"7200", 291=>x"7000", 292=>x"6c00",
---- 293=>x"7200", 294=>x"7500", 295=>x"7000", 296=>x"6f00",
---- 297=>x"7200", 298=>x"7900", 299=>x"7700", 300=>x"6f00",
---- 301=>x"7300", 302=>x"6400", 303=>x"6c00", 304=>x"6d00",
---- 305=>x"6600", 306=>x"6300", 307=>x"7400", 308=>x"6800",
---- 309=>x"7400", 310=>x"6e00", 311=>x"7200", 312=>x"7000",
---- 313=>x"6b00", 314=>x"6e00", 315=>x"7b00", 316=>x"6100",
---- 317=>x"6900", 318=>x"7700", 319=>x"7400", 320=>x"5c00",
---- 321=>x"6f00", 322=>x"6f00", 323=>x"6d00", 324=>x"6e00",
---- 325=>x"6c00", 326=>x"6c00", 327=>x"6100", 328=>x"6b00",
---- 329=>x"6d00", 330=>x"6400", 331=>x"7c00", 332=>x"6700",
---- 333=>x"5e00", 334=>x"7600", 335=>x"8600", 336=>x"a400",
---- 337=>x"7300", 338=>x"8d00", 339=>x"8800", 340=>x"6500",
---- 341=>x"8600", 342=>x"8a00", 343=>x"8b00", 344=>x"7800",
---- 345=>x"8300", 346=>x"8100", 347=>x"8200", 348=>x"7a00",
---- 349=>x"7e00", 350=>x"7c00", 351=>x"7d00", 352=>x"7a00",
---- 353=>x"7600", 354=>x"7400", 355=>x"7c00", 356=>x"7300",
---- 357=>x"7c00", 358=>x"7200", 359=>x"7a00", 360=>x"7100",
---- 361=>x"7c00", 362=>x"7c00", 363=>x"8000", 364=>x"6f00",
---- 365=>x"7100", 366=>x"8400", 367=>x"7100", 368=>x"7400",
---- 369=>x"7600", 370=>x"7600", 371=>x"6700", 372=>x"8000",
---- 373=>x"6f00", 374=>x"6100", 375=>x"6f00", 376=>x"7200",
---- 377=>x"6600", 378=>x"6b00", 379=>x"7200", 380=>x"6400",
---- 381=>x"6900", 382=>x"7000", 383=>x"7500", 384=>x"6300",
---- 385=>x"7600", 386=>x"7700", 387=>x"8400", 388=>x"6d00",
---- 389=>x"8c00", 390=>x"8400", 391=>x"8b00", 392=>x"7a00",
---- 393=>x"7e00", 394=>x"8900", 395=>x"8500", 396=>x"8000",
---- 397=>x"8100", 398=>x"8b00", 399=>x"8800", 400=>x"8300",
---- 401=>x"7900", 402=>x"7f00", 403=>x"8a00", 404=>x"8200",
---- 405=>x"8300", 406=>x"7c00", 407=>x"8000", 408=>x"8100",
---- 409=>x"8400", 410=>x"8000", 411=>x"7400", 412=>x"8200",
---- 413=>x"8400", 414=>x"7d00", 415=>x"7400", 416=>x"7a00",
---- 417=>x"7d00", 418=>x"7100", 419=>x"7500", 420=>x"7600",
---- 421=>x"7000", 422=>x"6600", 423=>x"7600", 424=>x"7200",
---- 425=>x"6300", 426=>x"6d00", 427=>x"7900", 428=>x"7500",
---- 429=>x"9600", 430=>x"7700", 431=>x"7c00", 432=>x"7400",
---- 433=>x"7b00", 434=>x"7e00", 435=>x"7a00", 436=>x"7700",
---- 437=>x"7b00", 438=>x"7d00", 439=>x"7100", 440=>x"7500",
---- 441=>x"7800", 442=>x"7100", 443=>x"6c00", 444=>x"7200",
---- 445=>x"7500", 446=>x"6e00", 447=>x"7b00", 448=>x"6b00",
---- 449=>x"6800", 450=>x"8000", 451=>x"8800", 452=>x"6400",
---- 453=>x"7a00", 454=>x"8800", 455=>x"7e00", 456=>x"7800",
---- 457=>x"7e00", 458=>x"7f00", 459=>x"7d00", 460=>x"8200",
---- 461=>x"7900", 462=>x"7600", 463=>x"8500", 464=>x"7900",
---- 465=>x"8400", 466=>x"8400", 467=>x"7d00", 468=>x"8100",
---- 469=>x"8200", 470=>x"8800", 471=>x"8300", 472=>x"8a00",
---- 473=>x"7f00", 474=>x"7e00", 475=>x"7d00", 476=>x"7d00",
---- 477=>x"7f00", 478=>x"7c00", 479=>x"6700", 480=>x"7d00",
---- 481=>x"7400", 482=>x"7c00", 483=>x"7100", 484=>x"7800",
---- 485=>x"7600", 486=>x"8100", 487=>x"5700", 488=>x"7000",
---- 489=>x"7a00", 490=>x"7000", 491=>x"3800", 492=>x"6700",
---- 493=>x"6600", 494=>x"3b00", 495=>x"3300", 496=>x"4a00",
---- 497=>x"5200", 498=>x"3600", 499=>x"3a00", 500=>x"4a00",
---- 501=>x"5400", 502=>x"3600", 503=>x"4800", 504=>x"4600",
---- 505=>x"4000", 506=>x"3c00", 507=>x"5f00", 508=>x"2f00",
---- 509=>x"3600", 510=>x"4700", 511=>x"6e00", 512=>x"3400",
---- 513=>x"4d00", 514=>x"6500", 515=>x"6e00", 516=>x"5000",
---- 517=>x"5b00", 518=>x"8400", 519=>x"5100", 520=>x"4700",
---- 521=>x"7400", 522=>x"6700", 523=>x"5700", 524=>x"5800",
---- 525=>x"6100", 526=>x"3100", 527=>x"4f00", 528=>x"6a00",
---- 529=>x"2a00", 530=>x"2200", 531=>x"4100", 532=>x"4000",
---- 533=>x"d700", 534=>x"2900", 535=>x"4800", 536=>x"4700",
---- 537=>x"3800", 538=>x"2b00", 539=>x"4b00", 540=>x"4600",
---- 541=>x"4400", 542=>x"3c00", 543=>x"5e00", 544=>x"b000",
---- 545=>x"5a00", 546=>x"5000", 547=>x"6300", 548=>x"5800",
---- 549=>x"4e00", 550=>x"4b00", 551=>x"6800", 552=>x"5500",
---- 553=>x"4700", 554=>x"5100", 555=>x"6600", 556=>x"6500",
---- 557=>x"3700", 558=>x"4000", 559=>x"6800", 560=>x"6900",
---- 561=>x"4900", 562=>x"3600", 563=>x"6b00", 564=>x"5e00",
---- 565=>x"6e00", 566=>x"5100", 567=>x"5700", 568=>x"3700",
---- 569=>x"7000", 570=>x"7800", 571=>x"5600", 572=>x"3300",
---- 573=>x"3400", 574=>x"7900", 575=>x"9700", 576=>x"5900",
---- 577=>x"3c00", 578=>x"4900", 579=>x"6200", 580=>x"6b00",
---- 581=>x"6600", 582=>x"6900", 583=>x"5500", 584=>x"5300",
---- 585=>x"5300", 586=>x"7900", 587=>x"8300", 588=>x"4300",
---- 589=>x"5100", 590=>x"4200", 591=>x"4b00", 592=>x"2c00",
---- 593=>x"4900", 594=>x"5100", 595=>x"3100", 596=>x"2e00",
---- 597=>x"3900", 598=>x"3c00", 599=>x"3900", 600=>x"3200",
---- 601=>x"3a00", 602=>x"2e00", 603=>x"2b00", 604=>x"2f00",
---- 605=>x"3000", 606=>x"5600", 607=>x"3b00", 608=>x"2900",
---- 609=>x"2f00", 610=>x"5400", 611=>x"3b00", 612=>x"2b00",
---- 613=>x"3100", 614=>x"4b00", 615=>x"4900", 616=>x"3200",
---- 617=>x"4a00", 618=>x"6f00", 619=>x"5c00", 620=>x"3700",
---- 621=>x"4000", 622=>x"7100", 623=>x"6d00", 624=>x"3e00",
---- 625=>x"af00", 626=>x"5000", 627=>x"5e00", 628=>x"3500",
---- 629=>x"5d00", 630=>x"4100", 631=>x"4700", 632=>x"3c00",
---- 633=>x"4800", 634=>x"4f00", 635=>x"6c00", 636=>x"3e00",
---- 637=>x"4c00", 638=>x"8200", 639=>x"8500", 640=>x"2e00",
---- 641=>x"4400", 642=>x"4000", 643=>x"3000", 644=>x"2c00",
---- 645=>x"3600", 646=>x"3e00", 647=>x"3800", 648=>x"2200",
---- 649=>x"2100", 650=>x"2900", 651=>x"4700", 652=>x"2600",
---- 653=>x"2800", 654=>x"2200", 655=>x"2400", 656=>x"3200",
---- 657=>x"1f00", 658=>x"2300", 659=>x"2100", 660=>x"4100",
---- 661=>x"1900", 662=>x"1a00", 663=>x"4500", 664=>x"4400",
---- 665=>x"2500", 666=>x"3200", 667=>x"4d00", 668=>x"3c00",
---- 669=>x"3e00", 670=>x"4600", 671=>x"2b00", 672=>x"3c00",
---- 673=>x"3400", 674=>x"3d00", 675=>x"2300", 676=>x"3000",
---- 677=>x"1f00", 678=>x"3600", 679=>x"4100", 680=>x"3700",
---- 681=>x"3a00", 682=>x"4500", 683=>x"6400", 684=>x"2f00",
---- 685=>x"6d00", 686=>x"7200", 687=>x"6200", 688=>x"6a00",
---- 689=>x"8b00", 690=>x"9e00", 691=>x"9800", 692=>x"6f00",
---- 693=>x"7400", 694=>x"a200", 695=>x"c600", 696=>x"8800",
---- 697=>x"6c00", 698=>x"9f00", 699=>x"c200", 700=>x"8100",
---- 701=>x"8900", 702=>x"b800", 703=>x"bf00", 704=>x"7f00",
---- 705=>x"8900", 706=>x"bb00", 707=>x"2400", 708=>x"8900",
---- 709=>x"8400", 710=>x"9800", 711=>x"e200", 712=>x"8700",
---- 713=>x"7a00", 714=>x"7d00", 715=>x"d100", 716=>x"8000",
---- 717=>x"7800", 718=>x"a100", 719=>x"cd00", 720=>x"7500",
---- 721=>x"8300", 722=>x"d400", 723=>x"ac00", 724=>x"7300",
---- 725=>x"8300", 726=>x"c900", 727=>x"9200", 728=>x"7e00",
---- 729=>x"8a00", 730=>x"ca00", 731=>x"a600", 732=>x"7b00",
---- 733=>x"9f00", 734=>x"c900", 735=>x"9600", 736=>x"7100",
---- 737=>x"9b00", 738=>x"c900", 739=>x"a300", 740=>x"8000",
---- 741=>x"af00", 742=>x"da00", 743=>x"cc00", 744=>x"7300",
---- 745=>x"a000", 746=>x"d700", 747=>x"c200", 748=>x"6f00",
---- 749=>x"7600", 750=>x"c100", 751=>x"7d00", 752=>x"6800",
---- 753=>x"7900", 754=>x"b700", 755=>x"6500", 756=>x"5b00",
---- 757=>x"6200", 758=>x"5700", 759=>x"4700", 760=>x"6100",
---- 761=>x"6c00", 762=>x"3700", 763=>x"3f00", 764=>x"4800",
---- 765=>x"6200", 766=>x"5b00", 767=>x"3e00", 768=>x"7300",
---- 769=>x"7b00", 770=>x"7d00", 771=>x"4b00", 772=>x"9800",
---- 773=>x"a700", 774=>x"9b00", 775=>x"7f00", 776=>x"5100",
---- 777=>x"7600", 778=>x"9600", 779=>x"a600", 780=>x"5500",
---- 781=>x"3600", 782=>x"4900", 783=>x"9c00", 784=>x"7a00",
---- 785=>x"6500", 786=>x"3100", 787=>x"6300", 788=>x"6000",
---- 789=>x"6600", 790=>x"4a00", 791=>x"4900", 792=>x"7800",
---- 793=>x"3e00", 794=>x"6400", 795=>x"7f00", 796=>x"7300",
---- 797=>x"6000", 798=>x"6e00", 799=>x"9800", 800=>x"6f00",
---- 801=>x"6f00", 802=>x"7100", 803=>x"7600", 804=>x"7e00",
---- 805=>x"8e00", 806=>x"8200", 807=>x"7c00", 808=>x"9c00",
---- 809=>x"7a00", 810=>x"8600", 811=>x"7900", 812=>x"9500",
---- 813=>x"8b00", 814=>x"7f00", 815=>x"8600", 816=>x"8900",
---- 817=>x"8b00", 818=>x"8b00", 819=>x"9200", 820=>x"8700",
---- 821=>x"8100", 822=>x"9600", 823=>x"9500", 824=>x"9000",
---- 825=>x"8100", 826=>x"9000", 827=>x"8200", 828=>x"8f00",
---- 829=>x"8700", 830=>x"8500", 831=>x"7600", 832=>x"9300",
---- 833=>x"8200", 834=>x"8300", 835=>x"8500", 836=>x"7c00",
---- 837=>x"8c00", 838=>x"7300", 839=>x"8e00", 840=>x"6300",
---- 841=>x"6400", 842=>x"7a00", 843=>x"7e00", 844=>x"5d00",
---- 845=>x"6f00", 846=>x"8d00", 847=>x"6b00", 848=>x"5300",
---- 849=>x"6d00", 850=>x"8e00", 851=>x"8300", 852=>x"5100",
---- 853=>x"5c00", 854=>x"8f00", 855=>x"9d00", 856=>x"4f00",
---- 857=>x"5f00", 858=>x"8a00", 859=>x"6a00", 860=>x"4700",
---- 861=>x"6500", 862=>x"8500", 863=>x"9000", 864=>x"3d00",
---- 865=>x"5e00", 866=>x"9500", 867=>x"8700", 868=>x"3700",
---- 869=>x"5500", 870=>x"9900", 871=>x"8900", 872=>x"4e00",
---- 873=>x"6600", 874=>x"8f00", 875=>x"8900", 876=>x"6100",
---- 877=>x"6d00", 878=>x"8b00", 879=>x"8700", 880=>x"7a00",
---- 881=>x"7900", 882=>x"8400", 883=>x"8f00", 884=>x"8b00",
---- 885=>x"8600", 886=>x"7900", 887=>x"8800", 888=>x"9100",
---- 889=>x"8800", 890=>x"7800", 891=>x"8400", 892=>x"8500",
---- 893=>x"6300", 894=>x"8900", 895=>x"7500", 896=>x"7900",
---- 897=>x"6800", 898=>x"7800", 899=>x"7c00", 900=>x"6100",
---- 901=>x"7800", 902=>x"7300", 903=>x"6a00", 904=>x"5300",
---- 905=>x"6600", 906=>x"7300", 907=>x"7400", 908=>x"8300",
---- 909=>x"8100", 910=>x"7700", 911=>x"7c00", 912=>x"6000",
---- 913=>x"7c00", 914=>x"7900", 915=>x"7700", 916=>x"3500",
---- 917=>x"3b00", 918=>x"5b00", 919=>x"8b00", 920=>x"3700",
---- 921=>x"2800", 922=>x"2800", 923=>x"6600", 924=>x"3500",
---- 925=>x"2500", 926=>x"2e00", 927=>x"4100", 928=>x"4300",
---- 929=>x"4700", 930=>x"2d00", 931=>x"3b00", 932=>x"3300",
---- 933=>x"4900", 934=>x"4000", 935=>x"4000", 936=>x"6700",
---- 937=>x"3400", 938=>x"3d00", 939=>x"5b00", 940=>x"9300",
---- 941=>x"6b00", 942=>x"6500", 943=>x"6b00", 944=>x"7100",
---- 945=>x"8500", 946=>x"7b00", 947=>x"6600", 948=>x"8b00",
---- 949=>x"7a00", 950=>x"8200", 951=>x"5400", 952=>x"8900",
---- 953=>x"8d00", 954=>x"8600", 955=>x"6400", 956=>x"7500",
---- 957=>x"7200", 958=>x"a700", 959=>x"8b00", 960=>x"4a00",
---- 961=>x"5400", 962=>x"7600", 963=>x"8a00", 964=>x"4e00",
---- 965=>x"4b00", 966=>x"5c00", 967=>x"5000", 968=>x"4700",
---- 969=>x"7800", 970=>x"8100", 971=>x"4200", 972=>x"4800",
---- 973=>x"6400", 974=>x"9700", 975=>x"6600", 976=>x"5000",
---- 977=>x"4a00", 978=>x"8a00", 979=>x"8200", 980=>x"5400",
---- 981=>x"6600", 982=>x"7400", 983=>x"9d00", 984=>x"4d00",
---- 985=>x"7300", 986=>x"6e00", 987=>x"8500", 988=>x"3d00",
---- 989=>x"7100", 990=>x"7800", 991=>x"6300", 992=>x"4400",
---- 993=>x"5f00", 994=>x"7100", 995=>x"7500", 996=>x"2a00",
---- 997=>x"4c00", 998=>x"6c00", 999=>x"7800", 1000=>x"3300",
---- 1001=>x"2900", 1002=>x"4c00", 1003=>x"5d00", 1004=>x"6b00",
---- 1005=>x"2400", 1006=>x"3c00", 1007=>x"4a00", 1008=>x"6800",
---- 1009=>x"4200", 1010=>x"3800", 1011=>x"4c00", 1012=>x"4400",
---- 1013=>x"4a00", 1014=>x"2e00", 1015=>x"4300", 1016=>x"4900",
---- 1017=>x"3d00", 1018=>x"3300", 1019=>x"2e00", 1020=>x"4e00",
---- 1021=>x"4700", 1022=>x"3f00", 1023=>x"2c00"),
----
---- 20 => (0=>x"8100", 1=>x"8600", 2=>x"8500", 3=>x"8600", 4=>x"8200",
---- 5=>x"8400", 6=>x"8500", 7=>x"8600", 8=>x"8300",
---- 9=>x"7900", 10=>x"8600", 11=>x"8700", 12=>x"8300",
---- 13=>x"8500", 14=>x"8700", 15=>x"8700", 16=>x"8400",
---- 17=>x"8300", 18=>x"8300", 19=>x"8500", 20=>x"8200",
---- 21=>x"8300", 22=>x"7b00", 23=>x"8600", 24=>x"8000",
---- 25=>x"8300", 26=>x"8500", 27=>x"8400", 28=>x"8100",
---- 29=>x"8300", 30=>x"8000", 31=>x"8200", 32=>x"8400",
---- 33=>x"8600", 34=>x"8700", 35=>x"8400", 36=>x"8300",
---- 37=>x"8300", 38=>x"8600", 39=>x"8200", 40=>x"8200",
---- 41=>x"8000", 42=>x"8300", 43=>x"8300", 44=>x"8100",
---- 45=>x"8300", 46=>x"8400", 47=>x"8400", 48=>x"8100",
---- 49=>x"8100", 50=>x"8300", 51=>x"8200", 52=>x"8100",
---- 53=>x"8300", 54=>x"8100", 55=>x"8000", 56=>x"8200",
---- 57=>x"8200", 58=>x"8100", 59=>x"8400", 60=>x"8000",
---- 61=>x"8300", 62=>x"8200", 63=>x"8100", 64=>x"8400",
---- 65=>x"8200", 66=>x"8300", 67=>x"8300", 68=>x"8400",
---- 69=>x"8200", 70=>x"8100", 71=>x"7f00", 72=>x"8000",
---- 73=>x"7d00", 74=>x"8100", 75=>x"7f00", 76=>x"8200",
---- 77=>x"7f00", 78=>x"8200", 79=>x"7f00", 80=>x"8300",
---- 81=>x"8100", 82=>x"8100", 83=>x"8000", 84=>x"8000",
---- 85=>x"7d00", 86=>x"7f00", 87=>x"8000", 88=>x"8000",
---- 89=>x"7f00", 90=>x"7d00", 91=>x"7a00", 92=>x"8200",
---- 93=>x"8000", 94=>x"7d00", 95=>x"7d00", 96=>x"8100",
---- 97=>x"7f00", 98=>x"7e00", 99=>x"8000", 100=>x"8200",
---- 101=>x"7f00", 102=>x"7f00", 103=>x"7f00", 104=>x"8200",
---- 105=>x"8300", 106=>x"8000", 107=>x"7f00", 108=>x"8000",
---- 109=>x"7e00", 110=>x"7f00", 111=>x"7c00", 112=>x"8000",
---- 113=>x"7e00", 114=>x"7c00", 115=>x"7d00", 116=>x"7d00",
---- 117=>x"7a00", 118=>x"7b00", 119=>x"7a00", 120=>x"7900",
---- 121=>x"7d00", 122=>x"a300", 123=>x"9900", 124=>x"8600",
---- 125=>x"8000", 126=>x"8d00", 127=>x"8d00", 128=>x"9000",
---- 129=>x"6f00", 130=>x"7b00", 131=>x"7b00", 132=>x"5b00",
---- 133=>x"6700", 134=>x"7b00", 135=>x"7900", 136=>x"6000",
---- 137=>x"6e00", 138=>x"7600", 139=>x"7600", 140=>x"7300",
---- 141=>x"7000", 142=>x"7400", 143=>x"7700", 144=>x"7200",
---- 145=>x"7500", 146=>x"7600", 147=>x"7400", 148=>x"7500",
---- 149=>x"7000", 150=>x"6f00", 151=>x"6d00", 152=>x"6c00",
---- 153=>x"6e00", 154=>x"6900", 155=>x"6c00", 156=>x"6a00",
---- 157=>x"9400", 158=>x"6c00", 159=>x"7000", 160=>x"6a00",
---- 161=>x"6d00", 162=>x"6f00", 163=>x"7100", 164=>x"7100",
---- 165=>x"7100", 166=>x"7500", 167=>x"7700", 168=>x"6f00",
---- 169=>x"8900", 170=>x"7800", 171=>x"7600", 172=>x"7300",
---- 173=>x"7700", 174=>x"7200", 175=>x"7400", 176=>x"7300",
---- 177=>x"7100", 178=>x"6f00", 179=>x"7a00", 180=>x"6f00",
---- 181=>x"7300", 182=>x"7d00", 183=>x"7500", 184=>x"7200",
---- 185=>x"7900", 186=>x"7800", 187=>x"7600", 188=>x"7700",
---- 189=>x"7500", 190=>x"7300", 191=>x"8700", 192=>x"7800",
---- 193=>x"7500", 194=>x"7700", 195=>x"7000", 196=>x"7400",
---- 197=>x"7600", 198=>x"6f00", 199=>x"7400", 200=>x"7600",
---- 201=>x"7700", 202=>x"7100", 203=>x"7800", 204=>x"7100",
---- 205=>x"7000", 206=>x"7200", 207=>x"7400", 208=>x"7400",
---- 209=>x"7200", 210=>x"8d00", 211=>x"7100", 212=>x"7200",
---- 213=>x"7200", 214=>x"6f00", 215=>x"6f00", 216=>x"6f00",
---- 217=>x"7100", 218=>x"7200", 219=>x"7500", 220=>x"7400",
---- 221=>x"7900", 222=>x"7700", 223=>x"7a00", 224=>x"7600",
---- 225=>x"7800", 226=>x"7b00", 227=>x"7600", 228=>x"6d00",
---- 229=>x"7800", 230=>x"7700", 231=>x"7800", 232=>x"7100",
---- 233=>x"7700", 234=>x"7500", 235=>x"7500", 236=>x"7300",
---- 237=>x"7c00", 238=>x"8900", 239=>x"7500", 240=>x"7600",
---- 241=>x"7800", 242=>x"7700", 243=>x"7900", 244=>x"7800",
---- 245=>x"7000", 246=>x"7600", 247=>x"7e00", 248=>x"7000",
---- 249=>x"7700", 250=>x"8000", 251=>x"8500", 252=>x"7d00",
---- 253=>x"8200", 254=>x"7e00", 255=>x"8200", 256=>x"7b00",
---- 257=>x"7f00", 258=>x"7800", 259=>x"7900", 260=>x"7900",
---- 261=>x"7900", 262=>x"7c00", 263=>x"7a00", 264=>x"7d00",
---- 265=>x"7d00", 266=>x"6d00", 267=>x"7200", 268=>x"7a00",
---- 269=>x"6a00", 270=>x"7400", 271=>x"8000", 272=>x"7200",
---- 273=>x"7500", 274=>x"7a00", 275=>x"7a00", 276=>x"7100",
---- 277=>x"7100", 278=>x"7c00", 279=>x"7d00", 280=>x"6800",
---- 281=>x"7600", 282=>x"7800", 283=>x"7c00", 284=>x"7700",
---- 285=>x"7a00", 286=>x"7c00", 287=>x"7300", 288=>x"7300",
---- 289=>x"7b00", 290=>x"7100", 291=>x"6d00", 292=>x"7800",
---- 293=>x"7400", 294=>x"6f00", 295=>x"7c00", 296=>x"7600",
---- 297=>x"7e00", 298=>x"7a00", 299=>x"7c00", 300=>x"7900",
---- 301=>x"7700", 302=>x"7a00", 303=>x"7d00", 304=>x"7900",
---- 305=>x"7400", 306=>x"7900", 307=>x"7400", 308=>x"8100",
---- 309=>x"7100", 310=>x"6300", 311=>x"6600", 312=>x"7800",
---- 313=>x"6c00", 314=>x"6100", 315=>x"7200", 316=>x"7400",
---- 317=>x"6700", 318=>x"7400", 319=>x"8b00", 320=>x"6000",
---- 321=>x"7800", 322=>x"9200", 323=>x"8b00", 324=>x"6f00",
---- 325=>x"9100", 326=>x"9000", 327=>x"8b00", 328=>x"8f00",
---- 329=>x"9000", 330=>x"8c00", 331=>x"8700", 332=>x"8a00",
---- 333=>x"8e00", 334=>x"8800", 335=>x"8600", 336=>x"7900",
---- 337=>x"8700", 338=>x"8700", 339=>x"7f00", 340=>x"8300",
---- 341=>x"7b00", 342=>x"8400", 343=>x"8900", 344=>x"8500",
---- 345=>x"7c00", 346=>x"8800", 347=>x"8d00", 348=>x"7d00",
---- 349=>x"8800", 350=>x"8700", 351=>x"7200", 352=>x"7f00",
---- 353=>x"8900", 354=>x"7000", 355=>x"6f00", 356=>x"8600",
---- 357=>x"6e00", 358=>x"6800", 359=>x"7800", 360=>x"6d00",
---- 361=>x"6200", 362=>x"7700", 363=>x"8500", 364=>x"6300",
---- 365=>x"7100", 366=>x"7700", 367=>x"8800", 368=>x"7300",
---- 369=>x"7700", 370=>x"8300", 371=>x"8c00", 372=>x"7400",
---- 373=>x"8000", 374=>x"8800", 375=>x"8b00", 376=>x"7e00",
---- 377=>x"8600", 378=>x"8900", 379=>x"8500", 380=>x"8900",
---- 381=>x"8400", 382=>x"8500", 383=>x"8900", 384=>x"8700",
---- 385=>x"8800", 386=>x"8500", 387=>x"8900", 388=>x"8700",
---- 389=>x"8600", 390=>x"8500", 391=>x"7900", 392=>x"8800",
---- 393=>x"8700", 394=>x"7200", 395=>x"6000", 396=>x"8600",
---- 397=>x"8300", 398=>x"6b00", 399=>x"7400", 400=>x"7c00",
---- 401=>x"6900", 402=>x"7300", 403=>x"8200", 404=>x"7200",
---- 405=>x"6900", 406=>x"7c00", 407=>x"7f00", 408=>x"6d00",
---- 409=>x"7900", 410=>x"7f00", 411=>x"8500", 412=>x"7500",
---- 413=>x"7c00", 414=>x"8200", 415=>x"8000", 416=>x"8100",
---- 417=>x"7e00", 418=>x"8500", 419=>x"7e00", 420=>x"7f00",
---- 421=>x"8100", 422=>x"8300", 423=>x"7600", 424=>x"8000",
---- 425=>x"8100", 426=>x"7800", 427=>x"7000", 428=>x"7b00",
---- 429=>x"7500", 430=>x"7000", 431=>x"7c00", 432=>x"6a00",
---- 433=>x"6b00", 434=>x"7b00", 435=>x"8600", 436=>x"6700",
---- 437=>x"7400", 438=>x"8800", 439=>x"8900", 440=>x"7800",
---- 441=>x"8100", 442=>x"7e00", 443=>x"8500", 444=>x"8000",
---- 445=>x"8200", 446=>x"8300", 447=>x"6d00", 448=>x"7800",
---- 449=>x"7900", 450=>x"7d00", 451=>x"6500", 452=>x"8300",
---- 453=>x"7900", 454=>x"5c00", 455=>x"5d00", 456=>x"8500",
---- 457=>x"8900", 458=>x"7900", 459=>x"7000", 460=>x"8300",
---- 461=>x"8000", 462=>x"6d00", 463=>x"6700", 464=>x"8100",
---- 465=>x"6900", 466=>x"6200", 467=>x"5a00", 468=>x"7900",
---- 469=>x"6200", 470=>x"4400", 471=>x"3100", 472=>x"6300",
---- 473=>x"4600", 474=>x"2e00", 475=>x"4300", 476=>x"5500",
---- 477=>x"3100", 478=>x"3800", 479=>x"5200", 480=>x"5000",
---- 481=>x"2c00", 482=>x"5700", 483=>x"5300", 484=>x"2d00",
---- 485=>x"3800", 486=>x"6400", 487=>x"4900", 488=>x"3700",
---- 489=>x"5200", 490=>x"6400", 491=>x"3100", 492=>x"5000",
---- 493=>x"5b00", 494=>x"5700", 495=>x"2400", 496=>x"5200",
---- 497=>x"7000", 498=>x"4100", 499=>x"2500", 500=>x"5e00",
---- 501=>x"5300", 502=>x"d600", 503=>x"2b00", 504=>x"5800",
---- 505=>x"3000", 506=>x"2b00", 507=>x"3e00", 508=>x"5f00",
---- 509=>x"3d00", 510=>x"3f00", 511=>x"6200", 512=>x"3700",
---- 513=>x"4f00", 514=>x"4d00", 515=>x"6400", 516=>x"3100",
---- 517=>x"5700", 518=>x"5200", 519=>x"6800", 520=>x"4800",
---- 521=>x"5b00", 522=>x"4f00", 523=>x"7b00", 524=>x"5800",
---- 525=>x"4f00", 526=>x"5b00", 527=>x"8f00", 528=>x"6b00",
---- 529=>x"6100", 530=>x"6800", 531=>x"7400", 532=>x"7700",
---- 533=>x"5b00", 534=>x"6300", 535=>x"6600", 536=>x"7700",
---- 537=>x"4f00", 538=>x"7300", 539=>x"7000", 540=>x"8300",
---- 541=>x"5b00", 542=>x"7c00", 543=>x"7600", 544=>x"7700",
---- 545=>x"4d00", 546=>x"7300", 547=>x"8000", 548=>x"8200",
---- 549=>x"4200", 550=>x"7700", 551=>x"8a00", 552=>x"8c00",
---- 553=>x"5900", 554=>x"8500", 555=>x"8400", 556=>x"7a00",
---- 557=>x"6b00", 558=>x"8200", 559=>x"6a00", 560=>x"6500",
---- 561=>x"7900", 562=>x"7f00", 563=>x"7600", 564=>x"4700",
---- 565=>x"6d00", 566=>x"7700", 567=>x"8900", 568=>x"5d00",
---- 569=>x"6400", 570=>x"5800", 571=>x"7700", 572=>x"8300",
---- 573=>x"5200", 574=>x"4800", 575=>x"5400", 576=>x"7a00",
---- 577=>x"5400", 578=>x"5800", 579=>x"8500", 580=>x"a600",
---- 581=>x"8100", 582=>x"a000", 583=>x"9200", 584=>x"7900",
---- 585=>x"6000", 586=>x"4d00", 587=>x"3500", 588=>x"6d00",
---- 589=>x"3800", 590=>x"1a00", 591=>x"2500", 592=>x"4e00",
---- 593=>x"3300", 594=>x"2300", 595=>x"2400", 596=>x"4c00",
---- 597=>x"c200", 598=>x"2100", 599=>x"2200", 600=>x"4400",
---- 601=>x"4100", 602=>x"1d00", 603=>x"3200", 604=>x"2700",
---- 605=>x"3e00", 606=>x"2a00", 607=>x"2a00", 608=>x"2d00",
---- 609=>x"3b00", 610=>x"2d00", 611=>x"2f00", 612=>x"4d00",
---- 613=>x"3900", 614=>x"3900", 615=>x"4f00", 616=>x"4e00",
---- 617=>x"3100", 618=>x"4900", 619=>x"5c00", 620=>x"3d00",
---- 621=>x"3a00", 622=>x"5000", 623=>x"7400", 624=>x"3e00",
---- 625=>x"6c00", 626=>x"8500", 627=>x"7400", 628=>x"5400",
---- 629=>x"8b00", 630=>x"7b00", 631=>x"5b00", 632=>x"5600",
---- 633=>x"9200", 634=>x"9200", 635=>x"7300", 636=>x"3e00",
---- 637=>x"3f00", 638=>x"6700", 639=>x"7e00", 640=>x"2800",
---- 641=>x"2800", 642=>x"4200", 643=>x"7400", 644=>x"2800",
---- 645=>x"5400", 646=>x"8800", 647=>x"4c00", 648=>x"4300",
---- 649=>x"7200", 650=>x"a700", 651=>x"3d00", 652=>x"5200",
---- 653=>x"7e00", 654=>x"5500", 655=>x"2b00", 656=>x"6700",
---- 657=>x"6c00", 658=>x"3600", 659=>x"1d00", 660=>x"5d00",
---- 661=>x"3d00", 662=>x"4600", 663=>x"3600", 664=>x"2e00",
---- 665=>x"3b00", 666=>x"5e00", 667=>x"6b00", 668=>x"2500",
---- 669=>x"3c00", 670=>x"7e00", 671=>x"8400", 672=>x"2e00",
---- 673=>x"7900", 674=>x"a200", 675=>x"8e00", 676=>x"5600",
---- 677=>x"9200", 678=>x"9d00", 679=>x"9600", 680=>x"9500",
---- 681=>x"7400", 682=>x"8e00", 683=>x"6100", 684=>x"6100",
---- 685=>x"7c00", 686=>x"9700", 687=>x"a000", 688=>x"8400",
---- 689=>x"8f00", 690=>x"b400", 691=>x"b900", 692=>x"c200",
---- 693=>x"c100", 694=>x"cb00", 695=>x"c500", 696=>x"2e00",
---- 697=>x"cf00", 698=>x"cc00", 699=>x"9200", 700=>x"ce00",
---- 701=>x"d100", 702=>x"ac00", 703=>x"5900", 704=>x"d600",
---- 705=>x"cc00", 706=>x"8000", 707=>x"5a00", 708=>x"d600",
---- 709=>x"a200", 710=>x"6300", 711=>x"6600", 712=>x"bb00",
---- 713=>x"6d00", 714=>x"6300", 715=>x"6f00", 716=>x"7600",
---- 717=>x"6000", 718=>x"7800", 719=>x"9800", 720=>x"5900",
---- 721=>x"8100", 722=>x"9b00", 723=>x"bf00", 724=>x"7900",
---- 725=>x"9e00", 726=>x"b900", 727=>x"ba00", 728=>x"a000",
---- 729=>x"b000", 730=>x"cf00", 731=>x"6a00", 732=>x"a300",
---- 733=>x"c500", 734=>x"8900", 735=>x"2c00", 736=>x"c800",
---- 737=>x"a100", 738=>x"3200", 739=>x"3200", 740=>x"be00",
---- 741=>x"5100", 742=>x"2c00", 743=>x"2d00", 744=>x"5d00",
---- 745=>x"2e00", 746=>x"3200", 747=>x"3200", 748=>x"2600",
---- 749=>x"3b00", 750=>x"3000", 751=>x"3000", 752=>x"3900",
---- 753=>x"4500", 754=>x"2c00", 755=>x"3200", 756=>x"5200",
---- 757=>x"3900", 758=>x"3200", 759=>x"3500", 760=>x"3f00",
---- 761=>x"3500", 762=>x"3100", 763=>x"3200", 764=>x"3400",
---- 765=>x"3800", 766=>x"3300", 767=>x"3200", 768=>x"2e00",
---- 769=>x"2e00", 770=>x"2f00", 771=>x"3400", 772=>x"3600",
---- 773=>x"2e00", 774=>x"2f00", 775=>x"3200", 776=>x"6e00",
---- 777=>x"4100", 778=>x"2d00", 779=>x"2c00", 780=>x"ae00",
---- 781=>x"9000", 782=>x"4400", 783=>x"2300", 784=>x"ae00",
---- 785=>x"ae00", 786=>x"9100", 787=>x"4300", 788=>x"8b00",
---- 789=>x"8800", 790=>x"9b00", 791=>x"9600", 792=>x"9700",
---- 793=>x"7a00", 794=>x"5b00", 795=>x"9b00", 796=>x"b300",
---- 797=>x"7e00", 798=>x"5300", 799=>x"4e00", 800=>x"a700",
---- 801=>x"5f00", 802=>x"5100", 803=>x"4600", 804=>x"8600",
---- 805=>x"9700", 806=>x"5600", 807=>x"3000", 808=>x"5d00",
---- 809=>x"8700", 810=>x"8e00", 811=>x"3500", 812=>x"5100",
---- 813=>x"3c00", 814=>x"7700", 815=>x"7800", 816=>x"6c00",
---- 817=>x"1d00", 818=>x"3e00", 819=>x"ab00", 820=>x"9600",
---- 821=>x"3600", 822=>x"2000", 823=>x"8500", 824=>x"8400",
---- 825=>x"7000", 826=>x"3500", 827=>x"5300", 828=>x"6d00",
---- 829=>x"8d00", 830=>x"6e00", 831=>x"6400", 832=>x"7a00",
---- 833=>x"9300", 834=>x"6600", 835=>x"6a00", 836=>x"8500",
---- 837=>x"a200", 838=>x"8e00", 839=>x"7d00", 840=>x"7f00",
---- 841=>x"a900", 842=>x"a500", 843=>x"7700", 844=>x"7c00",
---- 845=>x"9f00", 846=>x"a700", 847=>x"7700", 848=>x"8a00",
---- 849=>x"9400", 850=>x"8e00", 851=>x"4500", 852=>x"8d00",
---- 853=>x"9400", 854=>x"9300", 855=>x"4300", 856=>x"9000",
---- 857=>x"8900", 858=>x"a600", 859=>x"6400", 860=>x"7300",
---- 861=>x"8b00", 862=>x"9b00", 863=>x"6f00", 864=>x"7100",
---- 865=>x"9800", 866=>x"8c00", 867=>x"8000", 868=>x"8a00",
---- 869=>x"9d00", 870=>x"6900", 871=>x"5300", 872=>x"9200",
---- 873=>x"a400", 874=>x"8f00", 875=>x"5300", 876=>x"9200",
---- 877=>x"7a00", 878=>x"8600", 879=>x"8a00", 880=>x"8c00",
---- 881=>x"4b00", 882=>x"5700", 883=>x"8a00", 884=>x"8400",
---- 885=>x"6e00", 886=>x"5a00", 887=>x"5a00", 888=>x"8300",
---- 889=>x"6900", 890=>x"6100", 891=>x"2c00", 892=>x"6c00",
---- 893=>x"8000", 894=>x"6700", 895=>x"4e00", 896=>x"6500",
---- 897=>x"7b00", 898=>x"8400", 899=>x"7c00", 900=>x"6900",
---- 901=>x"6c00", 902=>x"8700", 903=>x"9500", 904=>x"5900",
---- 905=>x"4300", 906=>x"5e00", 907=>x"7f00", 908=>x"6600",
---- 909=>x"4c00", 910=>x"3a00", 911=>x"6900", 912=>x"5200",
---- 913=>x"3f00", 914=>x"3500", 915=>x"5a00", 916=>x"6d00",
---- 917=>x"3800", 918=>x"2f00", 919=>x"3f00", 920=>x"9400",
---- 921=>x"3d00", 922=>x"3300", 923=>x"5700", 924=>x"6200",
---- 925=>x"4600", 926=>x"2b00", 927=>x"5c00", 928=>x"3500",
---- 929=>x"3300", 930=>x"d100", 931=>x"5f00", 932=>x"4900",
---- 933=>x"4300", 934=>x"4800", 935=>x"8f00", 936=>x"6a00",
---- 937=>x"7700", 938=>x"b500", 939=>x"5300", 940=>x"5e00",
---- 941=>x"7300", 942=>x"5c00", 943=>x"2f00", 944=>x"5800",
---- 945=>x"4700", 946=>x"6300", 947=>x"5600", 948=>x"5b00",
---- 949=>x"6e00", 950=>x"8800", 951=>x"5c00", 952=>x"6800",
---- 953=>x"6700", 954=>x"6600", 955=>x"7c00", 956=>x"6200",
---- 957=>x"5700", 958=>x"7000", 959=>x"8300", 960=>x"7a00",
---- 961=>x"6300", 962=>x"6100", 963=>x"4500", 964=>x"7c00",
---- 965=>x"9400", 966=>x"5e00", 967=>x"2600", 968=>x"4b00",
---- 969=>x"6300", 970=>x"6c00", 971=>x"3a00", 972=>x"4800",
---- 973=>x"2800", 974=>x"5000", 975=>x"4d00", 976=>x"4a00",
---- 977=>x"3700", 978=>x"4500", 979=>x"4a00", 980=>x"7700",
---- 981=>x"3800", 982=>x"3600", 983=>x"c400", 984=>x"6400",
---- 985=>x"5f00", 986=>x"3300", 987=>x"3500", 988=>x"5f00",
---- 989=>x"7900", 990=>x"5a00", 991=>x"3300", 992=>x"4500",
---- 993=>x"6200", 994=>x"6800", 995=>x"3e00", 996=>x"6f00",
---- 997=>x"5100", 998=>x"4b00", 999=>x"4100", 1000=>x"7200",
---- 1001=>x"5200", 1002=>x"2a00", 1003=>x"3700", 1004=>x"6b00",
---- 1005=>x"6900", 1006=>x"4000", 1007=>x"3c00", 1008=>x"5d00",
---- 1009=>x"6500", 1010=>x"5f00", 1011=>x"7100", 1012=>x"5900",
---- 1013=>x"6c00", 1014=>x"4f00", 1015=>x"7800", 1016=>x"3b00",
---- 1017=>x"5700", 1018=>x"4a00", 1019=>x"5300", 1020=>x"2f00",
---- 1021=>x"5400", 1022=>x"5a00", 1023=>x"2e00"),
----
---- 21 => (0=>x"8600", 1=>x"8500", 2=>x"8600", 3=>x"8600", 4=>x"8500",
---- 5=>x"8600", 6=>x"8600", 7=>x"8400", 8=>x"8600",
---- 9=>x"8400", 10=>x"8600", 11=>x"8500", 12=>x"8500",
---- 13=>x"8400", 14=>x"8500", 15=>x"7800", 16=>x"8500",
---- 17=>x"8500", 18=>x"8600", 19=>x"8500", 20=>x"8400",
---- 21=>x"8400", 22=>x"8500", 23=>x"8500", 24=>x"8400",
---- 25=>x"8300", 26=>x"8400", 27=>x"8400", 28=>x"8100",
---- 29=>x"8500", 30=>x"8600", 31=>x"8500", 32=>x"8300",
---- 33=>x"8700", 34=>x"8400", 35=>x"8600", 36=>x"8300",
---- 37=>x"8400", 38=>x"8600", 39=>x"8500", 40=>x"8300",
---- 41=>x"8100", 42=>x"8400", 43=>x"8400", 44=>x"8100",
---- 45=>x"8300", 46=>x"8300", 47=>x"8400", 48=>x"8000",
---- 49=>x"8300", 50=>x"8600", 51=>x"8500", 52=>x"7e00",
---- 53=>x"8100", 54=>x"8000", 55=>x"8200", 56=>x"8100",
---- 57=>x"8100", 58=>x"8000", 59=>x"8400", 60=>x"8200",
---- 61=>x"8200", 62=>x"8000", 63=>x"8300", 64=>x"8300",
---- 65=>x"7d00", 66=>x"8300", 67=>x"8200", 68=>x"8100",
---- 69=>x"8300", 70=>x"8400", 71=>x"7f00", 72=>x"8000",
---- 73=>x"7f00", 74=>x"7e00", 75=>x"8000", 76=>x"7c00",
---- 77=>x"7d00", 78=>x"8000", 79=>x"8000", 80=>x"7e00",
---- 81=>x"8100", 82=>x"8200", 83=>x"8000", 84=>x"7c00",
---- 85=>x"8100", 86=>x"8000", 87=>x"7f00", 88=>x"7e00",
---- 89=>x"8100", 90=>x"8100", 91=>x"8000", 92=>x"7f00",
---- 93=>x"8900", 94=>x"8500", 95=>x"8000", 96=>x"7f00",
---- 97=>x"7f00", 98=>x"8000", 99=>x"8200", 100=>x"7f00",
---- 101=>x"7f00", 102=>x"8100", 103=>x"8200", 104=>x"8000",
---- 105=>x"8100", 106=>x"7f00", 107=>x"8000", 108=>x"7e00",
---- 109=>x"7f00", 110=>x"7f00", 111=>x"7f00", 112=>x"7c00",
---- 113=>x"7d00", 114=>x"8000", 115=>x"8200", 116=>x"7e00",
---- 117=>x"9100", 118=>x"9100", 119=>x"9400", 120=>x"9300",
---- 121=>x"9f00", 122=>x"9400", 123=>x"8e00", 124=>x"8d00",
---- 125=>x"8500", 126=>x"8200", 127=>x"7b00", 128=>x"7e00",
---- 129=>x"7c00", 130=>x"7900", 131=>x"7700", 132=>x"7800",
---- 133=>x"7700", 134=>x"7b00", 135=>x"7600", 136=>x"7d00",
---- 137=>x"7700", 138=>x"7900", 139=>x"7900", 140=>x"7a00",
---- 141=>x"7500", 142=>x"7700", 143=>x"7b00", 144=>x"6e00",
---- 145=>x"7000", 146=>x"7900", 147=>x"7600", 148=>x"6e00",
---- 149=>x"7200", 150=>x"7400", 151=>x"7600", 152=>x"7100",
---- 153=>x"7700", 154=>x"7800", 155=>x"7600", 156=>x"7600",
---- 157=>x"7800", 158=>x"7400", 159=>x"7400", 160=>x"7900",
---- 161=>x"7500", 162=>x"7200", 163=>x"7400", 164=>x"7a00",
---- 165=>x"7500", 166=>x"7200", 167=>x"7c00", 168=>x"7400",
---- 169=>x"7600", 170=>x"7d00", 171=>x"7800", 172=>x"7a00",
---- 173=>x"7b00", 174=>x"7a00", 175=>x"7700", 176=>x"7b00",
---- 177=>x"7500", 178=>x"7200", 179=>x"7b00", 180=>x"7500",
---- 181=>x"7200", 182=>x"7200", 183=>x"7a00", 184=>x"7700",
---- 185=>x"7600", 186=>x"7600", 187=>x"7500", 188=>x"7100",
---- 189=>x"6f00", 190=>x"6e00", 191=>x"6a00", 192=>x"6e00",
---- 193=>x"7100", 194=>x"6e00", 195=>x"7300", 196=>x"7500",
---- 197=>x"7900", 198=>x"7800", 199=>x"7b00", 200=>x"7900",
---- 201=>x"7a00", 202=>x"7600", 203=>x"7600", 204=>x"7100",
---- 205=>x"7600", 206=>x"7700", 207=>x"7700", 208=>x"7500",
---- 209=>x"7500", 210=>x"7400", 211=>x"7b00", 212=>x"7300",
---- 213=>x"8500", 214=>x"7b00", 215=>x"7b00", 216=>x"7800",
---- 217=>x"7c00", 218=>x"8000", 219=>x"7600", 220=>x"7a00",
---- 221=>x"7a00", 222=>x"7d00", 223=>x"7f00", 224=>x"7700",
---- 225=>x"7d00", 226=>x"7f00", 227=>x"7b00", 228=>x"7d00",
---- 229=>x"7c00", 230=>x"8200", 231=>x"8000", 232=>x"7d00",
---- 233=>x"8200", 234=>x"8100", 235=>x"8400", 236=>x"7d00",
---- 237=>x"8000", 238=>x"8400", 239=>x"7f00", 240=>x"8200",
---- 241=>x"7c00", 242=>x"8600", 243=>x"8300", 244=>x"8400",
---- 245=>x"8500", 246=>x"8100", 247=>x"7600", 248=>x"8400",
---- 249=>x"7d00", 250=>x"7900", 251=>x"7a00", 252=>x"7e00",
---- 253=>x"7800", 254=>x"7800", 255=>x"7400", 256=>x"7d00",
---- 257=>x"7100", 258=>x"7100", 259=>x"7b00", 260=>x"7600",
---- 261=>x"7700", 262=>x"7900", 263=>x"8600", 264=>x"7b00",
---- 265=>x"8300", 266=>x"7800", 267=>x"7e00", 268=>x"7a00",
---- 269=>x"7b00", 270=>x"8100", 271=>x"7d00", 272=>x"8100",
---- 273=>x"8100", 274=>x"8200", 275=>x"7f00", 276=>x"8100",
---- 277=>x"8000", 278=>x"7300", 279=>x"7000", 280=>x"7d00",
---- 281=>x"7000", 282=>x"6d00", 283=>x"7a00", 284=>x"6e00",
---- 285=>x"7400", 286=>x"7d00", 287=>x"7e00", 288=>x"7900",
---- 289=>x"8100", 290=>x"8200", 291=>x"7a00", 292=>x"8000",
---- 293=>x"7d00", 294=>x"7800", 295=>x"6b00", 296=>x"8200",
---- 297=>x"7800", 298=>x"6500", 299=>x"7300", 300=>x"7b00",
---- 301=>x"7000", 302=>x"7000", 303=>x"8a00", 304=>x"6c00",
---- 305=>x"7400", 306=>x"8e00", 307=>x"8900", 308=>x"7800",
---- 309=>x"9000", 310=>x"8c00", 311=>x"8e00", 312=>x"9000",
---- 313=>x"9400", 314=>x"8a00", 315=>x"8800", 316=>x"8e00",
---- 317=>x"8d00", 318=>x"8e00", 319=>x"8300", 320=>x"8600",
---- 321=>x"8a00", 322=>x"8700", 323=>x"8700", 324=>x"8a00",
---- 325=>x"8000", 326=>x"8400", 327=>x"8e00", 328=>x"8600",
---- 329=>x"7e00", 330=>x"8600", 331=>x"8f00", 332=>x"7c00",
---- 333=>x"8d00", 334=>x"8400", 335=>x"8f00", 336=>x"8e00",
---- 337=>x"8b00", 338=>x"7000", 339=>x"7700", 340=>x"8800",
---- 341=>x"6e00", 342=>x"7e00", 343=>x"7b00", 344=>x"6c00",
---- 345=>x"7500", 346=>x"7d00", 347=>x"8100", 348=>x"6c00",
---- 349=>x"7e00", 350=>x"7f00", 351=>x"8f00", 352=>x"7600",
---- 353=>x"8200", 354=>x"9000", 355=>x"8c00", 356=>x"7e00",
---- 357=>x"8c00", 358=>x"8d00", 359=>x"8900", 360=>x"8d00",
---- 361=>x"8a00", 362=>x"8600", 363=>x"8500", 364=>x"8b00",
---- 365=>x"8700", 366=>x"8600", 367=>x"8600", 368=>x"8600",
---- 369=>x"8700", 370=>x"8600", 371=>x"8a00", 372=>x"7500",
---- 373=>x"8800", 374=>x"8600", 375=>x"7b00", 376=>x"8a00",
---- 377=>x"8900", 378=>x"7800", 379=>x"7300", 380=>x"8400",
---- 381=>x"7f00", 382=>x"7000", 383=>x"7f00", 384=>x"7700",
---- 385=>x"6d00", 386=>x"7b00", 387=>x"8100", 388=>x"6a00",
---- 389=>x"7700", 390=>x"7f00", 391=>x"7d00", 392=>x"7000",
---- 393=>x"7d00", 394=>x"7f00", 395=>x"7f00", 396=>x"7b00",
---- 397=>x"7d00", 398=>x"8000", 399=>x"7f00", 400=>x"7d00",
---- 401=>x"8000", 402=>x"7b00", 403=>x"7800", 404=>x"8000",
---- 405=>x"7c00", 406=>x"7a00", 407=>x"7800", 408=>x"8200",
---- 409=>x"7d00", 410=>x"7a00", 411=>x"7a00", 412=>x"8500",
---- 413=>x"8700", 414=>x"7e00", 415=>x"8100", 416=>x"7d00",
---- 417=>x"8100", 418=>x"7500", 419=>x"7d00", 420=>x"7300",
---- 421=>x"6a00", 422=>x"7100", 423=>x"7d00", 424=>x"6b00",
---- 425=>x"7a00", 426=>x"8600", 427=>x"8700", 428=>x"8200",
---- 429=>x"8d00", 430=>x"8500", 431=>x"7f00", 432=>x"8b00",
---- 433=>x"8600", 434=>x"8600", 435=>x"8300", 436=>x"8500",
---- 437=>x"8300", 438=>x"7d00", 439=>x"7900", 440=>x"8100",
---- 441=>x"8200", 442=>x"7500", 443=>x"7b00", 444=>x"7000",
---- 445=>x"7900", 446=>x"7100", 447=>x"7200", 448=>x"5000",
---- 449=>x"5f00", 450=>x"5a00", 451=>x"4b00", 452=>x"4600",
---- 453=>x"4500", 454=>x"5500", 455=>x"3c00", 456=>x"6900",
---- 457=>x"5900", 458=>x"4700", 459=>x"2e00", 460=>x"5700",
---- 461=>x"4000", 462=>x"3400", 463=>x"3700", 464=>x"3a00",
---- 465=>x"3000", 466=>x"3800", 467=>x"5300", 468=>x"3400",
---- 469=>x"3400", 470=>x"6000", 471=>x"5d00", 472=>x"3400",
---- 473=>x"2200", 474=>x"4d00", 475=>x"5200", 476=>x"2700",
---- 477=>x"1e00", 478=>x"5100", 479=>x"5300", 480=>x"2200",
---- 481=>x"1f00", 482=>x"5700", 483=>x"6300", 484=>x"1f00",
---- 485=>x"2100", 486=>x"5300", 487=>x"7200", 488=>x"2200",
---- 489=>x"2c00", 490=>x"6200", 491=>x"6b00", 492=>x"2700",
---- 493=>x"3b00", 494=>x"8000", 495=>x"6100", 496=>x"2e00",
---- 497=>x"4f00", 498=>x"7e00", 499=>x"6800", 500=>x"4800",
---- 501=>x"5c00", 502=>x"5900", 503=>x"7000", 504=>x"6c00",
---- 505=>x"4500", 506=>x"3800", 507=>x"7f00", 508=>x"6500",
---- 509=>x"2200", 510=>x"2800", 511=>x"6e00", 512=>x"5800",
---- 513=>x"1c00", 514=>x"2400", 515=>x"4e00", 516=>x"5100",
---- 517=>x"2200", 518=>x"2c00", 519=>x"4b00", 520=>x"5300",
---- 521=>x"2100", 522=>x"2d00", 523=>x"4b00", 524=>x"4700",
---- 525=>x"2000", 526=>x"2e00", 527=>x"4900", 528=>x"3200",
---- 529=>x"d900", 530=>x"2e00", 531=>x"3a00", 532=>x"3100",
---- 533=>x"2f00", 534=>x"3000", 535=>x"2b00", 536=>x"2e00",
---- 537=>x"3000", 538=>x"2d00", 539=>x"2e00", 540=>x"2b00",
---- 541=>x"2900", 542=>x"3300", 543=>x"2f00", 544=>x"3300",
---- 545=>x"2e00", 546=>x"3500", 547=>x"2a00", 548=>x"5700",
---- 549=>x"3f00", 550=>x"3300", 551=>x"2c00", 552=>x"6000",
---- 553=>x"3b00", 554=>x"5300", 555=>x"3300", 556=>x"5600",
---- 557=>x"7b00", 558=>x"5000", 559=>x"2100", 560=>x"8700",
---- 561=>x"6900", 562=>x"2100", 563=>x"2b00", 564=>x"8000",
---- 565=>x"4e00", 566=>x"3c00", 567=>x"3c00", 568=>x"4500",
---- 569=>x"5e00", 570=>x"4a00", 571=>x"3e00", 572=>x"7400",
---- 573=>x"7400", 574=>x"2100", 575=>x"2a00", 576=>x"9e00",
---- 577=>x"4300", 578=>x"3200", 579=>x"3600", 580=>x"4e00",
---- 581=>x"5900", 582=>x"5f00", 583=>x"4e00", 584=>x"3600",
---- 585=>x"8300", 586=>x"8300", 587=>x"6700", 588=>x"4700",
---- 589=>x"7c00", 590=>x"8c00", 591=>x"7300", 592=>x"5100",
---- 593=>x"7500", 594=>x"8e00", 595=>x"6b00", 596=>x"4d00",
---- 597=>x"7700", 598=>x"8800", 599=>x"8700", 600=>x"5600",
---- 601=>x"7500", 602=>x"6f00", 603=>x"7000", 604=>x"5000",
---- 605=>x"7600", 606=>x"5d00", 607=>x"6600", 608=>x"5600",
---- 609=>x"7b00", 610=>x"7e00", 611=>x"4e00", 612=>x"5f00",
---- 613=>x"9300", 614=>x"9e00", 615=>x"6100", 616=>x"7900",
---- 617=>x"aa00", 618=>x"b600", 619=>x"8400", 620=>x"7400",
---- 621=>x"a400", 622=>x"c900", 623=>x"9c00", 624=>x"5800",
---- 625=>x"5300", 626=>x"9300", 627=>x"8200", 628=>x"4500",
---- 629=>x"4900", 630=>x"5b00", 631=>x"3a00", 632=>x"5800",
---- 633=>x"6600", 634=>x"5e00", 635=>x"3100", 636=>x"5000",
---- 637=>x"2b00", 638=>x"2700", 639=>x"2300", 640=>x"5800",
---- 641=>x"2b00", 642=>x"2300", 643=>x"2200", 644=>x"2700",
---- 645=>x"2800", 646=>x"d600", 647=>x"2b00", 648=>x"2500",
---- 649=>x"2c00", 650=>x"2e00", 651=>x"2e00", 652=>x"3200",
---- 653=>x"3800", 654=>x"3400", 655=>x"2d00", 656=>x"3f00",
---- 657=>x"4f00", 658=>x"5900", 659=>x"5f00", 660=>x"5500",
---- 661=>x"6700", 662=>x"6e00", 663=>x"8200", 664=>x"6d00",
---- 665=>x"6f00", 666=>x"8700", 667=>x"aa00", 668=>x"8400",
---- 669=>x"9c00", 670=>x"a700", 671=>x"bc00", 672=>x"a200",
---- 673=>x"a800", 674=>x"b500", 675=>x"ae00", 676=>x"ab00",
---- 677=>x"b800", 678=>x"c500", 679=>x"8400", 680=>x"ac00",
---- 681=>x"c600", 682=>x"a200", 683=>x"5b00", 684=>x"bf00",
---- 685=>x"b800", 686=>x"6400", 687=>x"5e00", 688=>x"c400",
---- 689=>x"7300", 690=>x"5f00", 691=>x"6200", 692=>x"8100",
---- 693=>x"5a00", 694=>x"6100", 695=>x"5b00", 696=>x"5900",
---- 697=>x"6a00", 698=>x"5a00", 699=>x"7000", 700=>x"6900",
---- 701=>x"6200", 702=>x"6200", 703=>x"ae00", 704=>x"5f00",
---- 705=>x"5e00", 706=>x"9b00", 707=>x"b800", 708=>x"5e00",
---- 709=>x"8d00", 710=>x"c500", 711=>x"6700", 712=>x"8f00",
---- 713=>x"c400", 714=>x"8d00", 715=>x"2e00", 716=>x"b300",
---- 717=>x"9d00", 718=>x"3c00", 719=>x"2e00", 720=>x"a000",
---- 721=>x"4400", 722=>x"2d00", 723=>x"3600", 724=>x"6100",
---- 725=>x"d200", 726=>x"3a00", 727=>x"3400", 728=>x"3000",
---- 729=>x"3600", 730=>x"3400", 731=>x"3600", 732=>x"3100",
---- 733=>x"3300", 734=>x"3100", 735=>x"3200", 736=>x"3300",
---- 737=>x"3400", 738=>x"3500", 739=>x"3300", 740=>x"3000",
---- 741=>x"3400", 742=>x"3000", 743=>x"3000", 744=>x"3300",
---- 745=>x"3800", 746=>x"3500", 747=>x"3200", 748=>x"3400",
---- 749=>x"3200", 750=>x"3300", 751=>x"3300", 752=>x"3200",
---- 753=>x"3400", 754=>x"3300", 755=>x"3300", 756=>x"3b00",
---- 757=>x"3500", 758=>x"3100", 759=>x"3500", 760=>x"c600",
---- 761=>x"3500", 762=>x"3000", 763=>x"3000", 764=>x"3500",
---- 765=>x"cb00", 766=>x"3400", 767=>x"3200", 768=>x"3100",
---- 769=>x"3400", 770=>x"3600", 771=>x"3300", 772=>x"3400",
---- 773=>x"3400", 774=>x"3700", 775=>x"3300", 776=>x"2d00",
---- 777=>x"3000", 778=>x"3200", 779=>x"3000", 780=>x"2b00",
---- 781=>x"2c00", 782=>x"3000", 783=>x"3100", 784=>x"2b00",
---- 785=>x"3300", 786=>x"3000", 787=>x"3400", 788=>x"3800",
---- 789=>x"2b00", 790=>x"3000", 791=>x"3500", 792=>x"8700",
---- 793=>x"2e00", 794=>x"2e00", 795=>x"3500", 796=>x"a800",
---- 797=>x"5f00", 798=>x"2200", 799=>x"3300", 800=>x"5900",
---- 801=>x"8400", 802=>x"3e00", 803=>x"3200", 804=>x"5800",
---- 805=>x"8500", 806=>x"7f00", 807=>x"2e00", 808=>x"3900",
---- 809=>x"6400", 810=>x"9400", 811=>x"4f00", 812=>x"2400",
---- 813=>x"3b00", 814=>x"8100", 815=>x"8900", 816=>x"6200",
---- 817=>x"2800", 818=>x"5300", 819=>x"9d00", 820=>x"b600",
---- 821=>x"4700", 822=>x"4800", 823=>x"8100", 824=>x"b600",
---- 825=>x"9400", 826=>x"5900", 827=>x"5600", 828=>x"7800",
---- 829=>x"9600", 830=>x"6100", 831=>x"2800", 832=>x"5200",
---- 833=>x"6d00", 834=>x"a700", 835=>x"2400", 836=>x"4200",
---- 837=>x"3500", 838=>x"b400", 839=>x"6200", 840=>x"2f00",
---- 841=>x"1c00", 842=>x"6000", 843=>x"8100", 844=>x"4000",
---- 845=>x"2000", 846=>x"2f00", 847=>x"7600", 848=>x"4700",
---- 849=>x"2b00", 850=>x"3300", 851=>x"8500", 852=>x"2500",
---- 853=>x"4d00", 854=>x"3400", 855=>x"7500", 856=>x"2200",
---- 857=>x"4100", 858=>x"2c00", 859=>x"6c00", 860=>x"3d00",
---- 861=>x"2400", 862=>x"2500", 863=>x"6300", 864=>x"7900",
---- 865=>x"3d00", 866=>x"2900", 867=>x"6f00", 868=>x"9b00",
---- 869=>x"6a00", 870=>x"6400", 871=>x"a200", 872=>x"7d00",
---- 873=>x"5100", 874=>x"7500", 875=>x"af00", 876=>x"8700",
---- 877=>x"8a00", 878=>x"b000", 879=>x"a000", 880=>x"8d00",
---- 881=>x"a300", 882=>x"b500", 883=>x"9300", 884=>x"6a00",
---- 885=>x"8a00", 886=>x"7c00", 887=>x"9e00", 888=>x"2100",
---- 889=>x"4400", 890=>x"5500", 891=>x"4200", 892=>x"1d00",
---- 893=>x"3000", 894=>x"5c00", 895=>x"2300", 896=>x"3300",
---- 897=>x"2b00", 898=>x"6300", 899=>x"3100", 900=>x"6500",
---- 901=>x"2500", 902=>x"6200", 903=>x"3e00", 904=>x"8f00",
---- 905=>x"5100", 906=>x"5300", 907=>x"4300", 908=>x"8000",
---- 909=>x"8000", 910=>x"6800", 911=>x"4e00", 912=>x"7900",
---- 913=>x"9100", 914=>x"8800", 915=>x"8500", 916=>x"ab00",
---- 917=>x"8300", 918=>x"a900", 919=>x"4f00", 920=>x"5400",
---- 921=>x"4d00", 922=>x"8100", 923=>x"8c00", 924=>x"7c00",
---- 925=>x"5800", 926=>x"6200", 927=>x"7200", 928=>x"6100",
---- 929=>x"5600", 930=>x"7a00", 931=>x"5600", 932=>x"4d00",
---- 933=>x"3600", 934=>x"a300", 935=>x"3e00", 936=>x"3300",
---- 937=>x"2d00", 938=>x"2b00", 939=>x"3400", 940=>x"2600",
---- 941=>x"2e00", 942=>x"2d00", 943=>x"3300", 944=>x"2e00",
---- 945=>x"2600", 946=>x"2e00", 947=>x"3600", 948=>x"2d00",
---- 949=>x"2600", 950=>x"3300", 951=>x"3500", 952=>x"3900",
---- 953=>x"2600", 954=>x"3400", 955=>x"3100", 956=>x"3f00",
---- 957=>x"2d00", 958=>x"3200", 959=>x"2c00", 960=>x"2f00",
---- 961=>x"3100", 962=>x"2e00", 963=>x"d500", 964=>x"3000",
---- 965=>x"2f00", 966=>x"2e00", 967=>x"2e00", 968=>x"2f00",
---- 969=>x"2e00", 970=>x"2d00", 971=>x"2d00", 972=>x"2a00",
---- 973=>x"2c00", 974=>x"2b00", 975=>x"d400", 976=>x"2d00",
---- 977=>x"2500", 978=>x"2900", 979=>x"3000", 980=>x"3700",
---- 981=>x"2300", 982=>x"2b00", 983=>x"3100", 984=>x"3400",
---- 985=>x"2500", 986=>x"2c00", 987=>x"2c00", 988=>x"3100",
---- 989=>x"2d00", 990=>x"3000", 991=>x"2e00", 992=>x"2c00",
---- 993=>x"2b00", 994=>x"3400", 995=>x"3600", 996=>x"2600",
---- 997=>x"2700", 998=>x"2d00", 999=>x"3100", 1000=>x"2f00",
---- 1001=>x"2b00", 1002=>x"2c00", 1003=>x"3000", 1004=>x"3800",
---- 1005=>x"2600", 1006=>x"2900", 1007=>x"2b00", 1008=>x"3b00",
---- 1009=>x"2000", 1010=>x"2100", 1011=>x"2400", 1012=>x"7500",
---- 1013=>x"3600", 1014=>x"2100", 1015=>x"2700", 1016=>x"7f00",
---- 1017=>x"7400", 1018=>x"3c00", 1019=>x"3000", 1020=>x"5b00",
---- 1021=>x"5b00", 1022=>x"6600", 1023=>x"3d00"),
----
---- 22 => (0=>x"8600", 1=>x"8600", 2=>x"8500", 3=>x"8300", 4=>x"8600",
---- 5=>x"8500", 6=>x"8600", 7=>x"8300", 8=>x"8700",
---- 9=>x"8600", 10=>x"8500", 11=>x"7c00", 12=>x"8400",
---- 13=>x"8500", 14=>x"8500", 15=>x"8300", 16=>x"8200",
---- 17=>x"8400", 18=>x"8700", 19=>x"8600", 20=>x"7b00",
---- 21=>x"8600", 22=>x"8600", 23=>x"8100", 24=>x"8500",
---- 25=>x"8400", 26=>x"8200", 27=>x"8300", 28=>x"8300",
---- 29=>x"8200", 30=>x"8200", 31=>x"8500", 32=>x"8700",
---- 33=>x"8600", 34=>x"8500", 35=>x"8400", 36=>x"8600",
---- 37=>x"8700", 38=>x"8500", 39=>x"8300", 40=>x"8400",
---- 41=>x"8200", 42=>x"8100", 43=>x"8500", 44=>x"8300",
---- 45=>x"8200", 46=>x"8200", 47=>x"8200", 48=>x"8400",
---- 49=>x"8100", 50=>x"8200", 51=>x"8100", 52=>x"8300",
---- 53=>x"8300", 54=>x"8100", 55=>x"8000", 56=>x"8300",
---- 57=>x"8200", 58=>x"8000", 59=>x"7d00", 60=>x"8100",
---- 61=>x"8200", 62=>x"8000", 63=>x"8000", 64=>x"7f00",
---- 65=>x"8100", 66=>x"8400", 67=>x"8400", 68=>x"8000",
---- 69=>x"8100", 70=>x"8100", 71=>x"8100", 72=>x"8100",
---- 73=>x"8200", 74=>x"8300", 75=>x"8200", 76=>x"8100",
---- 77=>x"8100", 78=>x"8600", 79=>x"8400", 80=>x"8000",
---- 81=>x"8000", 82=>x"8200", 83=>x"7f00", 84=>x"8300",
---- 85=>x"8100", 86=>x"8000", 87=>x"8000", 88=>x"8000",
---- 89=>x"8100", 90=>x"8100", 91=>x"8200", 92=>x"8200",
---- 93=>x"8600", 94=>x"8200", 95=>x"7e00", 96=>x"8200",
---- 97=>x"8400", 98=>x"8100", 99=>x"8000", 100=>x"8700",
---- 101=>x"7f00", 102=>x"8000", 103=>x"8100", 104=>x"8200",
---- 105=>x"8000", 106=>x"7f00", 107=>x"7e00", 108=>x"7d00",
---- 109=>x"7c00", 110=>x"7d00", 111=>x"7f00", 112=>x"8800",
---- 113=>x"8900", 114=>x"8800", 115=>x"8100", 116=>x"9400",
---- 117=>x"8900", 118=>x"7d00", 119=>x"7500", 120=>x"8100",
---- 121=>x"7e00", 122=>x"7900", 123=>x"7a00", 124=>x"7f00",
---- 125=>x"7d00", 126=>x"7900", 127=>x"7a00", 128=>x"7c00",
---- 129=>x"7a00", 130=>x"7d00", 131=>x"7c00", 132=>x"7a00",
---- 133=>x"7900", 134=>x"7a00", 135=>x"7600", 136=>x"8000",
---- 137=>x"7a00", 138=>x"7600", 139=>x"7700", 140=>x"7b00",
---- 141=>x"7c00", 142=>x"7600", 143=>x"7b00", 144=>x"7900",
---- 145=>x"7c00", 146=>x"8000", 147=>x"7e00", 148=>x"7c00",
---- 149=>x"8300", 150=>x"7d00", 151=>x"7700", 152=>x"7b00",
---- 153=>x"7a00", 154=>x"7a00", 155=>x"8000", 156=>x"7100",
---- 157=>x"7b00", 158=>x"7e00", 159=>x"8100", 160=>x"7700",
---- 161=>x"7e00", 162=>x"7c00", 163=>x"7d00", 164=>x"7c00",
---- 165=>x"7600", 166=>x"7d00", 167=>x"7800", 168=>x"7600",
---- 169=>x"7900", 170=>x"7a00", 171=>x"7500", 172=>x"7a00",
---- 173=>x"7700", 174=>x"7800", 175=>x"7800", 176=>x"7800",
---- 177=>x"7400", 178=>x"7300", 179=>x"7100", 180=>x"6f00",
---- 181=>x"7100", 182=>x"7400", 183=>x"7a00", 184=>x"6b00",
---- 185=>x"6e00", 186=>x"7900", 187=>x"8000", 188=>x"7100",
---- 189=>x"7600", 190=>x"7800", 191=>x"8000", 192=>x"7700",
---- 193=>x"7800", 194=>x"7900", 195=>x"7c00", 196=>x"7500",
---- 197=>x"7c00", 198=>x"7e00", 199=>x"8400", 200=>x"7700",
---- 201=>x"7c00", 202=>x"8200", 203=>x"8200", 204=>x"8000",
---- 205=>x"8900", 206=>x"8400", 207=>x"8100", 208=>x"8400",
---- 209=>x"8200", 210=>x"7f00", 211=>x"8600", 212=>x"7b00",
---- 213=>x"8200", 214=>x"8900", 215=>x"8500", 216=>x"7d00",
---- 217=>x"8300", 218=>x"8700", 219=>x"8300", 220=>x"7e00",
---- 221=>x"7e00", 222=>x"8700", 223=>x"8d00", 224=>x"8400",
---- 225=>x"8600", 226=>x"8f00", 227=>x"8b00", 228=>x"8600",
---- 229=>x"8700", 230=>x"8300", 231=>x"8600", 232=>x"8b00",
---- 233=>x"8a00", 234=>x"8400", 235=>x"8500", 236=>x"8a00",
---- 237=>x"8d00", 238=>x"8300", 239=>x"8500", 240=>x"8000",
---- 241=>x"7d00", 242=>x"8700", 243=>x"7800", 244=>x"7c00",
---- 245=>x"7e00", 246=>x"6c00", 247=>x"7100", 248=>x"7700",
---- 249=>x"7100", 250=>x"8700", 251=>x"8700", 252=>x"7400",
---- 253=>x"8300", 254=>x"8d00", 255=>x"8600", 256=>x"8000",
---- 257=>x"8600", 258=>x"8800", 259=>x"7a00", 260=>x"8400",
---- 261=>x"8400", 262=>x"8600", 263=>x"8b00", 264=>x"8600",
---- 265=>x"8500", 266=>x"8300", 267=>x"8100", 268=>x"8300",
---- 269=>x"7700", 270=>x"7200", 271=>x"7d00", 272=>x"7400",
---- 273=>x"7600", 274=>x"7800", 275=>x"7400", 276=>x"7800",
---- 277=>x"7b00", 278=>x"7500", 279=>x"6900", 280=>x"7600",
---- 281=>x"7200", 282=>x"7100", 283=>x"7f00", 284=>x"7a00",
---- 285=>x"6f00", 286=>x"7e00", 287=>x"9c00", 288=>x"6b00",
---- 289=>x"7900", 290=>x"9400", 291=>x"9600", 292=>x"7800",
---- 293=>x"9500", 294=>x"9000", 295=>x"9400", 296=>x"9300",
---- 297=>x"9700", 298=>x"9300", 299=>x"9100", 300=>x"9200",
---- 301=>x"9400", 302=>x"9700", 303=>x"8c00", 304=>x"9000",
---- 305=>x"9700", 306=>x"8e00", 307=>x"8b00", 308=>x"9300",
---- 309=>x"8f00", 310=>x"8b00", 311=>x"8a00", 312=>x"8d00",
---- 313=>x"8900", 314=>x"9200", 315=>x"9900", 316=>x"8400",
---- 317=>x"8d00", 318=>x"9b00", 319=>x"7e00", 320=>x"8a00",
---- 321=>x"9400", 322=>x"7a00", 323=>x"7200", 324=>x"8c00",
---- 325=>x"7500", 326=>x"7100", 327=>x"7900", 328=>x"6d00",
---- 329=>x"7c00", 330=>x"7f00", 331=>x"8a00", 332=>x"7300",
---- 333=>x"8600", 334=>x"8800", 335=>x"9700", 336=>x"7800",
---- 337=>x"8800", 338=>x"8e00", 339=>x"8a00", 340=>x"8600",
---- 341=>x"9400", 342=>x"8b00", 343=>x"8700", 344=>x"6b00",
---- 345=>x"9000", 346=>x"8a00", 347=>x"8c00", 348=>x"7400",
---- 349=>x"8f00", 350=>x"8b00", 351=>x"8400", 352=>x"8800",
---- 353=>x"8500", 354=>x"8900", 355=>x"8800", 356=>x"8900",
---- 357=>x"8800", 358=>x"8900", 359=>x"7e00", 360=>x"8900",
---- 361=>x"8f00", 362=>x"7b00", 363=>x"7800", 364=>x"8900",
---- 365=>x"7d00", 366=>x"7500", 367=>x"8500", 368=>x"7c00",
---- 369=>x"6f00", 370=>x"7b00", 371=>x"8200", 372=>x"7400",
---- 373=>x"7f00", 374=>x"8000", 375=>x"8300", 376=>x"8200",
---- 377=>x"7c00", 378=>x"8200", 379=>x"8500", 380=>x"7f00",
---- 381=>x"7d00", 382=>x"8000", 383=>x"8700", 384=>x"8100",
---- 385=>x"8000", 386=>x"8000", 387=>x"8500", 388=>x"8400",
---- 389=>x"8300", 390=>x"7900", 391=>x"7e00", 392=>x"7d00",
---- 393=>x"8100", 394=>x"7f00", 395=>x"7800", 396=>x"7500",
---- 397=>x"7d00", 398=>x"8000", 399=>x"7500", 400=>x"7400",
---- 401=>x"8300", 402=>x"7800", 403=>x"7b00", 404=>x"7900",
---- 405=>x"7d00", 406=>x"8600", 407=>x"7500", 408=>x"7800",
---- 409=>x"7900", 410=>x"8600", 411=>x"8900", 412=>x"7700",
---- 413=>x"7600", 414=>x"8600", 415=>x"8100", 416=>x"8000",
---- 417=>x"7f00", 418=>x"7000", 419=>x"6b00", 420=>x"8200",
---- 421=>x"8400", 422=>x"8300", 423=>x"8300", 424=>x"8200",
---- 425=>x"7200", 426=>x"6300", 427=>x"8a00", 428=>x"8200",
---- 429=>x"6f00", 430=>x"6000", 431=>x"7a00", 432=>x"7700",
---- 433=>x"6400", 434=>x"5900", 435=>x"6500", 436=>x"7d00",
---- 437=>x"5a00", 438=>x"3300", 439=>x"3c00", 440=>x"7f00",
---- 441=>x"5d00", 442=>x"2a00", 443=>x"2a00", 444=>x"6f00",
---- 445=>x"6100", 446=>x"3200", 447=>x"2800", 448=>x"4700",
---- 449=>x"4e00", 450=>x"3c00", 451=>x"2d00", 452=>x"3f00",
---- 453=>x"4e00", 454=>x"3800", 455=>x"2800", 456=>x"3000",
---- 457=>x"2e00", 458=>x"2700", 459=>x"3000", 460=>x"3c00",
---- 461=>x"2800", 462=>x"2900", 463=>x"d600", 464=>x"3900",
---- 465=>x"2400", 466=>x"2900", 467=>x"2600", 468=>x"2a00",
---- 469=>x"2700", 470=>x"2c00", 471=>x"2700", 472=>x"2500",
---- 473=>x"3700", 474=>x"3900", 475=>x"2d00", 476=>x"2b00",
---- 477=>x"4c00", 478=>x"2e00", 479=>x"3400", 480=>x"3a00",
---- 481=>x"3100", 482=>x"2b00", 483=>x"3400", 484=>x"3900",
---- 485=>x"2100", 486=>x"3100", 487=>x"2700", 488=>x"2400",
---- 489=>x"2800", 490=>x"3300", 491=>x"3500", 492=>x"1c00",
---- 493=>x"3000", 494=>x"3200", 495=>x"3100", 496=>x"1c00",
---- 497=>x"2b00", 498=>x"2800", 499=>x"2e00", 500=>x"1e00",
---- 501=>x"2600", 502=>x"2c00", 503=>x"4800", 504=>x"3400",
---- 505=>x"2400", 506=>x"3000", 507=>x"4700", 508=>x"5000",
---- 509=>x"2600", 510=>x"2c00", 511=>x"4b00", 512=>x"5800",
---- 513=>x"2b00", 514=>x"2c00", 515=>x"5400", 516=>x"4c00",
---- 517=>x"3a00", 518=>x"2600", 519=>x"5800", 520=>x"3100",
---- 521=>x"4700", 522=>x"3000", 523=>x"5a00", 524=>x"2e00",
---- 525=>x"3b00", 526=>x"4200", 527=>x"5f00", 528=>x"3000",
---- 529=>x"2f00", 530=>x"2a00", 531=>x"5500", 532=>x"2600",
---- 533=>x"3100", 534=>x"2600", 535=>x"3f00", 536=>x"2d00",
---- 537=>x"2f00", 538=>x"2700", 539=>x"3000", 540=>x"3500",
---- 541=>x"3200", 542=>x"2800", 543=>x"2b00", 544=>x"3800",
---- 545=>x"3000", 546=>x"2c00", 547=>x"2c00", 548=>x"3300",
---- 549=>x"2700", 550=>x"2500", 551=>x"2c00", 552=>x"2c00",
---- 553=>x"2700", 554=>x"2800", 555=>x"2d00", 556=>x"2d00",
---- 557=>x"2c00", 558=>x"2e00", 559=>x"2a00", 560=>x"3500",
---- 561=>x"2d00", 562=>x"3100", 563=>x"3000", 564=>x"2e00",
---- 565=>x"2c00", 566=>x"2f00", 567=>x"3000", 568=>x"2f00",
---- 569=>x"2a00", 570=>x"2c00", 571=>x"2d00", 572=>x"2f00",
---- 573=>x"2e00", 574=>x"3000", 575=>x"2d00", 576=>x"3400",
---- 577=>x"2f00", 578=>x"3400", 579=>x"3300", 580=>x"4c00",
---- 581=>x"2c00", 582=>x"2a00", 583=>x"3500", 584=>x"5b00",
---- 585=>x"3400", 586=>x"2e00", 587=>x"3200", 588=>x"4b00",
---- 589=>x"3500", 590=>x"2b00", 591=>x"2e00", 592=>x"5f00",
---- 593=>x"3e00", 594=>x"2b00", 595=>x"2b00", 596=>x"7b00",
---- 597=>x"3200", 598=>x"2d00", 599=>x"2a00", 600=>x"9700",
---- 601=>x"5100", 602=>x"2000", 603=>x"2500", 604=>x"ac00",
---- 605=>x"9200", 606=>x"4500", 607=>x"2800", 608=>x"7400",
---- 609=>x"9b00", 610=>x"9a00", 611=>x"3b00", 612=>x"3600",
---- 613=>x"7500", 614=>x"aa00", 615=>x"5e00", 616=>x"2f00",
---- 617=>x"4d00", 618=>x"8600", 619=>x"5400", 620=>x"3500",
---- 621=>x"3300", 622=>x"6400", 623=>x"3200", 624=>x"3b00",
---- 625=>x"2500", 626=>x"3700", 627=>x"2600", 628=>x"2a00",
---- 629=>x"2800", 630=>x"3300", 631=>x"2200", 632=>x"2300",
---- 633=>x"2900", 634=>x"2900", 635=>x"1d00", 636=>x"2400",
---- 637=>x"2b00", 638=>x"1c00", 639=>x"3800", 640=>x"2900",
---- 641=>x"2400", 642=>x"1600", 643=>x"6300", 644=>x"2700",
---- 645=>x"1f00", 646=>x"1d00", 647=>x"8e00", 648=>x"2300",
---- 649=>x"1800", 650=>x"3d00", 651=>x"a100", 652=>x"3200",
---- 653=>x"3400", 654=>x"6700", 655=>x"8f00", 656=>x"6300",
---- 657=>x"7700", 658=>x"7200", 659=>x"7400", 660=>x"9f00",
---- 661=>x"9c00", 662=>x"6800", 663=>x"6800", 664=>x"b700",
---- 665=>x"6e00", 666=>x"6500", 667=>x"6b00", 668=>x"8800",
---- 669=>x"5700", 670=>x"5e00", 671=>x"7300", 672=>x"5d00",
---- 673=>x"5e00", 674=>x"5700", 675=>x"6900", 676=>x"5d00",
---- 677=>x"a200", 678=>x"5900", 679=>x"9900", 680=>x"5e00",
---- 681=>x"5700", 682=>x"7a00", 683=>x"b300", 684=>x"5800",
---- 685=>x"6500", 686=>x"b400", 687=>x"5e00", 688=>x"6400",
---- 689=>x"5f00", 690=>x"8e00", 691=>x"2500", 692=>x"8c00",
---- 693=>x"ae00", 694=>x"3500", 695=>x"2700", 696=>x"ba00",
---- 697=>x"5c00", 698=>x"1c00", 699=>x"2700", 700=>x"9a00",
---- 701=>x"2300", 702=>x"2f00", 703=>x"3000", 704=>x"4000",
---- 705=>x"2600", 706=>x"2f00", 707=>x"3200", 708=>x"2200",
---- 709=>x"3400", 710=>x"3500", 711=>x"3300", 712=>x"3400",
---- 713=>x"3400", 714=>x"3600", 715=>x"3500", 716=>x"3300",
---- 717=>x"3300", 718=>x"3300", 719=>x"3500", 720=>x"3000",
---- 721=>x"3200", 722=>x"3700", 723=>x"3800", 724=>x"3500",
---- 725=>x"3600", 726=>x"3b00", 727=>x"3700", 728=>x"3600",
---- 729=>x"3700", 730=>x"3a00", 731=>x"3b00", 732=>x"3300",
---- 733=>x"3400", 734=>x"3700", 735=>x"3900", 736=>x"3100",
---- 737=>x"3800", 738=>x"3900", 739=>x"3900", 740=>x"2e00",
---- 741=>x"3400", 742=>x"3900", 743=>x"3500", 744=>x"3200",
---- 745=>x"3400", 746=>x"3900", 747=>x"3b00", 748=>x"3000",
---- 749=>x"3500", 750=>x"4000", 751=>x"3800", 752=>x"2f00",
---- 753=>x"3e00", 754=>x"4700", 755=>x"3800", 756=>x"3200",
---- 757=>x"3900", 758=>x"c000", 759=>x"3d00", 760=>x"3000",
---- 761=>x"3900", 762=>x"3e00", 763=>x"c000", 764=>x"3600",
---- 765=>x"3d00", 766=>x"4200", 767=>x"4800", 768=>x"3700",
---- 769=>x"3d00", 770=>x"4800", 771=>x"4a00", 772=>x"3800",
---- 773=>x"4800", 774=>x"b300", 775=>x"4a00", 776=>x"3600",
---- 777=>x"4c00", 778=>x"4d00", 779=>x"4c00", 780=>x"3400",
---- 781=>x"4500", 782=>x"4e00", 783=>x"4700", 784=>x"3a00",
---- 785=>x"4600", 786=>x"5500", 787=>x"4300", 788=>x"4200",
---- 789=>x"4600", 790=>x"5800", 791=>x"4000", 792=>x"c600",
---- 793=>x"4100", 794=>x"5100", 795=>x"3b00", 796=>x"3700",
---- 797=>x"4000", 798=>x"ac00", 799=>x"3800", 800=>x"3700",
---- 801=>x"c000", 802=>x"5100", 803=>x"3600", 804=>x"3400",
---- 805=>x"4200", 806=>x"4900", 807=>x"3400", 808=>x"3100",
---- 809=>x"4400", 810=>x"4000", 811=>x"3100", 812=>x"3000",
---- 813=>x"3d00", 814=>x"3e00", 815=>x"3600", 816=>x"5400",
---- 817=>x"3300", 818=>x"3a00", 819=>x"2f00", 820=>x"8100",
---- 821=>x"2c00", 822=>x"3300", 823=>x"2c00", 824=>x"9b00",
---- 825=>x"3f00", 826=>x"2f00", 827=>x"2e00", 828=>x"9800",
---- 829=>x"6800", 830=>x"d800", 831=>x"3000", 832=>x"8300",
---- 833=>x"9d00", 834=>x"2200", 835=>x"2800", 836=>x"6b00",
---- 837=>x"c000", 838=>x"2e00", 839=>x"2200", 840=>x"6600",
---- 841=>x"c700", 842=>x"3b00", 843=>x"1d00", 844=>x"7700",
---- 845=>x"d300", 846=>x"4f00", 847=>x"2100", 848=>x"9d00",
---- 849=>x"cf00", 850=>x"5e00", 851=>x"1f00", 852=>x"ba00",
---- 853=>x"c800", 854=>x"4f00", 855=>x"1d00", 856=>x"c200",
---- 857=>x"ba00", 858=>x"3f00", 859=>x"1f00", 860=>x"c600",
---- 861=>x"9000", 862=>x"2d00", 863=>x"2200", 864=>x"b500",
---- 865=>x"5700", 866=>x"5e00", 867=>x"3900", 868=>x"9800",
---- 869=>x"6e00", 870=>x"c100", 871=>x"5500", 872=>x"9000",
---- 873=>x"8b00", 874=>x"9d00", 875=>x"3f00", 876=>x"4900",
---- 877=>x"2900", 878=>x"2800", 879=>x"2d00", 880=>x"5d00",
---- 881=>x"3000", 882=>x"2500", 883=>x"4f00", 884=>x"b400",
---- 885=>x"8700", 886=>x"7b00", 887=>x"7700", 888=>x"5400",
---- 889=>x"6000", 890=>x"8100", 891=>x"7200", 892=>x"2200",
---- 893=>x"4000", 894=>x"2f00", 895=>x"2000", 896=>x"3000",
---- 897=>x"4200", 898=>x"1f00", 899=>x"2800", 900=>x"2e00",
---- 901=>x"2f00", 902=>x"2800", 903=>x"3900", 904=>x"2e00",
---- 905=>x"2400", 906=>x"2c00", 907=>x"4100", 908=>x"7500",
---- 909=>x"3900", 910=>x"2400", 911=>x"3e00", 912=>x"a000",
---- 913=>x"3000", 914=>x"2b00", 915=>x"3400", 916=>x"6300",
---- 917=>x"2300", 918=>x"3300", 919=>x"3700", 920=>x"2d00",
---- 921=>x"2900", 922=>x"3500", 923=>x"3600", 924=>x"2700",
---- 925=>x"2f00", 926=>x"3900", 927=>x"3600", 928=>x"2200",
---- 929=>x"3100", 930=>x"3500", 931=>x"2b00", 932=>x"2a00",
---- 933=>x"3100", 934=>x"3100", 935=>x"2400", 936=>x"3900",
---- 937=>x"3800", 938=>x"2c00", 939=>x"2900", 940=>x"3a00",
---- 941=>x"3400", 942=>x"2b00", 943=>x"2d00", 944=>x"3200",
---- 945=>x"2c00", 946=>x"2f00", 947=>x"3200", 948=>x"2800",
---- 949=>x"2a00", 950=>x"2d00", 951=>x"2f00", 952=>x"2b00",
---- 953=>x"2c00", 954=>x"2b00", 955=>x"2600", 956=>x"2b00",
---- 957=>x"2a00", 958=>x"2c00", 959=>x"2a00", 960=>x"2c00",
---- 961=>x"2b00", 962=>x"2b00", 963=>x"2e00", 964=>x"3300",
---- 965=>x"2d00", 966=>x"2a00", 967=>x"2d00", 968=>x"2e00",
---- 969=>x"2f00", 970=>x"2900", 971=>x"2800", 972=>x"3300",
---- 973=>x"2a00", 974=>x"2700", 975=>x"2700", 976=>x"2d00",
---- 977=>x"2700", 978=>x"2600", 979=>x"2d00", 980=>x"2a00",
---- 981=>x"2f00", 982=>x"2e00", 983=>x"2a00", 984=>x"2900",
---- 985=>x"3100", 986=>x"3100", 987=>x"2c00", 988=>x"3000",
---- 989=>x"2c00", 990=>x"2a00", 991=>x"2900", 992=>x"2b00",
---- 993=>x"2700", 994=>x"2700", 995=>x"2800", 996=>x"2500",
---- 997=>x"2c00", 998=>x"3200", 999=>x"2f00", 1000=>x"3300",
---- 1001=>x"2e00", 1002=>x"3100", 1003=>x"3100", 1004=>x"2f00",
---- 1005=>x"3200", 1006=>x"3400", 1007=>x"3700", 1008=>x"2a00",
---- 1009=>x"3200", 1010=>x"3c00", 1011=>x"4b00", 1012=>x"2b00",
---- 1013=>x"3600", 1014=>x"4300", 1015=>x"4d00", 1016=>x"3900",
---- 1017=>x"4b00", 1018=>x"5000", 1019=>x"5300", 1020=>x"4500",
---- 1021=>x"5400", 1022=>x"5100", 1023=>x"5a00"),
----
---- 23 => (0=>x"8500", 1=>x"8800", 2=>x"8400", 3=>x"7b00", 4=>x"8500",
---- 5=>x"8800", 6=>x"8500", 7=>x"8400", 8=>x"8500",
---- 9=>x"8600", 10=>x"8500", 11=>x"8400", 12=>x"8200",
---- 13=>x"8200", 14=>x"8200", 15=>x"8300", 16=>x"8100",
---- 17=>x"8600", 18=>x"8500", 19=>x"8400", 20=>x"8200",
---- 21=>x"8500", 22=>x"8400", 23=>x"8300", 24=>x"8500",
---- 25=>x"8300", 26=>x"8300", 27=>x"8400", 28=>x"8500",
---- 29=>x"8400", 30=>x"8700", 31=>x"8200", 32=>x"8400",
---- 33=>x"8500", 34=>x"8600", 35=>x"8400", 36=>x"8300",
---- 37=>x"8300", 38=>x"8500", 39=>x"8400", 40=>x"8200",
---- 41=>x"8200", 42=>x"8400", 43=>x"8200", 44=>x"8100",
---- 45=>x"8000", 46=>x"8500", 47=>x"8200", 48=>x"8200",
---- 49=>x"8000", 50=>x"8300", 51=>x"8300", 52=>x"8100",
---- 53=>x"8300", 54=>x"8400", 55=>x"8500", 56=>x"8100",
---- 57=>x"8200", 58=>x"8100", 59=>x"8400", 60=>x"8200",
---- 61=>x"7c00", 62=>x"8100", 63=>x"8400", 64=>x"8100",
---- 65=>x"7f00", 66=>x"8300", 67=>x"8200", 68=>x"8000",
---- 69=>x"8100", 70=>x"8000", 71=>x"8100", 72=>x"8100",
---- 73=>x"8100", 74=>x"7f00", 75=>x"8100", 76=>x"8300",
---- 77=>x"8000", 78=>x"8000", 79=>x"7f00", 80=>x"8000",
---- 81=>x"8100", 82=>x"7f00", 83=>x"8000", 84=>x"8200",
---- 85=>x"8000", 86=>x"7f00", 87=>x"8100", 88=>x"8000",
---- 89=>x"8100", 90=>x"7e00", 91=>x"7e00", 92=>x"8000",
---- 93=>x"7f00", 94=>x"8100", 95=>x"7f00", 96=>x"8000",
---- 97=>x"8000", 98=>x"8000", 99=>x"7e00", 100=>x"7f00",
---- 101=>x"7f00", 102=>x"7c00", 103=>x"7a00", 104=>x"7e00",
---- 105=>x"7d00", 106=>x"8100", 107=>x"8800", 108=>x"8000",
---- 109=>x"8000", 110=>x"8a00", 111=>x"9500", 112=>x"7f00",
---- 113=>x"8600", 114=>x"9500", 115=>x"9100", 116=>x"7e00",
---- 117=>x"8600", 118=>x"8b00", 119=>x"8a00", 120=>x"7b00",
---- 121=>x"7d00", 122=>x"8400", 123=>x"8700", 124=>x"7900",
---- 125=>x"7e00", 126=>x"8a00", 127=>x"8700", 128=>x"7e00",
---- 129=>x"8200", 130=>x"8800", 131=>x"8300", 132=>x"7900",
---- 133=>x"8500", 134=>x"8500", 135=>x"8400", 136=>x"7b00",
---- 137=>x"7e00", 138=>x"8100", 139=>x"8500", 140=>x"8000",
---- 141=>x"8400", 142=>x"8800", 143=>x"8600", 144=>x"7900",
---- 145=>x"8700", 146=>x"8100", 147=>x"8200", 148=>x"8500",
---- 149=>x"8100", 150=>x"7500", 151=>x"8100", 152=>x"7e00",
---- 153=>x"7a00", 154=>x"7f00", 155=>x"8300", 156=>x"7900",
---- 157=>x"7c00", 158=>x"8300", 159=>x"8300", 160=>x"7900",
---- 161=>x"7f00", 162=>x"8000", 163=>x"8100", 164=>x"7600",
---- 165=>x"7d00", 166=>x"7800", 167=>x"7c00", 168=>x"7800",
---- 169=>x"7800", 170=>x"7800", 171=>x"7a00", 172=>x"7400",
---- 173=>x"7700", 174=>x"8000", 175=>x"7d00", 176=>x"7400",
---- 177=>x"7d00", 178=>x"7d00", 179=>x"8400", 180=>x"7700",
---- 181=>x"7f00", 182=>x"8300", 183=>x"7900", 184=>x"8000",
---- 185=>x"8000", 186=>x"7d00", 187=>x"7f00", 188=>x"8400",
---- 189=>x"7e00", 190=>x"8100", 191=>x"8200", 192=>x"8100",
---- 193=>x"8100", 194=>x"7f00", 195=>x"8500", 196=>x"7f00",
---- 197=>x"7a00", 198=>x"8100", 199=>x"8000", 200=>x"8000",
---- 201=>x"7f00", 202=>x"7d00", 203=>x"8600", 204=>x"7f00",
---- 205=>x"8800", 206=>x"8900", 207=>x"8b00", 208=>x"8900",
---- 209=>x"8c00", 210=>x"9100", 211=>x"9000", 212=>x"8700",
---- 213=>x"9000", 214=>x"9000", 215=>x"8c00", 216=>x"8c00",
---- 217=>x"9400", 218=>x"8d00", 219=>x"8200", 220=>x"9200",
---- 221=>x"8900", 222=>x"7f00", 223=>x"8200", 224=>x"8500",
---- 225=>x"8200", 226=>x"8800", 227=>x"8200", 228=>x"8b00",
---- 229=>x"8d00", 230=>x"8800", 231=>x"8800", 232=>x"8f00",
---- 233=>x"8d00", 234=>x"8000", 235=>x"7f00", 236=>x"8500",
---- 237=>x"7d00", 238=>x"8100", 239=>x"8700", 240=>x"7300",
---- 241=>x"8300", 242=>x"8900", 243=>x"8800", 244=>x"8700",
---- 245=>x"8d00", 246=>x"8800", 247=>x"7b00", 248=>x"8b00",
---- 249=>x"8300", 250=>x"7b00", 251=>x"7f00", 252=>x"7900",
---- 253=>x"7700", 254=>x"8200", 255=>x"8100", 256=>x"7900",
---- 257=>x"8600", 258=>x"8300", 259=>x"7600", 260=>x"8600",
---- 261=>x"8400", 262=>x"7700", 263=>x"6700", 264=>x"8000",
---- 265=>x"7800", 266=>x"5f00", 267=>x"6a00", 268=>x"7900",
---- 269=>x"6100", 270=>x"6d00", 271=>x"8d00", 272=>x"6600",
---- 273=>x"7400", 274=>x"9300", 275=>x"a000", 276=>x"7600",
---- 277=>x"8c00", 278=>x"9700", 279=>x"9d00", 280=>x"9500",
---- 281=>x"9000", 282=>x"9400", 283=>x"9a00", 284=>x"9300",
---- 285=>x"9700", 286=>x"9300", 287=>x"9200", 288=>x"9400",
---- 289=>x"9c00", 290=>x"9600", 291=>x"8600", 292=>x"9900",
---- 293=>x"9700", 294=>x"8e00", 295=>x"8700", 296=>x"9100",
---- 297=>x"8d00", 298=>x"8e00", 299=>x"9800", 300=>x"8200",
---- 301=>x"8b00", 302=>x"9f00", 303=>x"8e00", 304=>x"8900",
---- 305=>x"9a00", 306=>x"8b00", 307=>x"7200", 308=>x"9c00",
---- 309=>x"8400", 310=>x"6e00", 311=>x"8100", 312=>x"7800",
---- 313=>x"7100", 314=>x"8200", 315=>x"9300", 316=>x"6b00",
---- 317=>x"7e00", 318=>x"8f00", 319=>x"9400", 320=>x"7e00",
---- 321=>x"8c00", 322=>x"8a00", 323=>x"9200", 324=>x"8b00",
---- 325=>x"9300", 326=>x"8c00", 327=>x"8e00", 328=>x"8e00",
---- 329=>x"8f00", 330=>x"9600", 331=>x"8d00", 332=>x"8f00",
---- 333=>x"8e00", 334=>x"9600", 335=>x"8d00", 336=>x"9000",
---- 337=>x"9700", 338=>x"8b00", 339=>x"8c00", 340=>x"8e00",
---- 341=>x"8c00", 342=>x"8800", 343=>x"8d00", 344=>x"8b00",
---- 345=>x"8f00", 346=>x"8c00", 347=>x"7300", 348=>x"8e00",
---- 349=>x"8700", 350=>x"7800", 351=>x"8000", 352=>x"8000",
---- 353=>x"7500", 354=>x"7800", 355=>x"8500", 356=>x"7000",
---- 357=>x"8100", 358=>x"8300", 359=>x"8100", 360=>x"8000",
---- 361=>x"8200", 362=>x"8100", 363=>x"8800", 364=>x"8300",
---- 365=>x"8600", 366=>x"8300", 367=>x"8400", 368=>x"8600",
---- 369=>x"8800", 370=>x"8800", 371=>x"8300", 372=>x"8700",
---- 373=>x"8600", 374=>x"8400", 375=>x"8300", 376=>x"8300",
---- 377=>x"8500", 378=>x"8000", 379=>x"7700", 380=>x"8400",
---- 381=>x"7d00", 382=>x"7800", 383=>x"8200", 384=>x"8100",
---- 385=>x"7900", 386=>x"7800", 387=>x"8a00", 388=>x"7d00",
---- 389=>x"7300", 390=>x"8700", 391=>x"8d00", 392=>x"7300",
---- 393=>x"7b00", 394=>x"7f00", 395=>x"6e00", 396=>x"7e00",
---- 397=>x"8f00", 398=>x"8900", 399=>x"8400", 400=>x"8800",
---- 401=>x"8d00", 402=>x"8f00", 403=>x"8c00", 404=>x"8700",
---- 405=>x"8400", 406=>x"8100", 407=>x"7700", 408=>x"7800",
---- 409=>x"6c00", 410=>x"6a00", 411=>x"6f00", 412=>x"8000",
---- 413=>x"8000", 414=>x"7f00", 415=>x"7000", 416=>x"7d00",
---- 417=>x"7b00", 418=>x"6e00", 419=>x"5300", 420=>x"7100",
---- 421=>x"6600", 422=>x"4b00", 423=>x"4100", 424=>x"8300",
---- 425=>x"6c00", 426=>x"4800", 427=>x"4200", 428=>x"6f00",
---- 429=>x"6100", 430=>x"4800", 431=>x"4600", 432=>x"4a00",
---- 433=>x"3f00", 434=>x"5500", 435=>x"5000", 436=>x"3000",
---- 437=>x"3700", 438=>x"5a00", 439=>x"3e00", 440=>x"3300",
---- 441=>x"4900", 442=>x"4900", 443=>x"3100", 444=>x"4000",
---- 445=>x"5f00", 446=>x"3800", 447=>x"2800", 448=>x"5000",
---- 449=>x"5d00", 450=>x"2e00", 451=>x"2900", 452=>x"5f00",
---- 453=>x"5200", 454=>x"2a00", 455=>x"2a00", 456=>x"6100",
---- 457=>x"b500", 458=>x"2500", 459=>x"2b00", 460=>x"5500",
---- 461=>x"4800", 462=>x"2400", 463=>x"3100", 464=>x"4a00",
---- 465=>x"5800", 466=>x"3c00", 467=>x"4300", 468=>x"3300",
---- 469=>x"6200", 470=>x"4700", 471=>x"2e00", 472=>x"2800",
---- 473=>x"3800", 474=>x"5200", 475=>x"2c00", 476=>x"2900",
---- 477=>x"2600", 478=>x"3600", 479=>x"5100", 480=>x"3d00",
---- 481=>x"3700", 482=>x"4d00", 483=>x"6600", 484=>x"3e00",
---- 485=>x"5a00", 486=>x"6800", 487=>x"5100", 488=>x"4600",
---- 489=>x"4500", 490=>x"3900", 491=>x"3a00", 492=>x"3500",
---- 493=>x"2f00", 494=>x"3200", 495=>x"3b00", 496=>x"4000",
---- 497=>x"4500", 498=>x"3200", 499=>x"4200", 500=>x"4600",
---- 501=>x"3d00", 502=>x"4300", 503=>x"3d00", 504=>x"3d00",
---- 505=>x"2f00", 506=>x"3600", 507=>x"4200", 508=>x"3900",
---- 509=>x"2500", 510=>x"2500", 511=>x"3700", 512=>x"3d00",
---- 513=>x"2700", 514=>x"2500", 515=>x"3000", 516=>x"3b00",
---- 517=>x"2300", 518=>x"2500", 519=>x"2a00", 520=>x"4300",
---- 521=>x"2400", 522=>x"2700", 523=>x"2400", 524=>x"5300",
---- 525=>x"2600", 526=>x"2f00", 527=>x"2700", 528=>x"6500",
---- 529=>x"2900", 530=>x"2f00", 531=>x"2d00", 532=>x"7400",
---- 533=>x"3800", 534=>x"3300", 535=>x"2600", 536=>x"6f00",
---- 537=>x"5200", 538=>x"2e00", 539=>x"2900", 540=>x"5900",
---- 541=>x"4f00", 542=>x"2800", 543=>x"3400", 544=>x"3c00",
---- 545=>x"3500", 546=>x"2e00", 547=>x"3b00", 548=>x"3300",
---- 549=>x"2f00", 550=>x"3900", 551=>x"3a00", 552=>x"3100",
---- 553=>x"2e00", 554=>x"3100", 555=>x"2e00", 556=>x"2d00",
---- 557=>x"2f00", 558=>x"3000", 559=>x"2b00", 560=>x"2d00",
---- 561=>x"3000", 562=>x"2e00", 563=>x"2d00", 564=>x"2e00",
---- 565=>x"2e00", 566=>x"3400", 567=>x"3000", 568=>x"2c00",
---- 569=>x"2a00", 570=>x"3200", 571=>x"3200", 572=>x"2b00",
---- 573=>x"2b00", 574=>x"2f00", 575=>x"3600", 576=>x"2b00",
---- 577=>x"2c00", 578=>x"2d00", 579=>x"3100", 580=>x"2c00",
---- 581=>x"2c00", 582=>x"2d00", 583=>x"2e00", 584=>x"3000",
---- 585=>x"2e00", 586=>x"2f00", 587=>x"2f00", 588=>x"2e00",
---- 589=>x"2e00", 590=>x"2d00", 591=>x"2d00", 592=>x"2d00",
---- 593=>x"2a00", 594=>x"2e00", 595=>x"2d00", 596=>x"2800",
---- 597=>x"2600", 598=>x"2c00", 599=>x"2700", 600=>x"2700",
---- 601=>x"2200", 602=>x"2600", 603=>x"2100", 604=>x"2700",
---- 605=>x"2300", 606=>x"2500", 607=>x"2300", 608=>x"2200",
---- 609=>x"2700", 610=>x"2900", 611=>x"2300", 612=>x"1c00",
---- 613=>x"2500", 614=>x"1e00", 615=>x"2f00", 616=>x"1b00",
---- 617=>x"1e00", 618=>x"1900", 619=>x"5d00", 620=>x"1c00",
---- 621=>x"1b00", 622=>x"2900", 623=>x"8000", 624=>x"2300",
---- 625=>x"1a00", 626=>x"4a00", 627=>x"9000", 628=>x"2400",
---- 629=>x"4000", 630=>x"6f00", 631=>x"7d00", 632=>x"5000",
---- 633=>x"8400", 634=>x"7f00", 635=>x"6d00", 636=>x"9f00",
---- 637=>x"a600", 638=>x"9800", 639=>x"8f00", 640=>x"ac00",
---- 641=>x"a500", 642=>x"ab00", 643=>x"ac00", 644=>x"b400",
---- 645=>x"b200", 646=>x"b600", 647=>x"b500", 648=>x"aa00",
---- 649=>x"b900", 650=>x"be00", 651=>x"c000", 652=>x"9a00",
---- 653=>x"a900", 654=>x"af00", 655=>x"b700", 656=>x"8200",
---- 657=>x"7d00", 658=>x"9e00", 659=>x"bf00", 660=>x"6800",
---- 661=>x"7f00", 662=>x"2f00", 663=>x"af00", 664=>x"7b00",
---- 665=>x"b100", 666=>x"cf00", 667=>x"4d00", 668=>x"a300",
---- 669=>x"d100", 670=>x"7500", 671=>x"2800", 672=>x"c300",
---- 673=>x"8b00", 674=>x"2600", 675=>x"2a00", 676=>x"a800",
---- 677=>x"3000", 678=>x"2300", 679=>x"2d00", 680=>x"4a00",
---- 681=>x"2300", 682=>x"2f00", 683=>x"3100", 684=>x"1f00",
---- 685=>x"2700", 686=>x"3100", 687=>x"4400", 688=>x"2c00",
---- 689=>x"2400", 690=>x"4100", 691=>x"5c00", 692=>x"2900",
---- 693=>x"2500", 694=>x"4100", 695=>x"6600", 696=>x"2c00",
---- 697=>x"2900", 698=>x"3000", 699=>x"5200", 700=>x"3500",
---- 701=>x"d600", 702=>x"2a00", 703=>x"4800", 704=>x"2f00",
---- 705=>x"2c00", 706=>x"2b00", 707=>x"3b00", 708=>x"3100",
---- 709=>x"2a00", 710=>x"2a00", 711=>x"3c00", 712=>x"3000",
---- 713=>x"2a00", 714=>x"2a00", 715=>x"3600", 716=>x"3200",
---- 717=>x"2e00", 718=>x"2c00", 719=>x"2b00", 720=>x"3600",
---- 721=>x"2f00", 722=>x"2c00", 723=>x"3100", 724=>x"c100",
---- 725=>x"3500", 726=>x"3300", 727=>x"3700", 728=>x"3b00",
---- 729=>x"3100", 730=>x"3200", 731=>x"3a00", 732=>x"3700",
---- 733=>x"d200", 734=>x"2b00", 735=>x"3700", 736=>x"3b00",
---- 737=>x"3100", 738=>x"3200", 739=>x"3900", 740=>x"3a00",
---- 741=>x"2e00", 742=>x"2d00", 743=>x"3a00", 744=>x"3b00",
---- 745=>x"2e00", 746=>x"2e00", 747=>x"3b00", 748=>x"3900",
---- 749=>x"2d00", 750=>x"3100", 751=>x"3c00", 752=>x"3500",
---- 753=>x"2a00", 754=>x"2f00", 755=>x"3b00", 756=>x"3800",
---- 757=>x"2d00", 758=>x"3200", 759=>x"3e00", 760=>x"3400",
---- 761=>x"2d00", 762=>x"3400", 763=>x"4300", 764=>x"3700",
---- 765=>x"2e00", 766=>x"3100", 767=>x"4200", 768=>x"3100",
---- 769=>x"2d00", 770=>x"3600", 771=>x"4600", 772=>x"2f00",
---- 773=>x"2800", 774=>x"3100", 775=>x"4b00", 776=>x"2f00",
---- 777=>x"2900", 778=>x"3200", 779=>x"4200", 780=>x"2900",
---- 781=>x"2600", 782=>x"3800", 783=>x"4800", 784=>x"3000",
---- 785=>x"2a00", 786=>x"4000", 787=>x"5000", 788=>x"2e00",
---- 789=>x"2d00", 790=>x"3a00", 791=>x"4a00", 792=>x"2c00",
---- 793=>x"2900", 794=>x"3b00", 795=>x"5200", 796=>x"2c00",
---- 797=>x"2c00", 798=>x"3f00", 799=>x"5300", 800=>x"2d00",
---- 801=>x"2700", 802=>x"3d00", 803=>x"5200", 804=>x"2b00",
---- 805=>x"2300", 806=>x"4100", 807=>x"4f00", 808=>x"2b00",
---- 809=>x"2700", 810=>x"4200", 811=>x"5400", 812=>x"3100",
---- 813=>x"2d00", 814=>x"4600", 815=>x"5200", 816=>x"2c00",
---- 817=>x"2a00", 818=>x"bf00", 819=>x"5200", 820=>x"2d00",
---- 821=>x"2900", 822=>x"3c00", 823=>x"4e00", 824=>x"3200",
---- 825=>x"3100", 826=>x"4200", 827=>x"4e00", 828=>x"2f00",
---- 829=>x"2d00", 830=>x"4300", 831=>x"4f00", 832=>x"2a00",
---- 833=>x"2400", 834=>x"4400", 835=>x"4c00", 836=>x"2b00",
---- 837=>x"2500", 838=>x"3c00", 839=>x"4800", 840=>x"2400",
---- 841=>x"2200", 842=>x"3900", 843=>x"4500", 844=>x"2800",
---- 845=>x"2400", 846=>x"3900", 847=>x"4700", 848=>x"2900",
---- 849=>x"2200", 850=>x"3e00", 851=>x"4800", 852=>x"2300",
---- 853=>x"2100", 854=>x"4300", 855=>x"4000", 856=>x"2a00",
---- 857=>x"2600", 858=>x"4700", 859=>x"4800", 860=>x"2500",
---- 861=>x"2b00", 862=>x"5200", 863=>x"4800", 864=>x"1d00",
---- 865=>x"2a00", 866=>x"5300", 867=>x"4500", 868=>x"1b00",
---- 869=>x"3000", 870=>x"4f00", 871=>x"4000", 872=>x"2100",
---- 873=>x"3400", 874=>x"4900", 875=>x"3500", 876=>x"3f00",
---- 877=>x"3a00", 878=>x"4700", 879=>x"3000", 880=>x"3500",
---- 881=>x"3900", 882=>x"3e00", 883=>x"3300", 884=>x"3e00",
---- 885=>x"5300", 886=>x"3f00", 887=>x"2f00", 888=>x"8200",
---- 889=>x"8800", 890=>x"7000", 891=>x"6f00", 892=>x"4c00",
---- 893=>x"5b00", 894=>x"4e00", 895=>x"7c00", 896=>x"4300",
---- 897=>x"3a00", 898=>x"2c00", 899=>x"4100", 900=>x"4200",
---- 901=>x"3d00", 902=>x"3200", 903=>x"4200", 904=>x"3a00",
---- 905=>x"3000", 906=>x"2d00", 907=>x"3f00", 908=>x"3b00",
---- 909=>x"3400", 910=>x"3200", 911=>x"3c00", 912=>x"ca00",
---- 913=>x"2b00", 914=>x"3500", 915=>x"3800", 916=>x"3100",
---- 917=>x"d400", 918=>x"3b00", 919=>x"3900", 920=>x"2700",
---- 921=>x"2b00", 922=>x"3b00", 923=>x"3400", 924=>x"2b00",
---- 925=>x"2e00", 926=>x"2f00", 927=>x"3100", 928=>x"2900",
---- 929=>x"3400", 930=>x"2f00", 931=>x"2f00", 932=>x"3000",
---- 933=>x"3500", 934=>x"2900", 935=>x"2e00", 936=>x"3400",
---- 937=>x"3000", 938=>x"2800", 939=>x"2c00", 940=>x"3100",
---- 941=>x"2800", 942=>x"2700", 943=>x"2900", 944=>x"3200",
---- 945=>x"2a00", 946=>x"2c00", 947=>x"2a00", 948=>x"2f00",
---- 949=>x"2b00", 950=>x"2900", 951=>x"2800", 952=>x"2900",
---- 953=>x"2b00", 954=>x"2600", 955=>x"2a00", 956=>x"2b00",
---- 957=>x"2700", 958=>x"2300", 959=>x"2a00", 960=>x"2500",
---- 961=>x"2300", 962=>x"2500", 963=>x"2f00", 964=>x"2800",
---- 965=>x"2400", 966=>x"2900", 967=>x"2f00", 968=>x"2600",
---- 969=>x"2a00", 970=>x"3100", 971=>x"3200", 972=>x"2300",
---- 973=>x"2500", 974=>x"2a00", 975=>x"3200", 976=>x"2b00",
---- 977=>x"2700", 978=>x"2e00", 979=>x"4000", 980=>x"2f00",
---- 981=>x"2f00", 982=>x"3600", 983=>x"3900", 984=>x"2e00",
---- 985=>x"2d00", 986=>x"2700", 987=>x"2900", 988=>x"2800",
---- 989=>x"2800", 990=>x"2e00", 991=>x"3300", 992=>x"3300",
---- 993=>x"3600", 994=>x"4000", 995=>x"4a00", 996=>x"3400",
---- 997=>x"3a00", 998=>x"4300", 999=>x"5200", 1000=>x"3500",
---- 1001=>x"4800", 1002=>x"5400", 1003=>x"5f00", 1004=>x"4700",
---- 1005=>x"5500", 1006=>x"5d00", 1007=>x"6500", 1008=>x"5300",
---- 1009=>x"5900", 1010=>x"6300", 1011=>x"9500", 1012=>x"5700",
---- 1013=>x"5b00", 1014=>x"6300", 1015=>x"6800", 1016=>x"5700",
---- 1017=>x"5f00", 1018=>x"6800", 1019=>x"6b00", 1020=>x"5900",
---- 1021=>x"5f00", 1022=>x"6700", 1023=>x"6a00"),
----
---- 24 => (0=>x"8700", 1=>x"7900", 2=>x"8700", 3=>x"8700", 4=>x"8700",
---- 5=>x"8600", 6=>x"8700", 7=>x"8800", 8=>x"8700",
---- 9=>x"8500", 10=>x"8700", 11=>x"8700", 12=>x"8400",
---- 13=>x"8600", 14=>x"8500", 15=>x"8400", 16=>x"8500",
---- 17=>x"8500", 18=>x"8300", 19=>x"8400", 20=>x"8700",
---- 21=>x"8400", 22=>x"8200", 23=>x"8400", 24=>x"8200",
---- 25=>x"8500", 26=>x"8200", 27=>x"8300", 28=>x"7f00",
---- 29=>x"8400", 30=>x"8400", 31=>x"8600", 32=>x"8300",
---- 33=>x"8300", 34=>x"8300", 35=>x"8600", 36=>x"8500",
---- 37=>x"8200", 38=>x"8200", 39=>x"8800", 40=>x"8400",
---- 41=>x"8100", 42=>x"8300", 43=>x"8600", 44=>x"8200",
---- 45=>x"8400", 46=>x"8100", 47=>x"8200", 48=>x"8500",
---- 49=>x"8400", 50=>x"8100", 51=>x"8200", 52=>x"8a00",
---- 53=>x"8600", 54=>x"8500", 55=>x"8300", 56=>x"8500",
---- 57=>x"8a00", 58=>x"8700", 59=>x"8300", 60=>x"8600",
---- 61=>x"8400", 62=>x"7b00", 63=>x"8500", 64=>x"8400",
---- 65=>x"8300", 66=>x"8400", 67=>x"8100", 68=>x"8500",
---- 69=>x"8600", 70=>x"8400", 71=>x"8000", 72=>x"7f00",
---- 73=>x"8300", 74=>x"8100", 75=>x"7f00", 76=>x"8400",
---- 77=>x"7f00", 78=>x"7f00", 79=>x"8100", 80=>x"8200",
---- 81=>x"8100", 82=>x"7d00", 83=>x"8000", 84=>x"8100",
---- 85=>x"8000", 86=>x"7e00", 87=>x"8000", 88=>x"8200",
---- 89=>x"8300", 90=>x"7e00", 91=>x"8000", 92=>x"8100",
---- 93=>x"8800", 94=>x"8100", 95=>x"7b00", 96=>x"7d00",
---- 97=>x"7f00", 98=>x"8400", 99=>x"8600", 100=>x"8100",
---- 101=>x"8a00", 102=>x"8e00", 103=>x"9700", 104=>x"8f00",
---- 105=>x"9500", 106=>x"9400", 107=>x"9800", 108=>x"8b00",
---- 109=>x"8e00", 110=>x"9300", 111=>x"9b00", 112=>x"8a00",
---- 113=>x"9200", 114=>x"9400", 115=>x"9200", 116=>x"8b00",
---- 117=>x"9200", 118=>x"8e00", 119=>x"8e00", 120=>x"8900",
---- 121=>x"8200", 122=>x"8400", 123=>x"8300", 124=>x"8700",
---- 125=>x"8100", 126=>x"7e00", 127=>x"8400", 128=>x"8300",
---- 129=>x"8200", 130=>x"7e00", 131=>x"8800", 132=>x"8400",
---- 133=>x"7e00", 134=>x"7f00", 135=>x"8700", 136=>x"7e00",
---- 137=>x"8000", 138=>x"8100", 139=>x"8200", 140=>x"8000",
---- 141=>x"8600", 142=>x"8000", 143=>x"8600", 144=>x"8200",
---- 145=>x"8900", 146=>x"8200", 147=>x"8b00", 148=>x"8800",
---- 149=>x"8700", 150=>x"8600", 151=>x"8c00", 152=>x"8400",
---- 153=>x"8100", 154=>x"8300", 155=>x"8800", 156=>x"8000",
---- 157=>x"8000", 158=>x"7f00", 159=>x"8800", 160=>x"7e00",
---- 161=>x"7900", 162=>x"8100", 163=>x"8500", 164=>x"7f00",
---- 165=>x"7e00", 166=>x"8000", 167=>x"8700", 168=>x"8100",
---- 169=>x"8200", 170=>x"8600", 171=>x"8900", 172=>x"8500",
---- 173=>x"8200", 174=>x"7c00", 175=>x"8e00", 176=>x"8000",
---- 177=>x"8200", 178=>x"8700", 179=>x"8d00", 180=>x"7c00",
---- 181=>x"8700", 182=>x"8b00", 183=>x"8700", 184=>x"8100",
---- 185=>x"8c00", 186=>x"8d00", 187=>x"8900", 188=>x"8800",
---- 189=>x"8a00", 190=>x"7200", 191=>x"8a00", 192=>x"8400",
---- 193=>x"8700", 194=>x"8200", 195=>x"8500", 196=>x"8d00",
---- 197=>x"8900", 198=>x"8700", 199=>x"8c00", 200=>x"8a00",
---- 201=>x"8e00", 202=>x"8900", 203=>x"8700", 204=>x"8f00",
---- 205=>x"8800", 206=>x"8d00", 207=>x"8c00", 208=>x"8d00",
---- 209=>x"8a00", 210=>x"8c00", 211=>x"8e00", 212=>x"8600",
---- 213=>x"8400", 214=>x"8c00", 215=>x"9000", 216=>x"7b00",
---- 217=>x"8c00", 218=>x"8700", 219=>x"8c00", 220=>x"8a00",
---- 221=>x"8200", 222=>x"8c00", 223=>x"8c00", 224=>x"8600",
---- 225=>x"8a00", 226=>x"8a00", 227=>x"8800", 228=>x"8400",
---- 229=>x"8200", 230=>x"8b00", 231=>x"8e00", 232=>x"8400",
---- 233=>x"8b00", 234=>x"8d00", 235=>x"8200", 236=>x"8b00",
---- 237=>x"8b00", 238=>x"7f00", 239=>x"7300", 240=>x"8800",
---- 241=>x"7c00", 242=>x"8100", 243=>x"7e00", 244=>x"8000",
---- 245=>x"7d00", 246=>x"7900", 247=>x"6f00", 248=>x"7a00",
---- 249=>x"7100", 250=>x"6d00", 251=>x"6200", 252=>x"7100",
---- 253=>x"6f00", 254=>x"6b00", 255=>x"8100", 256=>x"6b00",
---- 257=>x"6900", 258=>x"8e00", 259=>x"a300", 260=>x"6c00",
---- 261=>x"8600", 262=>x"9e00", 263=>x"ab00", 264=>x"9500",
---- 265=>x"a300", 266=>x"9600", 267=>x"a400", 268=>x"9c00",
---- 269=>x"a300", 270=>x"a400", 271=>x"9700", 272=>x"9c00",
---- 273=>x"9d00", 274=>x"a100", 275=>x"9400", 276=>x"a400",
---- 277=>x"9400", 278=>x"9300", 279=>x"9200", 280=>x"9a00",
---- 281=>x"9100", 282=>x"8d00", 283=>x"9700", 284=>x"9000",
---- 285=>x"8c00", 286=>x"9b00", 287=>x"9700", 288=>x"8b00",
---- 289=>x"9700", 290=>x"9a00", 291=>x"8000", 292=>x"9000",
---- 293=>x"9700", 294=>x"7f00", 295=>x"8000", 296=>x"8a00",
---- 297=>x"7400", 298=>x"8300", 299=>x"9400", 300=>x"7b00",
---- 301=>x"8900", 302=>x"9800", 303=>x"9200", 304=>x"8500",
---- 305=>x"9600", 306=>x"9800", 307=>x"9600", 308=>x"9400",
---- 309=>x"9100", 310=>x"9300", 311=>x"9800", 312=>x"9500",
---- 313=>x"9400", 314=>x"9100", 315=>x"9b00", 316=>x"9400",
---- 317=>x"9a00", 318=>x"9400", 319=>x"8f00", 320=>x"9a00",
---- 321=>x"9400", 322=>x"6e00", 323=>x"8900", 324=>x"9400",
---- 325=>x"9000", 326=>x"8600", 327=>x"9400", 328=>x"8600",
---- 329=>x"8c00", 330=>x"9000", 331=>x"8f00", 332=>x"8600",
---- 333=>x"9300", 334=>x"8a00", 335=>x"7c00", 336=>x"8f00",
---- 337=>x"8200", 338=>x"7400", 339=>x"8100", 340=>x"7f00",
---- 341=>x"7d00", 342=>x"8400", 343=>x"8600", 344=>x"7b00",
---- 345=>x"8a00", 346=>x"8b00", 347=>x"8500", 348=>x"8200",
---- 349=>x"8500", 350=>x"8d00", 351=>x"9800", 352=>x"8300",
---- 353=>x"8700", 354=>x"8a00", 355=>x"9100", 356=>x"8700",
---- 357=>x"8500", 358=>x"8600", 359=>x"8000", 360=>x"8900",
---- 361=>x"8500", 362=>x"7a00", 363=>x"7f00", 364=>x"8800",
---- 365=>x"8300", 366=>x"7c00", 367=>x"8b00", 368=>x"7c00",
---- 369=>x"7b00", 370=>x"8700", 371=>x"8e00", 372=>x"7a00",
---- 373=>x"8200", 374=>x"8a00", 375=>x"8b00", 376=>x"8400",
---- 377=>x"8f00", 378=>x"8a00", 379=>x"8c00", 380=>x"9300",
---- 381=>x"8a00", 382=>x"8600", 383=>x"8600", 384=>x"8a00",
---- 385=>x"8800", 386=>x"8a00", 387=>x"8600", 388=>x"8300",
---- 389=>x"8800", 390=>x"8900", 391=>x"8d00", 392=>x"6600",
---- 393=>x"6e00", 394=>x"8100", 395=>x"9300", 396=>x"7500",
---- 397=>x"6300", 398=>x"5b00", 399=>x"6d00", 400=>x"7800",
---- 401=>x"6100", 402=>x"6200", 403=>x"5900", 404=>x"6500",
---- 405=>x"3b00", 406=>x"3b00", 407=>x"4500", 408=>x"6d00",
---- 409=>x"6500", 410=>x"5700", 411=>x"5000", 412=>x"6600",
---- 413=>x"5f00", 414=>x"5f00", 415=>x"ae00", 416=>x"3e00",
---- 417=>x"5400", 418=>x"4b00", 419=>x"4d00", 420=>x"4a00",
---- 421=>x"4700", 422=>x"4b00", 423=>x"5700", 424=>x"4800",
---- 425=>x"3a00", 426=>x"3d00", 427=>x"4400", 428=>x"bd00",
---- 429=>x"3900", 430=>x"3500", 431=>x"2e00", 432=>x"3800",
---- 433=>x"3200", 434=>x"2a00", 435=>x"2c00", 436=>x"2c00",
---- 437=>x"2f00", 438=>x"2e00", 439=>x"3000", 440=>x"2e00",
---- 441=>x"2c00", 442=>x"2e00", 443=>x"3200", 444=>x"2b00",
---- 445=>x"2f00", 446=>x"2f00", 447=>x"2e00", 448=>x"2700",
---- 449=>x"3600", 450=>x"3300", 451=>x"3700", 452=>x"2d00",
---- 453=>x"4300", 454=>x"3a00", 455=>x"3900", 456=>x"c100",
---- 457=>x"4600", 458=>x"3100", 459=>x"3900", 460=>x"3e00",
---- 461=>x"3300", 462=>x"3a00", 463=>x"3800", 464=>x"2d00",
---- 465=>x"3300", 466=>x"4000", 467=>x"3000", 468=>x"2f00",
---- 469=>x"4d00", 470=>x"4600", 471=>x"2c00", 472=>x"3d00",
---- 473=>x"5700", 474=>x"3600", 475=>x"2c00", 476=>x"6500",
---- 477=>x"4700", 478=>x"2f00", 479=>x"2600", 480=>x"4900",
---- 481=>x"3a00", 482=>x"2900", 483=>x"2800", 484=>x"4300",
---- 485=>x"3200", 486=>x"2a00", 487=>x"2c00", 488=>x"2c00",
---- 489=>x"2800", 490=>x"2900", 491=>x"2c00", 492=>x"2d00",
---- 493=>x"2b00", 494=>x"3300", 495=>x"3300", 496=>x"3c00",
---- 497=>x"2b00", 498=>x"3600", 499=>x"2e00", 500=>x"4d00",
---- 501=>x"2d00", 502=>x"3600", 503=>x"2700", 504=>x"6000",
---- 505=>x"4200", 506=>x"2c00", 507=>x"2400", 508=>x"6900",
---- 509=>x"5500", 510=>x"2500", 511=>x"2600", 512=>x"5800",
---- 513=>x"6700", 514=>x"3200", 515=>x"2600", 516=>x"3500",
---- 517=>x"6e00", 518=>x"6200", 519=>x"3100", 520=>x"2200",
---- 521=>x"4100", 522=>x"7a00", 523=>x"6e00", 524=>x"2800",
---- 525=>x"2500", 526=>x"4700", 527=>x"7600", 528=>x"d400",
---- 529=>x"2b00", 530=>x"2e00", 531=>x"3e00", 532=>x"2900",
---- 533=>x"2c00", 534=>x"3200", 535=>x"3000", 536=>x"2b00",
---- 537=>x"2b00", 538=>x"3400", 539=>x"3200", 540=>x"2e00",
---- 541=>x"2a00", 542=>x"3300", 543=>x"3100", 544=>x"2b00",
---- 545=>x"2a00", 546=>x"2f00", 547=>x"3100", 548=>x"2e00",
---- 549=>x"2f00", 550=>x"3600", 551=>x"cd00", 552=>x"2f00",
---- 553=>x"3300", 554=>x"3200", 555=>x"2c00", 556=>x"3300",
---- 557=>x"3500", 558=>x"2c00", 559=>x"2600", 560=>x"3200",
---- 561=>x"3400", 562=>x"2f00", 563=>x"2400", 564=>x"2e00",
---- 565=>x"2d00", 566=>x"2900", 567=>x"2500", 568=>x"2c00",
---- 569=>x"2e00", 570=>x"2900", 571=>x"2400", 572=>x"3100",
---- 573=>x"3300", 574=>x"2f00", 575=>x"2700", 576=>x"3400",
---- 577=>x"3000", 578=>x"3000", 579=>x"2400", 580=>x"2e00",
---- 581=>x"2d00", 582=>x"2600", 583=>x"4400", 584=>x"2d00",
---- 585=>x"2a00", 586=>x"2500", 587=>x"7200", 588=>x"2b00",
---- 589=>x"2800", 590=>x"4300", 591=>x"9100", 592=>x"2400",
---- 593=>x"2a00", 594=>x"7700", 595=>x"9300", 596=>x"1e00",
---- 597=>x"4300", 598=>x"9400", 599=>x"7b00", 600=>x"2100",
---- 601=>x"7200", 602=>x"8f00", 603=>x"6b00", 604=>x"3e00",
---- 605=>x"7200", 606=>x"7600", 607=>x"6f00", 608=>x"6300",
---- 609=>x"8f00", 610=>x"6600", 611=>x"7800", 612=>x"8700",
---- 613=>x"8000", 614=>x"6900", 615=>x"9200", 616=>x"9600",
---- 617=>x"6f00", 618=>x"7200", 619=>x"aa00", 620=>x"8100",
---- 621=>x"7000", 622=>x"8400", 623=>x"c100", 624=>x"7300",
---- 625=>x"7300", 626=>x"a600", 627=>x"d300", 628=>x"7600",
---- 629=>x"8800", 630=>x"c900", 631=>x"bd00", 632=>x"6400",
---- 633=>x"8800", 634=>x"ac00", 635=>x"9700", 636=>x"7e00",
---- 637=>x"7d00", 638=>x"9900", 639=>x"b400", 640=>x"ae00",
---- 641=>x"b200", 642=>x"be00", 643=>x"9600", 644=>x"b700",
---- 645=>x"b400", 646=>x"9400", 647=>x"4400", 648=>x"c500",
---- 649=>x"a700", 650=>x"3b00", 651=>x"1f00", 652=>x"be00",
---- 653=>x"6c00", 654=>x"1d00", 655=>x"2600", 656=>x"6b00",
---- 657=>x"2100", 658=>x"2500", 659=>x"2500", 660=>x"2900",
---- 661=>x"2500", 662=>x"2800", 663=>x"2a00", 664=>x"2800",
---- 665=>x"3300", 666=>x"3300", 667=>x"3100", 668=>x"3200",
---- 669=>x"3700", 670=>x"3a00", 671=>x"3500", 672=>x"2c00",
---- 673=>x"2d00", 674=>x"3100", 675=>x"3400", 676=>x"3500",
---- 677=>x"2e00", 678=>x"2f00", 679=>x"3100", 680=>x"3700",
---- 681=>x"3a00", 682=>x"3000", 683=>x"3300", 684=>x"3400",
---- 685=>x"3400", 686=>x"2f00", 687=>x"3500", 688=>x"3800",
---- 689=>x"3200", 690=>x"2a00", 691=>x"3400", 692=>x"3500",
---- 693=>x"2d00", 694=>x"2b00", 695=>x"3300", 696=>x"3300",
---- 697=>x"2b00", 698=>x"2e00", 699=>x"3000", 700=>x"3f00",
---- 701=>x"2700", 702=>x"2f00", 703=>x"2d00", 704=>x"4300",
---- 705=>x"2d00", 706=>x"2f00", 707=>x"3100", 708=>x"3e00",
---- 709=>x"3000", 710=>x"2c00", 711=>x"ca00", 712=>x"c600",
---- 713=>x"3400", 714=>x"2b00", 715=>x"3000", 716=>x"3700",
---- 717=>x"3700", 718=>x"3100", 719=>x"2d00", 720=>x"3500",
---- 721=>x"3600", 722=>x"3400", 723=>x"3100", 724=>x"3600",
---- 725=>x"3100", 726=>x"3500", 727=>x"3700", 728=>x"3600",
---- 729=>x"3300", 730=>x"3500", 731=>x"3e00", 732=>x"3200",
---- 733=>x"3200", 734=>x"3700", 735=>x"c900", 736=>x"3500",
---- 737=>x"3400", 738=>x"3500", 739=>x"3300", 740=>x"3200",
---- 741=>x"3300", 742=>x"3500", 743=>x"3100", 744=>x"3200",
---- 745=>x"3400", 746=>x"3900", 747=>x"3000", 748=>x"3400",
---- 749=>x"cf00", 750=>x"3800", 751=>x"3100", 752=>x"3500",
---- 753=>x"2d00", 754=>x"3500", 755=>x"3800", 756=>x"3300",
---- 757=>x"3100", 758=>x"3100", 759=>x"3a00", 760=>x"3400",
---- 761=>x"3200", 762=>x"3200", 763=>x"3a00", 764=>x"3400",
---- 765=>x"3000", 766=>x"3700", 767=>x"3500", 768=>x"3600",
---- 769=>x"3000", 770=>x"3300", 771=>x"3600", 772=>x"3300",
---- 773=>x"3100", 774=>x"3200", 775=>x"3000", 776=>x"3300",
---- 777=>x"3100", 778=>x"3300", 779=>x"2f00", 780=>x"3000",
---- 781=>x"3000", 782=>x"3000", 783=>x"cf00", 784=>x"2e00",
---- 785=>x"3000", 786=>x"3400", 787=>x"3000", 788=>x"3800",
---- 789=>x"3300", 790=>x"3800", 791=>x"3200", 792=>x"3600",
---- 793=>x"3000", 794=>x"3800", 795=>x"3200", 796=>x"3000",
---- 797=>x"3000", 798=>x"3600", 799=>x"2e00", 800=>x"3000",
---- 801=>x"2f00", 802=>x"3300", 803=>x"2d00", 804=>x"3200",
---- 805=>x"3100", 806=>x"3800", 807=>x"3000", 808=>x"3600",
---- 809=>x"3300", 810=>x"c700", 811=>x"3600", 812=>x"3900",
---- 813=>x"3700", 814=>x"3900", 815=>x"3400", 816=>x"3900",
---- 817=>x"3400", 818=>x"3800", 819=>x"3500", 820=>x"3500",
---- 821=>x"3500", 822=>x"3400", 823=>x"3400", 824=>x"3900",
---- 825=>x"3800", 826=>x"3900", 827=>x"3a00", 828=>x"3c00",
---- 829=>x"3f00", 830=>x"3900", 831=>x"3400", 832=>x"3500",
---- 833=>x"3b00", 834=>x"3600", 835=>x"2e00", 836=>x"3900",
---- 837=>x"3a00", 838=>x"3800", 839=>x"3500", 840=>x"3a00",
---- 841=>x"3e00", 842=>x"3700", 843=>x"3200", 844=>x"3600",
---- 845=>x"4400", 846=>x"3800", 847=>x"3000", 848=>x"3800",
---- 849=>x"4b00", 850=>x"3b00", 851=>x"3100", 852=>x"3700",
---- 853=>x"5800", 854=>x"3800", 855=>x"2f00", 856=>x"3600",
---- 857=>x"6000", 858=>x"3d00", 859=>x"3200", 860=>x"3600",
---- 861=>x"5300", 862=>x"3800", 863=>x"3600", 864=>x"3d00",
---- 865=>x"4e00", 866=>x"3600", 867=>x"3400", 868=>x"3d00",
---- 869=>x"4200", 870=>x"3800", 871=>x"3500", 872=>x"3800",
---- 873=>x"3a00", 874=>x"4300", 875=>x"3700", 876=>x"3b00",
---- 877=>x"3b00", 878=>x"3f00", 879=>x"3500", 880=>x"4400",
---- 881=>x"3500", 882=>x"3c00", 883=>x"3900", 884=>x"3700",
---- 885=>x"3100", 886=>x"4400", 887=>x"5200", 888=>x"6b00",
---- 889=>x"5c00", 890=>x"5b00", 891=>x"4400", 892=>x"9300",
---- 893=>x"6f00", 894=>x"6700", 895=>x"3f00", 896=>x"3f00",
---- 897=>x"3900", 898=>x"6200", 899=>x"7200", 900=>x"3700",
---- 901=>x"3c00", 902=>x"3200", 903=>x"4e00", 904=>x"4000",
---- 905=>x"3800", 906=>x"3200", 907=>x"3100", 908=>x"4000",
---- 909=>x"3400", 910=>x"3300", 911=>x"3200", 912=>x"3300",
---- 913=>x"3100", 914=>x"3300", 915=>x"3300", 916=>x"3400",
---- 917=>x"3100", 918=>x"3300", 919=>x"2e00", 920=>x"2f00",
---- 921=>x"2d00", 922=>x"ce00", 923=>x"2a00", 924=>x"3100",
---- 925=>x"2d00", 926=>x"2800", 927=>x"2800", 928=>x"2f00",
---- 929=>x"2c00", 930=>x"2800", 931=>x"2700", 932=>x"2e00",
---- 933=>x"2c00", 934=>x"2800", 935=>x"2900", 936=>x"2d00",
---- 937=>x"2a00", 938=>x"2e00", 939=>x"2b00", 940=>x"2800",
---- 941=>x"2900", 942=>x"2a00", 943=>x"2d00", 944=>x"2400",
---- 945=>x"2a00", 946=>x"2900", 947=>x"2c00", 948=>x"2600",
---- 949=>x"2b00", 950=>x"2d00", 951=>x"3800", 952=>x"2c00",
---- 953=>x"2a00", 954=>x"3100", 955=>x"4800", 956=>x"2d00",
---- 957=>x"2b00", 958=>x"3c00", 959=>x"4d00", 960=>x"3000",
---- 961=>x"3400", 962=>x"4500", 963=>x"4f00", 964=>x"3300",
---- 965=>x"4300", 966=>x"4b00", 967=>x"4d00", 968=>x"3b00",
---- 969=>x"4a00", 970=>x"4c00", 971=>x"5b00", 972=>x"4600",
---- 973=>x"4e00", 974=>x"5800", 975=>x"6700", 976=>x"4f00",
---- 977=>x"5600", 978=>x"5400", 979=>x"4f00", 980=>x"3600",
---- 981=>x"c400", 982=>x"2b00", 983=>x"2500", 984=>x"2900",
---- 985=>x"2b00", 986=>x"3500", 987=>x"3b00", 988=>x"3f00",
---- 989=>x"4300", 990=>x"5100", 991=>x"5500", 992=>x"5200",
---- 993=>x"5600", 994=>x"5a00", 995=>x"6200", 996=>x"5900",
---- 997=>x"5e00", 998=>x"6a00", 999=>x"7100", 1000=>x"6200",
---- 1001=>x"9500", 1002=>x"7000", 1003=>x"7300", 1004=>x"6900",
---- 1005=>x"6f00", 1006=>x"7100", 1007=>x"7400", 1008=>x"6a00",
---- 1009=>x"6f00", 1010=>x"6f00", 1011=>x"7000", 1012=>x"6800",
---- 1013=>x"7100", 1014=>x"7400", 1015=>x"7300", 1016=>x"7000",
---- 1017=>x"7400", 1018=>x"7600", 1019=>x"7400", 1020=>x"6e00",
---- 1021=>x"6f00", 1022=>x"7400", 1023=>x"7700"),
----
---- 25 => (0=>x"8800", 1=>x"7a00", 2=>x"8800", 3=>x"8500", 4=>x"8800",
---- 5=>x"8600", 6=>x"8800", 7=>x"8500", 8=>x"8700",
---- 9=>x"8600", 10=>x"8800", 11=>x"8500", 12=>x"8500",
---- 13=>x"8400", 14=>x"8400", 15=>x"8400", 16=>x"8400",
---- 17=>x"8200", 18=>x"8300", 19=>x"8200", 20=>x"8300",
---- 21=>x"8300", 22=>x"8400", 23=>x"8000", 24=>x"8300",
---- 25=>x"7d00", 26=>x"8400", 27=>x"8500", 28=>x"8400",
---- 29=>x"8400", 30=>x"8400", 31=>x"8300", 32=>x"8300",
---- 33=>x"8100", 34=>x"8400", 35=>x"8500", 36=>x"8600",
---- 37=>x"8300", 38=>x"8500", 39=>x"8500", 40=>x"8300",
---- 41=>x"8300", 42=>x"8100", 43=>x"8300", 44=>x"8400",
---- 45=>x"7f00", 46=>x"7f00", 47=>x"8400", 48=>x"8200",
---- 49=>x"8100", 50=>x"8000", 51=>x"8000", 52=>x"8300",
---- 53=>x"7f00", 54=>x"7c00", 55=>x"7e00", 56=>x"8000",
---- 57=>x"7b00", 58=>x"7c00", 59=>x"7e00", 60=>x"8200",
---- 61=>x"8000", 62=>x"7d00", 63=>x"7c00", 64=>x"8000",
---- 65=>x"8200", 66=>x"7f00", 67=>x"7c00", 68=>x"7d00",
---- 69=>x"7e00", 70=>x"7d00", 71=>x"7a00", 72=>x"7b00",
---- 73=>x"7f00", 74=>x"7e00", 75=>x"7c00", 76=>x"7e00",
---- 77=>x"7d00", 78=>x"7d00", 79=>x"7c00", 80=>x"7f00",
---- 81=>x"7d00", 82=>x"7f00", 83=>x"7c00", 84=>x"7f00",
---- 85=>x"7d00", 86=>x"8500", 87=>x"8100", 88=>x"7e00",
---- 89=>x"7d00", 90=>x"7f00", 91=>x"8100", 92=>x"7d00",
---- 93=>x"7b00", 94=>x"7e00", 95=>x"7e00", 96=>x"8500",
---- 97=>x"8500", 98=>x"9200", 99=>x"7400", 100=>x"9500",
---- 101=>x"9600", 102=>x"9900", 103=>x"9b00", 104=>x"9500",
---- 105=>x"8c00", 106=>x"9200", 107=>x"9400", 108=>x"8f00",
---- 109=>x"8c00", 110=>x"8a00", 111=>x"9100", 112=>x"9100",
---- 113=>x"9100", 114=>x"9000", 115=>x"9700", 116=>x"8b00",
---- 117=>x"9300", 118=>x"9900", 119=>x"9600", 120=>x"8d00",
---- 121=>x"9500", 122=>x"8d00", 123=>x"9300", 124=>x"8f00",
---- 125=>x"8600", 126=>x"8600", 127=>x"8e00", 128=>x"7400",
---- 129=>x"8a00", 130=>x"8900", 131=>x"8d00", 132=>x"8700",
---- 133=>x"8400", 134=>x"8b00", 135=>x"8700", 136=>x"8500",
---- 137=>x"8900", 138=>x"8a00", 139=>x"8400", 140=>x"8c00",
---- 141=>x"8900", 142=>x"8100", 143=>x"8100", 144=>x"8c00",
---- 145=>x"8200", 146=>x"7b00", 147=>x"8700", 148=>x"8100",
---- 149=>x"8200", 150=>x"8b00", 151=>x"8b00", 152=>x"8d00",
---- 153=>x"8b00", 154=>x"8d00", 155=>x"8800", 156=>x"8700",
---- 157=>x"8400", 158=>x"8900", 159=>x"8100", 160=>x"8300",
---- 161=>x"8600", 162=>x"8800", 163=>x"8a00", 164=>x"8200",
---- 165=>x"8100", 166=>x"8200", 167=>x"8400", 168=>x"8a00",
---- 169=>x"8700", 170=>x"7600", 171=>x"8700", 172=>x"8900",
---- 173=>x"8700", 174=>x"8c00", 175=>x"8700", 176=>x"8800",
---- 177=>x"8200", 178=>x"8900", 179=>x"8800", 180=>x"8100",
---- 181=>x"7400", 182=>x"8b00", 183=>x"8b00", 184=>x"9100",
---- 185=>x"8b00", 186=>x"8c00", 187=>x"8c00", 188=>x"8a00",
---- 189=>x"9000", 190=>x"9000", 191=>x"9000", 192=>x"8f00",
---- 193=>x"8c00", 194=>x"9000", 195=>x"9100", 196=>x"8200",
---- 197=>x"9000", 198=>x"8800", 199=>x"8e00", 200=>x"7100",
---- 201=>x"8f00", 202=>x"8c00", 203=>x"8d00", 204=>x"8600",
---- 205=>x"8f00", 206=>x"8800", 207=>x"8c00", 208=>x"8e00",
---- 209=>x"8700", 210=>x"8b00", 211=>x"8900", 212=>x"9100",
---- 213=>x"8b00", 214=>x"9000", 215=>x"8b00", 216=>x"8f00",
---- 217=>x"8900", 218=>x"8c00", 219=>x"8500", 220=>x"8900",
---- 221=>x"8d00", 222=>x"8300", 223=>x"8100", 224=>x"9000",
---- 225=>x"8800", 226=>x"8600", 227=>x"7c00", 228=>x"8a00",
---- 229=>x"7700", 230=>x"7900", 231=>x"7f00", 232=>x"7300",
---- 233=>x"7100", 234=>x"7900", 235=>x"7200", 236=>x"7600",
---- 237=>x"7100", 238=>x"6400", 239=>x"7200", 240=>x"7100",
---- 241=>x"6500", 242=>x"7400", 243=>x"9d00", 244=>x"6800",
---- 245=>x"7e00", 246=>x"9f00", 247=>x"a300", 248=>x"8100",
---- 249=>x"a700", 250=>x"ac00", 251=>x"a800", 252=>x"a100",
---- 253=>x"ab00", 254=>x"ae00", 255=>x"b600", 256=>x"9f00",
---- 257=>x"ac00", 258=>x"b200", 259=>x"ad00", 260=>x"a600",
---- 261=>x"a700", 262=>x"a400", 263=>x"a000", 264=>x"b300",
---- 265=>x"9d00", 266=>x"9000", 267=>x"9900", 268=>x"9600",
---- 269=>x"9e00", 270=>x"9200", 271=>x"9600", 272=>x"8900",
---- 273=>x"8d00", 274=>x"a600", 275=>x"a000", 276=>x"9500",
---- 277=>x"9a00", 278=>x"9000", 279=>x"8b00", 280=>x"a600",
---- 281=>x"8d00", 282=>x"7e00", 283=>x"9900", 284=>x"8500",
---- 285=>x"8200", 286=>x"9b00", 287=>x"a000", 288=>x"8200",
---- 289=>x"9900", 290=>x"a000", 291=>x"9d00", 292=>x"9800",
---- 293=>x"9500", 294=>x"9400", 295=>x"a200", 296=>x"9200",
---- 297=>x"9600", 298=>x"9700", 299=>x"9800", 300=>x"9300",
---- 301=>x"9200", 302=>x"5f00", 303=>x"9500", 304=>x"9800",
---- 305=>x"9b00", 306=>x"9d00", 307=>x"8900", 308=>x"9a00",
---- 309=>x"9a00", 310=>x"8e00", 311=>x"8500", 312=>x"9700",
---- 313=>x"9500", 314=>x"9000", 315=>x"8f00", 316=>x"8f00",
---- 317=>x"8c00", 318=>x"9a00", 319=>x"9e00", 320=>x"8d00",
---- 321=>x"9800", 322=>x"9500", 323=>x"9800", 324=>x"8a00",
---- 325=>x"8f00", 326=>x"8900", 327=>x"8a00", 328=>x"8700",
---- 329=>x"8300", 330=>x"9100", 331=>x"9200", 332=>x"8200",
---- 333=>x"9200", 334=>x"9800", 335=>x"9900", 336=>x"8f00",
---- 337=>x"9600", 338=>x"9300", 339=>x"9800", 340=>x"9600",
---- 341=>x"9b00", 342=>x"9100", 343=>x"8000", 344=>x"8e00",
---- 345=>x"9700", 346=>x"8100", 347=>x"8900", 348=>x"8600",
---- 349=>x"7d00", 350=>x"8800", 351=>x"9500", 352=>x"8200",
---- 353=>x"8000", 354=>x"9300", 355=>x"9400", 356=>x"8100",
---- 357=>x"9300", 358=>x"8b00", 359=>x"8d00", 360=>x"8e00",
---- 361=>x"9600", 362=>x"8d00", 363=>x"8b00", 364=>x"8f00",
---- 365=>x"8c00", 366=>x"8c00", 367=>x"7100", 368=>x"8900",
---- 369=>x"8900", 370=>x"8f00", 371=>x"7400", 372=>x"8a00",
---- 373=>x"8300", 374=>x"7700", 375=>x"6c00", 376=>x"8800",
---- 377=>x"7100", 378=>x"6900", 379=>x"7c00", 380=>x"8500",
---- 381=>x"6300", 382=>x"7200", 383=>x"8b00", 384=>x"8900",
---- 385=>x"6600", 386=>x"7400", 387=>x"8b00", 388=>x"9200",
---- 389=>x"6c00", 390=>x"7200", 391=>x"8700", 392=>x"9100",
---- 393=>x"6d00", 394=>x"9d00", 395=>x"5d00", 396=>x"7f00",
---- 397=>x"9000", 398=>x"4800", 399=>x"3a00", 400=>x"4a00",
---- 401=>x"5600", 402=>x"4c00", 403=>x"4400", 404=>x"4800",
---- 405=>x"4f00", 406=>x"4a00", 407=>x"4e00", 408=>x"4b00",
---- 409=>x"3d00", 410=>x"4300", 411=>x"5d00", 412=>x"4400",
---- 413=>x"4800", 414=>x"5f00", 415=>x"5e00", 416=>x"5500",
---- 417=>x"5d00", 418=>x"6500", 419=>x"5300", 420=>x"4e00",
---- 421=>x"6300", 422=>x"5b00", 423=>x"4400", 424=>x"4600",
---- 425=>x"5e00", 426=>x"5400", 427=>x"4800", 428=>x"4200",
---- 429=>x"5600", 430=>x"4c00", 431=>x"4300", 432=>x"3200",
---- 433=>x"4900", 434=>x"4d00", 435=>x"4400", 436=>x"2d00",
---- 437=>x"4900", 438=>x"5900", 439=>x"3f00", 440=>x"2e00",
---- 441=>x"3700", 442=>x"5900", 443=>x"4b00", 444=>x"3100",
---- 445=>x"3100", 446=>x"3c00", 447=>x"5300", 448=>x"3300",
---- 449=>x"2f00", 450=>x"2e00", 451=>x"4100", 452=>x"3000",
---- 453=>x"2e00", 454=>x"3400", 455=>x"3300", 456=>x"2e00",
---- 457=>x"3400", 458=>x"3b00", 459=>x"3000", 460=>x"2c00",
---- 461=>x"3600", 462=>x"3800", 463=>x"2f00", 464=>x"cd00",
---- 465=>x"3900", 466=>x"3400", 467=>x"3200", 468=>x"3400",
---- 469=>x"3700", 470=>x"2a00", 471=>x"3800", 472=>x"3300",
---- 473=>x"3300", 474=>x"2700", 475=>x"4300", 476=>x"3600",
---- 477=>x"3100", 478=>x"2600", 479=>x"5000", 480=>x"3700",
---- 481=>x"2d00", 482=>x"2800", 483=>x"5a00", 484=>x"3800",
---- 485=>x"3000", 486=>x"3400", 487=>x"5800", 488=>x"3200",
---- 489=>x"3100", 490=>x"3800", 491=>x"4300", 492=>x"2f00",
---- 493=>x"3800", 494=>x"3e00", 495=>x"4000", 496=>x"2b00",
---- 497=>x"3000", 498=>x"4600", 499=>x"6200", 500=>x"2800",
---- 501=>x"2200", 502=>x"2700", 503=>x"5200", 504=>x"2900",
---- 505=>x"2800", 506=>x"2700", 507=>x"3300", 508=>x"2700",
---- 509=>x"2e00", 510=>x"2b00", 511=>x"2800", 512=>x"2a00",
---- 513=>x"d100", 514=>x"2e00", 515=>x"2c00", 516=>x"2500",
---- 517=>x"2c00", 518=>x"2f00", 519=>x"3000", 520=>x"4300",
---- 521=>x"2200", 522=>x"2300", 523=>x"2d00", 524=>x"6900",
---- 525=>x"4c00", 526=>x"3500", 527=>x"2700", 528=>x"3500",
---- 529=>x"4400", 530=>x"5800", 531=>x"3600", 532=>x"2700",
---- 533=>x"2b00", 534=>x"3900", 535=>x"2e00", 536=>x"2700",
---- 537=>x"2c00", 538=>x"2a00", 539=>x"2400", 540=>x"2800",
---- 541=>x"2500", 542=>x"2600", 543=>x"2c00", 544=>x"2600",
---- 545=>x"2700", 546=>x"2200", 547=>x"2c00", 548=>x"2700",
---- 549=>x"2500", 550=>x"2300", 551=>x"2800", 552=>x"2300",
---- 553=>x"2300", 554=>x"1b00", 555=>x"4200", 556=>x"2400",
---- 557=>x"2000", 558=>x"2600", 559=>x"7a00", 560=>x"2100",
---- 561=>x"1c00", 562=>x"5700", 563=>x"9900", 564=>x"1f00",
---- 565=>x"2f00", 566=>x"8a00", 567=>x"8700", 568=>x"2200",
---- 569=>x"6200", 570=>x"9800", 571=>x"6600", 572=>x"3c00",
---- 573=>x"9000", 574=>x"7700", 575=>x"6200", 576=>x"6f00",
---- 577=>x"9400", 578=>x"6200", 579=>x"8400", 580=>x"9800",
---- 581=>x"7400", 582=>x"6400", 583=>x"a300", 584=>x"9600",
---- 585=>x"6400", 586=>x"7e00", 587=>x"b600", 588=>x"7d00",
---- 589=>x"6f00", 590=>x"9500", 591=>x"b500", 592=>x"6d00",
---- 593=>x"8200", 594=>x"bb00", 595=>x"b700", 596=>x"6f00",
---- 597=>x"a200", 598=>x"c600", 599=>x"be00", 600=>x"7b00",
---- 601=>x"bc00", 602=>x"bd00", 603=>x"c200", 604=>x"9a00",
---- 605=>x"c200", 606=>x"c000", 607=>x"cb00", 608=>x"b800",
---- 609=>x"c800", 610=>x"c700", 611=>x"da00", 612=>x"ca00",
---- 613=>x"ca00", 614=>x"d000", 615=>x"c000", 616=>x"cb00",
---- 617=>x"cb00", 618=>x"3100", 619=>x"5b00", 620=>x"ca00",
---- 621=>x"d500", 622=>x"8200", 623=>x"1d00", 624=>x"d400",
---- 625=>x"a700", 626=>x"2800", 627=>x"2400", 628=>x"a700",
---- 629=>x"5300", 630=>x"1900", 631=>x"2500", 632=>x"9200",
---- 633=>x"4f00", 634=>x"2700", 635=>x"2100", 636=>x"8b00",
---- 637=>x"3500", 638=>x"2100", 639=>x"2700", 640=>x"4a00",
---- 641=>x"2500", 642=>x"2200", 643=>x"2700", 644=>x"2700",
---- 645=>x"2100", 646=>x"2200", 647=>x"2700", 648=>x"2700",
---- 649=>x"2400", 650=>x"2500", 651=>x"2b00", 652=>x"2b00",
---- 653=>x"2b00", 654=>x"d300", 655=>x"2c00", 656=>x"3a00",
---- 657=>x"4900", 658=>x"3f00", 659=>x"2f00", 660=>x"3400",
---- 661=>x"4100", 662=>x"3c00", 663=>x"3000", 664=>x"3400",
---- 665=>x"3700", 666=>x"3a00", 667=>x"3500", 668=>x"3700",
---- 669=>x"3a00", 670=>x"3e00", 671=>x"3900", 672=>x"3300",
---- 673=>x"3800", 674=>x"4100", 675=>x"3f00", 676=>x"2d00",
---- 677=>x"3300", 678=>x"4300", 679=>x"3d00", 680=>x"2e00",
---- 681=>x"3700", 682=>x"4300", 683=>x"4400", 684=>x"3300",
---- 685=>x"3400", 686=>x"4300", 687=>x"4a00", 688=>x"3200",
---- 689=>x"3300", 690=>x"3f00", 691=>x"4e00", 692=>x"3600",
---- 693=>x"3700", 694=>x"4400", 695=>x"4b00", 696=>x"3400",
---- 697=>x"3c00", 698=>x"ba00", 699=>x"4500", 700=>x"3200",
---- 701=>x"3b00", 702=>x"3a00", 703=>x"4400", 704=>x"3500",
---- 705=>x"3900", 706=>x"3a00", 707=>x"3e00", 708=>x"3b00",
---- 709=>x"3c00", 710=>x"c200", 711=>x"3900", 712=>x"3d00",
---- 713=>x"3800", 714=>x"3d00", 715=>x"3900", 716=>x"3400",
---- 717=>x"3900", 718=>x"3c00", 719=>x"3d00", 720=>x"3100",
---- 721=>x"4000", 722=>x"3a00", 723=>x"3b00", 724=>x"3500",
---- 725=>x"3800", 726=>x"3f00", 727=>x"3b00", 728=>x"3e00",
---- 729=>x"3800", 730=>x"4200", 731=>x"3d00", 732=>x"3c00",
---- 733=>x"3f00", 734=>x"3700", 735=>x"3e00", 736=>x"3900",
---- 737=>x"3b00", 738=>x"3900", 739=>x"3900", 740=>x"3200",
---- 741=>x"3800", 742=>x"c300", 743=>x"3800", 744=>x"2f00",
---- 745=>x"2f00", 746=>x"3a00", 747=>x"3800", 748=>x"2b00",
---- 749=>x"2f00", 750=>x"3300", 751=>x"3900", 752=>x"2e00",
---- 753=>x"3200", 754=>x"3100", 755=>x"cc00", 756=>x"3100",
---- 757=>x"2d00", 758=>x"3100", 759=>x"3100", 760=>x"3800",
---- 761=>x"2d00", 762=>x"3000", 763=>x"2f00", 764=>x"3700",
---- 765=>x"3000", 766=>x"3200", 767=>x"3400", 768=>x"3a00",
---- 769=>x"3400", 770=>x"3100", 771=>x"3500", 772=>x"3a00",
---- 773=>x"3200", 774=>x"2f00", 775=>x"3400", 776=>x"3600",
---- 777=>x"3500", 778=>x"2e00", 779=>x"3400", 780=>x"3500",
---- 781=>x"3500", 782=>x"2f00", 783=>x"3200", 784=>x"3300",
---- 785=>x"3900", 786=>x"cd00", 787=>x"2f00", 788=>x"2e00",
---- 789=>x"3200", 790=>x"3600", 791=>x"3400", 792=>x"d100",
---- 793=>x"2f00", 794=>x"3900", 795=>x"3600", 796=>x"3000",
---- 797=>x"2c00", 798=>x"3600", 799=>x"3700", 800=>x"3000",
---- 801=>x"2d00", 802=>x"3700", 803=>x"3900", 804=>x"3000",
---- 805=>x"2b00", 806=>x"3400", 807=>x"3b00", 808=>x"3500",
---- 809=>x"2f00", 810=>x"3300", 811=>x"3700", 812=>x"3100",
---- 813=>x"3000", 814=>x"3500", 815=>x"3800", 816=>x"3500",
---- 817=>x"2f00", 818=>x"3200", 819=>x"3500", 820=>x"3700",
---- 821=>x"3300", 822=>x"3500", 823=>x"3400", 824=>x"3900",
---- 825=>x"3500", 826=>x"3700", 827=>x"3a00", 828=>x"3500",
---- 829=>x"3000", 830=>x"3100", 831=>x"3900", 832=>x"3300",
---- 833=>x"2b00", 834=>x"3200", 835=>x"3400", 836=>x"3400",
---- 837=>x"2f00", 838=>x"3200", 839=>x"3400", 840=>x"3200",
---- 841=>x"2b00", 842=>x"2d00", 843=>x"3100", 844=>x"3000",
---- 845=>x"2b00", 846=>x"3200", 847=>x"cd00", 848=>x"3300",
---- 849=>x"2e00", 850=>x"3400", 851=>x"3200", 852=>x"3100",
---- 853=>x"2b00", 854=>x"3200", 855=>x"3400", 856=>x"3200",
---- 857=>x"3300", 858=>x"3200", 859=>x"2e00", 860=>x"3700",
---- 861=>x"3300", 862=>x"3300", 863=>x"3300", 864=>x"3300",
---- 865=>x"3100", 866=>x"2f00", 867=>x"3300", 868=>x"3800",
---- 869=>x"3d00", 870=>x"2f00", 871=>x"3200", 872=>x"3700",
---- 873=>x"4000", 874=>x"3200", 875=>x"3700", 876=>x"3400",
---- 877=>x"3900", 878=>x"3200", 879=>x"3c00", 880=>x"3800",
---- 881=>x"3a00", 882=>x"2f00", 883=>x"3b00", 884=>x"3d00",
---- 885=>x"3500", 886=>x"3600", 887=>x"3e00", 888=>x"3b00",
---- 889=>x"3200", 890=>x"3000", 891=>x"3700", 892=>x"3e00",
---- 893=>x"3400", 894=>x"3800", 895=>x"3800", 896=>x"4700",
---- 897=>x"3400", 898=>x"3400", 899=>x"3400", 900=>x"4900",
---- 901=>x"3600", 902=>x"2e00", 903=>x"2c00", 904=>x"3900",
---- 905=>x"3700", 906=>x"2f00", 907=>x"2e00", 908=>x"3500",
---- 909=>x"3400", 910=>x"2a00", 911=>x"2e00", 912=>x"2e00",
---- 913=>x"3000", 914=>x"2e00", 915=>x"2e00", 916=>x"2c00",
---- 917=>x"2f00", 918=>x"2e00", 919=>x"3100", 920=>x"2900",
---- 921=>x"3100", 922=>x"3300", 923=>x"3300", 924=>x"2b00",
---- 925=>x"3200", 926=>x"3c00", 927=>x"4100", 928=>x"2f00",
---- 929=>x"3200", 930=>x"4500", 931=>x"4800", 932=>x"3300",
---- 933=>x"3600", 934=>x"4400", 935=>x"4f00", 936=>x"3500",
---- 937=>x"3b00", 938=>x"4a00", 939=>x"5100", 940=>x"3800",
---- 941=>x"4000", 942=>x"5300", 943=>x"5a00", 944=>x"3c00",
---- 945=>x"4800", 946=>x"5600", 947=>x"6100", 948=>x"4800",
---- 949=>x"4c00", 950=>x"5c00", 951=>x"6800", 952=>x"4e00",
---- 953=>x"5400", 954=>x"6300", 955=>x"6f00", 956=>x"4b00",
---- 957=>x"5800", 958=>x"6b00", 959=>x"7300", 960=>x"5000",
---- 961=>x"6200", 962=>x"6d00", 963=>x"7800", 964=>x"5e00",
---- 965=>x"6600", 966=>x"6e00", 967=>x"7900", 968=>x"6700",
---- 969=>x"6800", 970=>x"7300", 971=>x"7500", 972=>x"6900",
---- 973=>x"6300", 974=>x"5300", 975=>x"4000", 976=>x"4000",
---- 977=>x"3800", 978=>x"2500", 979=>x"2500", 980=>x"2800",
---- 981=>x"2d00", 982=>x"3900", 983=>x"4d00", 984=>x"4600",
---- 985=>x"5100", 986=>x"5900", 987=>x"6200", 988=>x"5c00",
---- 989=>x"5a00", 990=>x"6500", 991=>x"6a00", 992=>x"6500",
---- 993=>x"6a00", 994=>x"7200", 995=>x"7600", 996=>x"7000",
---- 997=>x"7200", 998=>x"7200", 999=>x"7500", 1000=>x"7400",
---- 1001=>x"7200", 1002=>x"7300", 1003=>x"7600", 1004=>x"7600",
---- 1005=>x"7400", 1006=>x"7400", 1007=>x"7500", 1008=>x"7900",
---- 1009=>x"7700", 1010=>x"7700", 1011=>x"7600", 1012=>x"7800",
---- 1013=>x"7900", 1014=>x"7900", 1015=>x"7800", 1016=>x"7700",
---- 1017=>x"7a00", 1018=>x"7800", 1019=>x"7a00", 1020=>x"7800",
---- 1021=>x"7b00", 1022=>x"7900", 1023=>x"7c00"),
----
---- 26 => (0=>x"8700", 1=>x"8600", 2=>x"8700", 3=>x"8200", 4=>x"8700",
---- 5=>x"8600", 6=>x"8700", 7=>x"7d00", 8=>x"8600",
---- 9=>x"8600", 10=>x"8500", 11=>x"7e00", 12=>x"8600",
---- 13=>x"8500", 14=>x"8700", 15=>x"7e00", 16=>x"8300",
---- 17=>x"8200", 18=>x"8500", 19=>x"8500", 20=>x"8100",
---- 21=>x"8500", 22=>x"8200", 23=>x"8100", 24=>x"8600",
---- 25=>x"8500", 26=>x"8400", 27=>x"8400", 28=>x"8200",
---- 29=>x"8300", 30=>x"8300", 31=>x"8300", 32=>x"8600",
---- 33=>x"8500", 34=>x"8600", 35=>x"8200", 36=>x"8300",
---- 37=>x"8300", 38=>x"8500", 39=>x"8400", 40=>x"8700",
---- 41=>x"8200", 42=>x"8100", 43=>x"8200", 44=>x"8500",
---- 45=>x"7e00", 46=>x"8100", 47=>x"8100", 48=>x"7e00",
---- 49=>x"7f00", 50=>x"8000", 51=>x"7e00", 52=>x"7e00",
---- 53=>x"7d00", 54=>x"7c00", 55=>x"7e00", 56=>x"7c00",
---- 57=>x"7900", 58=>x"7b00", 59=>x"7b00", 60=>x"7b00",
---- 61=>x"7900", 62=>x"7b00", 63=>x"8500", 64=>x"7b00",
---- 65=>x"7a00", 66=>x"7c00", 67=>x"7900", 68=>x"7b00",
---- 69=>x"7d00", 70=>x"7900", 71=>x"7600", 72=>x"7c00",
---- 73=>x"7d00", 74=>x"7c00", 75=>x"7900", 76=>x"7c00",
---- 77=>x"7b00", 78=>x"7800", 79=>x"7a00", 80=>x"8100",
---- 81=>x"7b00", 82=>x"7a00", 83=>x"7c00", 84=>x"7e00",
---- 85=>x"7d00", 86=>x"7f00", 87=>x"7d00", 88=>x"7f00",
---- 89=>x"7c00", 90=>x"7a00", 91=>x"7b00", 92=>x"8700",
---- 93=>x"8a00", 94=>x"8800", 95=>x"8700", 96=>x"9700",
---- 97=>x"9100", 98=>x"9100", 99=>x"6900", 100=>x"9300",
---- 101=>x"9100", 102=>x"9a00", 103=>x"a800", 104=>x"9200",
---- 105=>x"9900", 106=>x"a400", 107=>x"ac00", 108=>x"9600",
---- 109=>x"9800", 110=>x"9d00", 111=>x"a800", 112=>x"9600",
---- 113=>x"9300", 114=>x"9800", 115=>x"9900", 116=>x"9500",
---- 117=>x"9300", 118=>x"9700", 119=>x"9c00", 120=>x"9700",
---- 121=>x"9500", 122=>x"9900", 123=>x"9900", 124=>x"9500",
---- 125=>x"9b00", 126=>x"9800", 127=>x"9600", 128=>x"9300",
---- 129=>x"9500", 130=>x"9000", 131=>x"9900", 132=>x"8c00",
---- 133=>x"9000", 134=>x"8f00", 135=>x"9400", 136=>x"8c00",
---- 137=>x"8c00", 138=>x"9200", 139=>x"8e00", 140=>x"8900",
---- 141=>x"8600", 142=>x"8200", 143=>x"8f00", 144=>x"8d00",
---- 145=>x"8d00", 146=>x"8c00", 147=>x"9100", 148=>x"8600",
---- 149=>x"8e00", 150=>x"8a00", 151=>x"8e00", 152=>x"8500",
---- 153=>x"8800", 154=>x"8500", 155=>x"8900", 156=>x"7400",
---- 157=>x"8f00", 158=>x"8400", 159=>x"8f00", 160=>x"8100",
---- 161=>x"7900", 162=>x"8700", 163=>x"9500", 164=>x"8700",
---- 165=>x"8200", 166=>x"8d00", 167=>x"8f00", 168=>x"8200",
---- 169=>x"8a00", 170=>x"8600", 171=>x"8c00", 172=>x"8800",
---- 173=>x"8400", 174=>x"8f00", 175=>x"8c00", 176=>x"8500",
---- 177=>x"9100", 178=>x"8b00", 179=>x"8d00", 180=>x"8d00",
---- 181=>x"8f00", 182=>x"8d00", 183=>x"8e00", 184=>x"8b00",
---- 185=>x"9300", 186=>x"9300", 187=>x"9100", 188=>x"9400",
---- 189=>x"9300", 190=>x"8f00", 191=>x"8100", 192=>x"9500",
---- 193=>x"9000", 194=>x"8600", 195=>x"8a00", 196=>x"9200",
---- 197=>x"8700", 198=>x"8e00", 199=>x"8b00", 200=>x"8800",
---- 201=>x"8c00", 202=>x"8400", 203=>x"8400", 204=>x"8700",
---- 205=>x"8500", 206=>x"8700", 207=>x"8100", 208=>x"8500",
---- 209=>x"8a00", 210=>x"8900", 211=>x"8500", 212=>x"8400",
---- 213=>x"8500", 214=>x"8200", 215=>x"7d00", 216=>x"8500",
---- 217=>x"8200", 218=>x"7800", 219=>x"8200", 220=>x"8300",
---- 221=>x"8000", 222=>x"7900", 223=>x"6f00", 224=>x"7e00",
---- 225=>x"7b00", 226=>x"6900", 227=>x"6e00", 228=>x"7900",
---- 229=>x"6a00", 230=>x"7500", 231=>x"9700", 232=>x"6e00",
---- 233=>x"7f00", 234=>x"a600", 235=>x"b300", 236=>x"9000",
---- 237=>x"a500", 238=>x"a500", 239=>x"b400", 240=>x"ad00",
---- 241=>x"ab00", 242=>x"ae00", 243=>x"bd00", 244=>x"af00",
---- 245=>x"b700", 246=>x"b500", 247=>x"b400", 248=>x"b500",
---- 249=>x"b800", 250=>x"a900", 251=>x"a900", 252=>x"af00",
---- 253=>x"a800", 254=>x"a400", 255=>x"a200", 256=>x"a900",
---- 257=>x"a100", 258=>x"9800", 259=>x"a700", 260=>x"9e00",
---- 261=>x"a600", 262=>x"ac00", 263=>x"a700", 264=>x"a300",
---- 265=>x"b300", 266=>x"aa00", 267=>x"9500", 268=>x"ae00",
---- 269=>x"9e00", 270=>x"9500", 271=>x"ac00", 272=>x"8600",
---- 273=>x"9500", 274=>x"ad00", 275=>x"b100", 276=>x"9600",
---- 277=>x"9f00", 278=>x"a900", 279=>x"ae00", 280=>x"a700",
---- 281=>x"a700", 282=>x"9800", 283=>x"a400", 284=>x"a000",
---- 285=>x"a200", 286=>x"a400", 287=>x"a700", 288=>x"9800",
---- 289=>x"a300", 290=>x"ae00", 291=>x"a200", 292=>x"a600",
---- 293=>x"a300", 294=>x"a100", 295=>x"a000", 296=>x"ae00",
---- 297=>x"9900", 298=>x"9400", 299=>x"9e00", 300=>x"8800",
---- 301=>x"9d00", 302=>x"9400", 303=>x"9a00", 304=>x"8900",
---- 305=>x"8d00", 306=>x"9a00", 307=>x"a100", 308=>x"8e00",
---- 309=>x"9300", 310=>x"9400", 311=>x"a200", 312=>x"9d00",
---- 313=>x"a200", 314=>x"9200", 315=>x"8800", 316=>x"9600",
---- 317=>x"9100", 318=>x"9100", 319=>x"8e00", 320=>x"8a00",
---- 321=>x"9900", 322=>x"9d00", 323=>x"9b00", 324=>x"9e00",
---- 325=>x"9d00", 326=>x"a000", 327=>x"9100", 328=>x"9900",
---- 329=>x"9500", 330=>x"8a00", 331=>x"8e00", 332=>x"9100",
---- 333=>x"8600", 334=>x"8900", 335=>x"9900", 336=>x"8700",
---- 337=>x"7200", 338=>x"9e00", 339=>x"a000", 340=>x"8200",
---- 341=>x"9400", 342=>x"9c00", 343=>x"a400", 344=>x"9500",
---- 345=>x"9100", 346=>x"9700", 347=>x"9a00", 348=>x"9d00",
---- 349=>x"9a00", 350=>x"9300", 351=>x"8400", 352=>x"9200",
---- 353=>x"9900", 354=>x"9200", 355=>x"6c00", 356=>x"9800",
---- 357=>x"8d00", 358=>x"7400", 359=>x"8300", 360=>x"8b00",
---- 361=>x"7300", 362=>x"8e00", 363=>x"8b00", 364=>x"6d00",
---- 365=>x"6800", 366=>x"8b00", 367=>x"8f00", 368=>x"6d00",
---- 369=>x"8400", 370=>x"8300", 371=>x"8300", 372=>x"8400",
---- 373=>x"8700", 374=>x"8500", 375=>x"7a00", 376=>x"8300",
---- 377=>x"8900", 378=>x"8500", 379=>x"7800", 380=>x"8500",
---- 381=>x"8200", 382=>x"7500", 383=>x"6100", 384=>x"7e00",
---- 385=>x"6600", 386=>x"5000", 387=>x"4000", 388=>x"5700",
---- 389=>x"4700", 390=>x"3800", 391=>x"3a00", 392=>x"4000",
---- 393=>x"3c00", 394=>x"4200", 395=>x"5f00", 396=>x"4200",
---- 397=>x"4f00", 398=>x"5300", 399=>x"4900", 400=>x"4500",
---- 401=>x"5800", 402=>x"4f00", 403=>x"4600", 404=>x"5600",
---- 405=>x"5700", 406=>x"4200", 407=>x"3f00", 408=>x"4900",
---- 409=>x"3600", 410=>x"3100", 411=>x"2d00", 412=>x"3e00",
---- 413=>x"2e00", 414=>x"2700", 415=>x"2500", 416=>x"3700",
---- 417=>x"3300", 418=>x"2f00", 419=>x"2900", 420=>x"3b00",
---- 421=>x"3a00", 422=>x"3600", 423=>x"2a00", 424=>x"3d00",
---- 425=>x"3100", 426=>x"2f00", 427=>x"3100", 428=>x"4900",
---- 429=>x"4200", 430=>x"3800", 431=>x"3300", 432=>x"4d00",
---- 433=>x"5800", 434=>x"4000", 435=>x"2b00", 436=>x"4900",
---- 437=>x"5d00", 438=>x"4300", 439=>x"2800", 440=>x"3e00",
---- 441=>x"5200", 442=>x"4f00", 443=>x"2a00", 444=>x"4400",
---- 445=>x"4200", 446=>x"4d00", 447=>x"3900", 448=>x"4d00",
---- 449=>x"4200", 450=>x"3d00", 451=>x"3e00", 452=>x"3600",
---- 453=>x"4100", 454=>x"3900", 455=>x"3400", 456=>x"2d00",
---- 457=>x"4000", 458=>x"3800", 459=>x"3100", 460=>x"3500",
---- 461=>x"3f00", 462=>x"2c00", 463=>x"3a00", 464=>x"4600",
---- 465=>x"3e00", 466=>x"2800", 467=>x"2a00", 468=>x"4a00",
---- 469=>x"3700", 470=>x"3100", 471=>x"2d00", 472=>x"4300",
---- 473=>x"4000", 474=>x"3d00", 475=>x"2d00", 476=>x"3b00",
---- 477=>x"3100", 478=>x"4700", 479=>x"3500", 480=>x"3100",
---- 481=>x"2b00", 482=>x"5a00", 483=>x"4900", 484=>x"2600",
---- 485=>x"2800", 486=>x"6100", 487=>x"4a00", 488=>x"1f00",
---- 489=>x"3100", 490=>x"6700", 491=>x"3e00", 492=>x"2a00",
---- 493=>x"3d00", 494=>x"5b00", 495=>x"4300", 496=>x"3a00",
---- 497=>x"4000", 498=>x"4a00", 499=>x"4600", 500=>x"5200",
---- 501=>x"5a00", 502=>x"3900", 503=>x"4b00", 504=>x"5300",
---- 505=>x"7300", 506=>x"3300", 507=>x"4300", 508=>x"2a00",
---- 509=>x"4000", 510=>x"5200", 511=>x"2a00", 512=>x"2b00",
---- 513=>x"2400", 514=>x"3000", 515=>x"3900", 516=>x"2b00",
---- 517=>x"2600", 518=>x"2500", 519=>x"2300", 520=>x"2e00",
---- 521=>x"2500", 522=>x"2800", 523=>x"1800", 524=>x"2900",
---- 525=>x"2500", 526=>x"1e00", 527=>x"3800", 528=>x"2600",
---- 529=>x"2000", 530=>x"1d00", 531=>x"7100", 532=>x"3200",
---- 533=>x"3d00", 534=>x"4700", 535=>x"9600", 536=>x"2500",
---- 537=>x"3400", 538=>x"7000", 539=>x"7300", 540=>x"2400",
---- 541=>x"4c00", 542=>x"7e00", 543=>x"5100", 544=>x"3f00",
---- 545=>x"8900", 546=>x"6c00", 547=>x"6d00", 548=>x"6d00",
---- 549=>x"8b00", 550=>x"5e00", 551=>x"af00", 552=>x"9500",
---- 553=>x"6300", 554=>x"8100", 555=>x"c800", 556=>x"8400",
---- 557=>x"5e00", 558=>x"5200", 559=>x"b100", 560=>x"6500",
---- 561=>x"7c00", 562=>x"b300", 563=>x"a300", 564=>x"6600",
---- 565=>x"a800", 566=>x"ad00", 567=>x"a600", 568=>x"7f00",
---- 569=>x"4800", 570=>x"af00", 571=>x"b300", 572=>x"9c00",
---- 573=>x"b000", 574=>x"b700", 575=>x"bd00", 576=>x"b400",
---- 577=>x"ae00", 578=>x"be00", 579=>x"4000", 580=>x"b400",
---- 581=>x"b800", 582=>x"bd00", 583=>x"c400", 584=>x"b400",
---- 585=>x"c000", 586=>x"c300", 587=>x"d600", 588=>x"bc00",
---- 589=>x"c000", 590=>x"cf00", 591=>x"bd00", 592=>x"bc00",
---- 593=>x"3e00", 594=>x"cf00", 595=>x"5700", 596=>x"bb00",
---- 597=>x"d000", 598=>x"8600", 599=>x"2000", 600=>x"cc00",
---- 601=>x"4d00", 602=>x"3600", 603=>x"2a00", 604=>x"d200",
---- 605=>x"5b00", 606=>x"1d00", 607=>x"2d00", 608=>x"9500",
---- 609=>x"2000", 610=>x"2500", 611=>x"2e00", 612=>x"3f00",
---- 613=>x"1e00", 614=>x"2500", 615=>x"2f00", 616=>x"1b00",
---- 617=>x"2600", 618=>x"2100", 619=>x"3000", 620=>x"2600",
---- 621=>x"2400", 622=>x"2300", 623=>x"3000", 624=>x"2900",
---- 625=>x"2800", 626=>x"2200", 627=>x"3100", 628=>x"2700",
---- 629=>x"2600", 630=>x"2300", 631=>x"3500", 632=>x"2700",
---- 633=>x"2800", 634=>x"2700", 635=>x"3500", 636=>x"2b00",
---- 637=>x"2800", 638=>x"2900", 639=>x"3600", 640=>x"2d00",
---- 641=>x"2d00", 642=>x"2400", 643=>x"3900", 644=>x"3000",
---- 645=>x"2900", 646=>x"2500", 647=>x"3800", 648=>x"3200",
---- 649=>x"3000", 650=>x"2700", 651=>x"3400", 652=>x"2d00",
---- 653=>x"2e00", 654=>x"2a00", 655=>x"3900", 656=>x"2b00",
---- 657=>x"2b00", 658=>x"3000", 659=>x"3a00", 660=>x"3000",
---- 661=>x"2a00", 662=>x"2500", 663=>x"3b00", 664=>x"3500",
---- 665=>x"3000", 666=>x"2a00", 667=>x"3c00", 668=>x"3300",
---- 669=>x"3000", 670=>x"2c00", 671=>x"3d00", 672=>x"3800",
---- 673=>x"3100", 674=>x"2e00", 675=>x"3500", 676=>x"3300",
---- 677=>x"3100", 678=>x"2800", 679=>x"3000", 680=>x"3300",
---- 681=>x"3200", 682=>x"2900", 683=>x"2d00", 684=>x"3b00",
---- 685=>x"3000", 686=>x"2a00", 687=>x"2b00", 688=>x"4400",
---- 689=>x"2d00", 690=>x"2a00", 691=>x"2a00", 692=>x"4200",
---- 693=>x"2e00", 694=>x"2c00", 695=>x"2b00", 696=>x"4900",
---- 697=>x"2f00", 698=>x"2c00", 699=>x"2c00", 700=>x"5100",
---- 701=>x"3300", 702=>x"2600", 703=>x"2900", 704=>x"5100",
---- 705=>x"3a00", 706=>x"2900", 707=>x"2a00", 708=>x"4b00",
---- 709=>x"4000", 710=>x"2c00", 711=>x"2b00", 712=>x"4500",
---- 713=>x"4200", 714=>x"2d00", 715=>x"3000", 716=>x"4500",
---- 717=>x"4700", 718=>x"3100", 719=>x"2c00", 720=>x"4300",
---- 721=>x"4500", 722=>x"3300", 723=>x"2e00", 724=>x"b900",
---- 725=>x"4600", 726=>x"3900", 727=>x"3100", 728=>x"3e00",
---- 729=>x"4700", 730=>x"3d00", 731=>x"3200", 732=>x"3b00",
---- 733=>x"3e00", 734=>x"3a00", 735=>x"3300", 736=>x"3b00",
---- 737=>x"3c00", 738=>x"4200", 739=>x"3900", 740=>x"3900",
---- 741=>x"3d00", 742=>x"4000", 743=>x"3800", 744=>x"3700",
---- 745=>x"3d00", 746=>x"4300", 747=>x"3600", 748=>x"3700",
---- 749=>x"3800", 750=>x"3e00", 751=>x"3800", 752=>x"3700",
---- 753=>x"3900", 754=>x"3700", 755=>x"3b00", 756=>x"3800",
---- 757=>x"3a00", 758=>x"3900", 759=>x"3400", 760=>x"3200",
---- 761=>x"3800", 762=>x"3c00", 763=>x"3400", 764=>x"3200",
---- 765=>x"3400", 766=>x"3d00", 767=>x"3800", 768=>x"2f00",
---- 769=>x"3000", 770=>x"3500", 771=>x"3700", 772=>x"2f00",
---- 773=>x"3000", 774=>x"3400", 775=>x"3400", 776=>x"3400",
---- 777=>x"2e00", 778=>x"3500", 779=>x"3200", 780=>x"3100",
---- 781=>x"2f00", 782=>x"3200", 783=>x"3200", 784=>x"3100",
---- 785=>x"2f00", 786=>x"3100", 787=>x"3200", 788=>x"3100",
---- 789=>x"3300", 790=>x"3400", 791=>x"3900", 792=>x"3000",
---- 793=>x"3400", 794=>x"3400", 795=>x"3200", 796=>x"3200",
---- 797=>x"3000", 798=>x"3100", 799=>x"3000", 800=>x"3500",
---- 801=>x"3400", 802=>x"3200", 803=>x"2d00", 804=>x"3900",
---- 805=>x"3900", 806=>x"3200", 807=>x"ce00", 808=>x"3c00",
---- 809=>x"4600", 810=>x"3300", 811=>x"3400", 812=>x"3900",
---- 813=>x"4000", 814=>x"3a00", 815=>x"3600", 816=>x"4000",
---- 817=>x"3d00", 818=>x"3900", 819=>x"3500", 820=>x"3e00",
---- 821=>x"4300", 822=>x"3500", 823=>x"3000", 824=>x"3e00",
---- 825=>x"4500", 826=>x"3c00", 827=>x"3600", 828=>x"3c00",
---- 829=>x"4600", 830=>x"3a00", 831=>x"3a00", 832=>x"3c00",
---- 833=>x"4800", 834=>x"3700", 835=>x"3100", 836=>x"3b00",
---- 837=>x"4200", 838=>x"3600", 839=>x"3800", 840=>x"4300",
---- 841=>x"4500", 842=>x"3700", 843=>x"3600", 844=>x"3f00",
---- 845=>x"5000", 846=>x"3300", 847=>x"3700", 848=>x"3e00",
---- 849=>x"4500", 850=>x"3100", 851=>x"3200", 852=>x"3c00",
---- 853=>x"4000", 854=>x"3000", 855=>x"2e00", 856=>x"4000",
---- 857=>x"3f00", 858=>x"2d00", 859=>x"2c00", 860=>x"3f00",
---- 861=>x"4100", 862=>x"3400", 863=>x"2a00", 864=>x"3900",
---- 865=>x"3800", 866=>x"3a00", 867=>x"3200", 868=>x"3500",
---- 869=>x"3300", 870=>x"3500", 871=>x"3a00", 872=>x"3500",
---- 873=>x"2f00", 874=>x"3100", 875=>x"3500", 876=>x"3500",
---- 877=>x"3100", 878=>x"3300", 879=>x"3500", 880=>x"3400",
---- 881=>x"3100", 882=>x"3200", 883=>x"3b00", 884=>x"3400",
---- 885=>x"2f00", 886=>x"3000", 887=>x"4100", 888=>x"3000",
---- 889=>x"3000", 890=>x"3200", 891=>x"4500", 892=>x"2f00",
---- 893=>x"3400", 894=>x"3c00", 895=>x"4700", 896=>x"2d00",
---- 897=>x"3400", 898=>x"4300", 899=>x"4e00", 900=>x"2c00",
---- 901=>x"3a00", 902=>x"4b00", 903=>x"5400", 904=>x"3100",
---- 905=>x"3c00", 906=>x"4f00", 907=>x"5600", 908=>x"3600",
---- 909=>x"4800", 910=>x"5200", 911=>x"5700", 912=>x"3900",
---- 913=>x"4a00", 914=>x"5900", 915=>x"6100", 916=>x"4000",
---- 917=>x"4b00", 918=>x"5900", 919=>x"6d00", 920=>x"4600",
---- 921=>x"4f00", 922=>x"5f00", 923=>x"6e00", 924=>x"4800",
---- 925=>x"5600", 926=>x"6900", 927=>x"7000", 928=>x"4e00",
---- 929=>x"5f00", 930=>x"7200", 931=>x"7300", 932=>x"5600",
---- 933=>x"6a00", 934=>x"7300", 935=>x"7800", 936=>x"5f00",
---- 937=>x"7100", 938=>x"7800", 939=>x"7800", 940=>x"6700",
---- 941=>x"7300", 942=>x"7400", 943=>x"7500", 944=>x"6d00",
---- 945=>x"7200", 946=>x"7300", 947=>x"7400", 948=>x"7100",
---- 949=>x"7400", 950=>x"7500", 951=>x"7500", 952=>x"7500",
---- 953=>x"7300", 954=>x"7500", 955=>x"7700", 956=>x"7600",
---- 957=>x"7500", 958=>x"7600", 959=>x"7a00", 960=>x"7400",
---- 961=>x"7300", 962=>x"7800", 963=>x"5f00", 964=>x"7800",
---- 965=>x"7500", 966=>x"5400", 967=>x"2c00", 968=>x"5e00",
---- 969=>x"3e00", 970=>x"2300", 971=>x"2100", 972=>x"2400",
---- 973=>x"2000", 974=>x"3200", 975=>x"4900", 976=>x"3200",
---- 977=>x"4500", 978=>x"5a00", 979=>x"6400", 980=>x"5a00",
---- 981=>x"6200", 982=>x"6700", 983=>x"6b00", 984=>x"6500",
---- 985=>x"7000", 986=>x"7300", 987=>x"7900", 988=>x"7000",
---- 989=>x"7600", 990=>x"7a00", 991=>x"7800", 992=>x"8800",
---- 993=>x"7a00", 994=>x"7a00", 995=>x"7700", 996=>x"7900",
---- 997=>x"7b00", 998=>x"7d00", 999=>x"7f00", 1000=>x"7a00",
---- 1001=>x"7d00", 1002=>x"7d00", 1003=>x"7d00", 1004=>x"7a00",
---- 1005=>x"7d00", 1006=>x"7d00", 1007=>x"7e00", 1008=>x"7900",
---- 1009=>x"7c00", 1010=>x"8100", 1011=>x"8000", 1012=>x"7900",
---- 1013=>x"7a00", 1014=>x"7e00", 1015=>x"8100", 1016=>x"7d00",
---- 1017=>x"7d00", 1018=>x"7d00", 1019=>x"7d00", 1020=>x"7b00",
---- 1021=>x"7d00", 1022=>x"7f00", 1023=>x"8000"),
----
---- 27 => (0=>x"8100", 1=>x"8200", 2=>x"7b00", 3=>x"8200", 4=>x"8300",
---- 5=>x"8200", 6=>x"8400", 7=>x"8100", 8=>x"8100",
---- 9=>x"8200", 10=>x"8600", 11=>x"8300", 12=>x"8200",
---- 13=>x"8100", 14=>x"8200", 15=>x"8200", 16=>x"8300",
---- 17=>x"8000", 18=>x"7f00", 19=>x"7f00", 20=>x"8200",
---- 21=>x"8200", 22=>x"8000", 23=>x"8000", 24=>x"8200",
---- 25=>x"8100", 26=>x"8200", 27=>x"8200", 28=>x"8200",
---- 29=>x"8100", 30=>x"8500", 31=>x"8200", 32=>x"8600",
---- 33=>x"8500", 34=>x"8400", 35=>x"7f00", 36=>x"8900",
---- 37=>x"8200", 38=>x"8200", 39=>x"8100", 40=>x"8300",
---- 41=>x"8200", 42=>x"8700", 43=>x"8300", 44=>x"8000",
---- 45=>x"8200", 46=>x"8100", 47=>x"8000", 48=>x"7f00",
---- 49=>x"7f00", 50=>x"7e00", 51=>x"8100", 52=>x"7f00",
---- 53=>x"8000", 54=>x"7e00", 55=>x"8000", 56=>x"7c00",
---- 57=>x"7e00", 58=>x"8200", 59=>x"8100", 60=>x"7c00",
---- 61=>x"7c00", 62=>x"7e00", 63=>x"8000", 64=>x"7c00",
---- 65=>x"7900", 66=>x"7900", 67=>x"8000", 68=>x"7a00",
---- 69=>x"7900", 70=>x"7c00", 71=>x"7d00", 72=>x"7d00",
---- 73=>x"7b00", 74=>x"7d00", 75=>x"7e00", 76=>x"7d00",
---- 77=>x"7900", 78=>x"7a00", 79=>x"7d00", 80=>x"7d00",
---- 81=>x"7b00", 82=>x"7600", 83=>x"7700", 84=>x"7b00",
---- 85=>x"7a00", 86=>x"7a00", 87=>x"7400", 88=>x"7900",
---- 89=>x"7b00", 90=>x"7e00", 91=>x"8b00", 92=>x"8500",
---- 93=>x"9000", 94=>x"9e00", 95=>x"ac00", 96=>x"a000",
---- 97=>x"a400", 98=>x"5500", 99=>x"aa00", 100=>x"5500",
---- 101=>x"a300", 102=>x"a700", 103=>x"ab00", 104=>x"aa00",
---- 105=>x"a700", 106=>x"a800", 107=>x"ac00", 108=>x"a000",
---- 109=>x"a300", 110=>x"aa00", 111=>x"ab00", 112=>x"a000",
---- 113=>x"9f00", 114=>x"a000", 115=>x"a500", 116=>x"9c00",
---- 117=>x"9f00", 118=>x"a600", 119=>x"a500", 120=>x"9800",
---- 121=>x"a100", 122=>x"aa00", 123=>x"a500", 124=>x"9c00",
---- 125=>x"a800", 126=>x"a000", 127=>x"a000", 128=>x"9e00",
---- 129=>x"a000", 130=>x"9e00", 131=>x"9800", 132=>x"9900",
---- 133=>x"9800", 134=>x"9800", 135=>x"9b00", 136=>x"9200",
---- 137=>x"9a00", 138=>x"9c00", 139=>x"a200", 140=>x"9100",
---- 141=>x"9900", 142=>x"9d00", 143=>x"a200", 144=>x"9300",
---- 145=>x"9000", 146=>x"9900", 147=>x"a000", 148=>x"8c00",
---- 149=>x"9700", 150=>x"9500", 151=>x"9900", 152=>x"9800",
---- 153=>x"6800", 154=>x"9300", 155=>x"9700", 156=>x"9400",
---- 157=>x"9100", 158=>x"9200", 159=>x"9600", 160=>x"8d00",
---- 161=>x"9000", 162=>x"9700", 163=>x"9800", 164=>x"8800",
---- 165=>x"8800", 166=>x"9300", 167=>x"9800", 168=>x"8600",
---- 169=>x"8b00", 170=>x"9300", 171=>x"8c00", 172=>x"8c00",
---- 173=>x"8d00", 174=>x"9000", 175=>x"9f00", 176=>x"8e00",
---- 177=>x"8d00", 178=>x"9500", 179=>x"9400", 180=>x"9300",
---- 181=>x"9800", 182=>x"9100", 183=>x"9100", 184=>x"8f00",
---- 185=>x"8d00", 186=>x"9000", 187=>x"9000", 188=>x"8e00",
---- 189=>x"8900", 190=>x"8d00", 191=>x"9400", 192=>x"9000",
---- 193=>x"8800", 194=>x"9100", 195=>x"6e00", 196=>x"8c00",
---- 197=>x"8e00", 198=>x"9100", 199=>x"9200", 200=>x"8800",
---- 201=>x"8800", 202=>x"8f00", 203=>x"8d00", 204=>x"8900",
---- 205=>x"8d00", 206=>x"8b00", 207=>x"9100", 208=>x"8700",
---- 209=>x"8d00", 210=>x"8d00", 211=>x"8200", 212=>x"8500",
---- 213=>x"8200", 214=>x"7e00", 215=>x"7a00", 216=>x"8200",
---- 217=>x"7600", 218=>x"7e00", 219=>x"9c00", 220=>x"6d00",
---- 221=>x"8100", 222=>x"a400", 223=>x"ad00", 224=>x"9000",
---- 225=>x"b100", 226=>x"b800", 227=>x"b000", 228=>x"a700",
---- 229=>x"b600", 230=>x"ba00", 231=>x"c100", 232=>x"a500",
---- 233=>x"b300", 234=>x"c700", 235=>x"c000", 236=>x"b900",
---- 237=>x"b200", 238=>x"c300", 239=>x"b300", 240=>x"b400",
---- 241=>x"a600", 242=>x"b100", 243=>x"b400", 244=>x"a800",
---- 245=>x"a000", 246=>x"a100", 247=>x"a900", 248=>x"a700",
---- 249=>x"a300", 250=>x"a300", 251=>x"b300", 252=>x"a400",
---- 253=>x"b000", 254=>x"b100", 255=>x"a700", 256=>x"4900",
---- 257=>x"ab00", 258=>x"a200", 259=>x"ad00", 260=>x"a300",
---- 261=>x"a000", 262=>x"b500", 263=>x"b700", 264=>x"a100",
---- 265=>x"5000", 266=>x"af00", 267=>x"b900", 268=>x"b300",
---- 269=>x"ac00", 270=>x"aa00", 271=>x"ab00", 272=>x"af00",
---- 273=>x"ab00", 274=>x"b000", 275=>x"b200", 276=>x"aa00",
---- 277=>x"b200", 278=>x"b300", 279=>x"b300", 280=>x"b400",
---- 281=>x"b300", 282=>x"4c00", 283=>x"a600", 284=>x"ae00",
---- 285=>x"b000", 286=>x"aa00", 287=>x"a900", 288=>x"9500",
---- 289=>x"a400", 290=>x"a900", 291=>x"a700", 292=>x"a000",
---- 293=>x"9c00", 294=>x"a100", 295=>x"ae00", 296=>x"9f00",
---- 297=>x"a500", 298=>x"aa00", 299=>x"aa00", 300=>x"ac00",
---- 301=>x"ad00", 302=>x"af00", 303=>x"ad00", 304=>x"a500",
---- 305=>x"b700", 306=>x"ae00", 307=>x"a900", 308=>x"9f00",
---- 309=>x"9e00", 310=>x"b100", 311=>x"a200", 312=>x"a300",
---- 313=>x"9c00", 314=>x"9600", 315=>x"9400", 316=>x"9800",
---- 317=>x"9f00", 318=>x"8900", 319=>x"9800", 320=>x"8b00",
---- 321=>x"8e00", 322=>x"a700", 323=>x"9d00", 324=>x"8b00",
---- 325=>x"9300", 326=>x"a400", 327=>x"a800", 328=>x"5f00",
---- 329=>x"a300", 330=>x"9900", 331=>x"9c00", 332=>x"9e00",
---- 333=>x"9f00", 334=>x"a000", 335=>x"6500", 336=>x"9a00",
---- 337=>x"9b00", 338=>x"9e00", 339=>x"9d00", 340=>x"a200",
---- 341=>x"9c00", 342=>x"9700", 343=>x"8800", 344=>x"9300",
---- 345=>x"7400", 346=>x"6900", 347=>x"6b00", 348=>x"6100",
---- 349=>x"6200", 350=>x"8800", 351=>x"8c00", 352=>x"7300",
---- 353=>x"8b00", 354=>x"9100", 355=>x"8900", 356=>x"9800",
---- 357=>x"8e00", 358=>x"8700", 359=>x"6b00", 360=>x"9400",
---- 361=>x"8300", 362=>x"6600", 363=>x"5f00", 364=>x"8500",
---- 365=>x"7200", 366=>x"6800", 367=>x"8000", 368=>x"7400",
---- 369=>x"6700", 370=>x"8000", 371=>x"7f00", 372=>x"6700",
---- 373=>x"7c00", 374=>x"8400", 375=>x"7400", 376=>x"6700",
---- 377=>x"7000", 378=>x"5700", 379=>x"4c00", 380=>x"5000",
---- 381=>x"4300", 382=>x"3e00", 383=>x"5200", 384=>x"3100",
---- 385=>x"4f00", 386=>x"6b00", 387=>x"5800", 388=>x"5d00",
---- 389=>x"6300", 390=>x"4300", 391=>x"2f00", 392=>x"5200",
---- 393=>x"3500", 394=>x"2f00", 395=>x"2b00", 396=>x"3800",
---- 397=>x"3d00", 398=>x"3500", 399=>x"3000", 400=>x"3e00",
---- 401=>x"3500", 402=>x"3300", 403=>x"5a00", 404=>x"3000",
---- 405=>x"2500", 406=>x"5300", 407=>x"6d00", 408=>x"2b00",
---- 409=>x"3e00", 410=>x"7400", 411=>x"6500", 412=>x"2e00",
---- 413=>x"4a00", 414=>x"7a00", 415=>x"5500", 416=>x"2b00",
---- 417=>x"5500", 418=>x"7800", 419=>x"4100", 420=>x"3600",
---- 421=>x"5100", 422=>x"5e00", 423=>x"4600", 424=>x"4100",
---- 425=>x"4400", 426=>x"b400", 427=>x"5800", 428=>x"4b00",
---- 429=>x"3b00", 430=>x"3c00", 431=>x"6e00", 432=>x"4a00",
---- 433=>x"3800", 434=>x"3300", 435=>x"6600", 436=>x"4a00",
---- 437=>x"4200", 438=>x"2300", 439=>x"4c00", 440=>x"4300",
---- 441=>x"4e00", 442=>x"2100", 443=>x"3200", 444=>x"4600",
---- 445=>x"5200", 446=>x"2800", 447=>x"3800", 448=>x"5100",
---- 449=>x"4600", 450=>x"3300", 451=>x"3f00", 452=>x"5800",
---- 453=>x"5800", 454=>x"5100", 455=>x"4600", 456=>x"4200",
---- 457=>x"6a00", 458=>x"7900", 459=>x"5800", 460=>x"4f00",
---- 461=>x"5900", 462=>x"5900", 463=>x"6200", 464=>x"6000",
---- 465=>x"5100", 466=>x"4900", 467=>x"4b00", 468=>x"4c00",
---- 469=>x"3700", 470=>x"4a00", 471=>x"3f00", 472=>x"2a00",
---- 473=>x"3600", 474=>x"5000", 475=>x"4600", 476=>x"3200",
---- 477=>x"2c00", 478=>x"6500", 479=>x"5e00", 480=>x"3100",
---- 481=>x"3a00", 482=>x"6300", 483=>x"2f00", 484=>x"1f00",
---- 485=>x"5700", 486=>x"3a00", 487=>x"2d00", 488=>x"2d00",
---- 489=>x"5b00", 490=>x"3c00", 491=>x"c700", 492=>x"3a00",
---- 493=>x"4900", 494=>x"2600", 495=>x"1d00", 496=>x"3600",
---- 497=>x"3900", 498=>x"1f00", 499=>x"2900", 500=>x"3b00",
---- 501=>x"2b00", 502=>x"1f00", 503=>x"5600", 504=>x"3500",
---- 505=>x"1800", 506=>x"3200", 507=>x"8f00", 508=>x"1e00",
---- 509=>x"2200", 510=>x"7200", 511=>x"9100", 512=>x"1800",
---- 513=>x"4900", 514=>x"9d00", 515=>x"6e00", 516=>x"2b00",
---- 517=>x"8900", 518=>x"8c00", 519=>x"6a00", 520=>x"5e00",
---- 521=>x"9f00", 522=>x"6a00", 523=>x"9d00", 524=>x"9600",
---- 525=>x"7800", 526=>x"7900", 527=>x"c400", 528=>x"9500",
---- 529=>x"6000", 530=>x"ac00", 531=>x"b900", 532=>x"6b00",
---- 533=>x"8c00", 534=>x"c800", 535=>x"a900", 536=>x"6700",
---- 537=>x"b400", 538=>x"ac00", 539=>x"9700", 540=>x"8e00",
---- 541=>x"a500", 542=>x"9700", 543=>x"a500", 544=>x"bb00",
---- 545=>x"9c00", 546=>x"a900", 547=>x"b600", 548=>x"be00",
---- 549=>x"9d00", 550=>x"af00", 551=>x"b800", 552=>x"a900",
---- 553=>x"ab00", 554=>x"b700", 555=>x"be00", 556=>x"a400",
---- 557=>x"b300", 558=>x"ba00", 559=>x"c500", 560=>x"af00",
---- 561=>x"b200", 562=>x"be00", 563=>x"c800", 564=>x"b500",
---- 565=>x"b900", 566=>x"c600", 567=>x"d200", 568=>x"bb00",
---- 569=>x"c400", 570=>x"d200", 571=>x"b000", 572=>x"c200",
---- 573=>x"d200", 574=>x"be00", 575=>x"5000", 576=>x"c600",
---- 577=>x"ca00", 578=>x"6000", 579=>x"3900", 580=>x"d100",
---- 581=>x"7900", 582=>x"2d00", 583=>x"4800", 584=>x"9800",
---- 585=>x"2700", 586=>x"3400", 587=>x"4c00", 588=>x"3800",
---- 589=>x"2300", 590=>x"3900", 591=>x"5200", 592=>x"2000",
---- 593=>x"3400", 594=>x"3b00", 595=>x"5400", 596=>x"2c00",
---- 597=>x"3100", 598=>x"4200", 599=>x"5800", 600=>x"3600",
---- 601=>x"3200", 602=>x"3f00", 603=>x"5800", 604=>x"3900",
---- 605=>x"3200", 606=>x"3f00", 607=>x"5400", 608=>x"4200",
---- 609=>x"3400", 610=>x"4300", 611=>x"5500", 612=>x"4a00",
---- 613=>x"3400", 614=>x"3d00", 615=>x"5400", 616=>x"4f00",
---- 617=>x"3800", 618=>x"3d00", 619=>x"5100", 620=>x"5600",
---- 621=>x"3b00", 622=>x"4300", 623=>x"4e00", 624=>x"5f00",
---- 625=>x"4500", 626=>x"4400", 627=>x"5100", 628=>x"6700",
---- 629=>x"4400", 630=>x"4200", 631=>x"5200", 632=>x"6900",
---- 633=>x"4800", 634=>x"4500", 635=>x"5000", 636=>x"6b00",
---- 637=>x"5600", 638=>x"4200", 639=>x"4e00", 640=>x"6900",
---- 641=>x"5500", 642=>x"4000", 643=>x"5000", 644=>x"6a00",
---- 645=>x"5700", 646=>x"4b00", 647=>x"5700", 648=>x"6c00",
---- 649=>x"6000", 650=>x"4b00", 651=>x"5d00", 652=>x"7100",
---- 653=>x"6300", 654=>x"4a00", 655=>x"5e00", 656=>x"7400",
---- 657=>x"6a00", 658=>x"5000", 659=>x"5900", 660=>x"7900",
---- 661=>x"6700", 662=>x"5200", 663=>x"5a00", 664=>x"7500",
---- 665=>x"6900", 666=>x"5400", 667=>x"5b00", 668=>x"6e00",
---- 669=>x"6b00", 670=>x"5d00", 671=>x"5f00", 672=>x"6a00",
---- 673=>x"6f00", 674=>x"5f00", 675=>x"5e00", 676=>x"6700",
---- 677=>x"6900", 678=>x"6500", 679=>x"5b00", 680=>x"5e00",
---- 681=>x"6500", 682=>x"6a00", 683=>x"5700", 684=>x"5e00",
---- 685=>x"6400", 686=>x"6900", 687=>x"5600", 688=>x"5700",
---- 689=>x"6000", 690=>x"6600", 691=>x"5900", 692=>x"5800",
---- 693=>x"5b00", 694=>x"6200", 695=>x"5700", 696=>x"5c00",
---- 697=>x"5c00", 698=>x"5c00", 699=>x"5300", 700=>x"5600",
---- 701=>x"5200", 702=>x"5700", 703=>x"5a00", 704=>x"5200",
---- 705=>x"5200", 706=>x"5500", 707=>x"5800", 708=>x"5200",
---- 709=>x"4e00", 710=>x"4f00", 711=>x"5300", 712=>x"5000",
---- 713=>x"4a00", 714=>x"4b00", 715=>x"5400", 716=>x"bb00",
---- 717=>x"4500", 718=>x"4b00", 719=>x"5400", 720=>x"4700",
---- 721=>x"4d00", 722=>x"4c00", 723=>x"5100", 724=>x"4400",
---- 725=>x"4f00", 726=>x"4900", 727=>x"4e00", 728=>x"3b00",
---- 729=>x"4c00", 730=>x"4600", 731=>x"5500", 732=>x"3600",
---- 733=>x"4900", 734=>x"4100", 735=>x"5200", 736=>x"3100",
---- 737=>x"3f00", 738=>x"3b00", 739=>x"4b00", 740=>x"2c00",
---- 741=>x"3a00", 742=>x"3d00", 743=>x"3e00", 744=>x"2f00",
---- 745=>x"3500", 746=>x"4000", 747=>x"3a00", 748=>x"3200",
---- 749=>x"3200", 750=>x"3e00", 751=>x"3b00", 752=>x"3600",
---- 753=>x"3500", 754=>x"3b00", 755=>x"3900", 756=>x"3800",
---- 757=>x"3900", 758=>x"3b00", 759=>x"3a00", 760=>x"3b00",
---- 761=>x"3300", 762=>x"3900", 763=>x"3d00", 764=>x"3c00",
---- 765=>x"3d00", 766=>x"3400", 767=>x"3a00", 768=>x"3e00",
---- 769=>x"3d00", 770=>x"3700", 771=>x"3b00", 772=>x"3a00",
---- 773=>x"3f00", 774=>x"3d00", 775=>x"3f00", 776=>x"3800",
---- 777=>x"3d00", 778=>x"3e00", 779=>x"3800", 780=>x"3400",
---- 781=>x"3b00", 782=>x"3b00", 783=>x"3600", 784=>x"3600",
---- 785=>x"3900", 786=>x"3d00", 787=>x"3900", 788=>x"3300",
---- 789=>x"3400", 790=>x"3d00", 791=>x"3f00", 792=>x"3600",
---- 793=>x"2f00", 794=>x"3a00", 795=>x"3c00", 796=>x"3200",
---- 797=>x"3300", 798=>x"3b00", 799=>x"4000", 800=>x"3100",
---- 801=>x"3a00", 802=>x"3900", 803=>x"3c00", 804=>x"3300",
---- 805=>x"3600", 806=>x"3600", 807=>x"3900", 808=>x"3100",
---- 809=>x"3500", 810=>x"3600", 811=>x"3800", 812=>x"3300",
---- 813=>x"3200", 814=>x"3e00", 815=>x"3e00", 816=>x"3400",
---- 817=>x"3000", 818=>x"3b00", 819=>x"3e00", 820=>x"3600",
---- 821=>x"3400", 822=>x"3e00", 823=>x"4500", 824=>x"3800",
---- 825=>x"3700", 826=>x"4600", 827=>x"4e00", 828=>x"3800",
---- 829=>x"3400", 830=>x"3f00", 831=>x"4a00", 832=>x"2e00",
---- 833=>x"2c00", 834=>x"3700", 835=>x"4700", 836=>x"3100",
---- 837=>x"2a00", 838=>x"3800", 839=>x"4800", 840=>x"3a00",
---- 841=>x"3000", 842=>x"3300", 843=>x"3e00", 844=>x"3900",
---- 845=>x"2d00", 846=>x"3700", 847=>x"3a00", 848=>x"3100",
---- 849=>x"2d00", 850=>x"3400", 851=>x"3600", 852=>x"3800",
---- 853=>x"3900", 854=>x"3500", 855=>x"3a00", 856=>x"3300",
---- 857=>x"3100", 858=>x"3900", 859=>x"4300", 860=>x"2d00",
---- 861=>x"3700", 862=>x"3600", 863=>x"4d00", 864=>x"3100",
---- 865=>x"3b00", 866=>x"3b00", 867=>x"4e00", 868=>x"3500",
---- 869=>x"3900", 870=>x"ba00", 871=>x"5c00", 872=>x"3b00",
---- 873=>x"3e00", 874=>x"5200", 875=>x"6e00", 876=>x"4300",
---- 877=>x"4600", 878=>x"5a00", 879=>x"7600", 880=>x"4600",
---- 881=>x"4c00", 882=>x"6200", 883=>x"7800", 884=>x"4800",
---- 885=>x"5000", 886=>x"6600", 887=>x"7900", 888=>x"4e00",
---- 889=>x"5800", 890=>x"6d00", 891=>x"7d00", 892=>x"5300",
---- 893=>x"6000", 894=>x"7400", 895=>x"7c00", 896=>x"5900",
---- 897=>x"6400", 898=>x"7600", 899=>x"7b00", 900=>x"5e00",
---- 901=>x"6b00", 902=>x"7800", 903=>x"7e00", 904=>x"6600",
---- 905=>x"6b00", 906=>x"7700", 907=>x"7a00", 908=>x"6a00",
---- 909=>x"7000", 910=>x"7600", 911=>x"7c00", 912=>x"6f00",
---- 913=>x"7700", 914=>x"7800", 915=>x"7c00", 916=>x"7100",
---- 917=>x"7400", 918=>x"7900", 919=>x"7f00", 920=>x"7200",
---- 921=>x"7500", 922=>x"7800", 923=>x"7e00", 924=>x"7500",
---- 925=>x"7400", 926=>x"7a00", 927=>x"7e00", 928=>x"7300",
---- 929=>x"7400", 930=>x"7800", 931=>x"7c00", 932=>x"7600",
---- 933=>x"7400", 934=>x"7500", 935=>x"7700", 936=>x"7700",
---- 937=>x"7700", 938=>x"7700", 939=>x"7700", 940=>x"7600",
---- 941=>x"7800", 942=>x"7800", 943=>x"6a00", 944=>x"8900",
---- 945=>x"7700", 946=>x"7200", 947=>x"4a00", 948=>x"7900",
---- 949=>x"7900", 950=>x"5200", 951=>x"2c00", 952=>x"7800",
---- 953=>x"6000", 954=>x"3400", 955=>x"2500", 956=>x"6200",
---- 957=>x"2f00", 958=>x"2a00", 959=>x"3400", 960=>x"2d00",
---- 961=>x"2000", 962=>x"2d00", 963=>x"b200", 964=>x"2300",
---- 965=>x"3000", 966=>x"4a00", 967=>x"6200", 968=>x"3700",
---- 969=>x"5500", 970=>x"6100", 971=>x"6c00", 972=>x"5f00",
---- 973=>x"6a00", 974=>x"6f00", 975=>x"7500", 976=>x"6a00",
---- 977=>x"7100", 978=>x"8700", 979=>x"7800", 980=>x"7200",
---- 981=>x"7600", 982=>x"8100", 983=>x"7b00", 984=>x"7e00",
---- 985=>x"7d00", 986=>x"7e00", 987=>x"7d00", 988=>x"7c00",
---- 989=>x"7900", 990=>x"7d00", 991=>x"7f00", 992=>x"7d00",
---- 993=>x"7c00", 994=>x"7d00", 995=>x"8000", 996=>x"7e00",
---- 997=>x"7f00", 998=>x"7f00", 999=>x"8100", 1000=>x"7f00",
---- 1001=>x"8000", 1002=>x"8200", 1003=>x"7f00", 1004=>x"8300",
---- 1005=>x"8000", 1006=>x"7f00", 1007=>x"7c00", 1008=>x"7c00",
---- 1009=>x"7e00", 1010=>x"7d00", 1011=>x"7c00", 1012=>x"7f00",
---- 1013=>x"7d00", 1014=>x"7f00", 1015=>x"8000", 1016=>x"7e00",
---- 1017=>x"7e00", 1018=>x"8100", 1019=>x"8100", 1020=>x"7e00",
---- 1021=>x"7f00", 1022=>x"8000", 1023=>x"8000"),
----
---- 28 => (0=>x"8200", 1=>x"8500", 2=>x"8700", 3=>x"8400", 4=>x"8200",
---- 5=>x"8500", 6=>x"8600", 7=>x"8400", 8=>x"8200",
---- 9=>x"8100", 10=>x"8600", 11=>x"8400", 12=>x"8100",
---- 13=>x"8300", 14=>x"8700", 15=>x"8200", 16=>x"8200",
---- 17=>x"8700", 18=>x"8500", 19=>x"8400", 20=>x"8200",
---- 21=>x"8100", 22=>x"8100", 23=>x"8200", 24=>x"8200",
---- 25=>x"8100", 26=>x"8300", 27=>x"8400", 28=>x"8100",
---- 29=>x"8400", 30=>x"8200", 31=>x"8200", 32=>x"7e00",
---- 33=>x"8400", 34=>x"8400", 35=>x"8400", 36=>x"7f00",
---- 37=>x"8400", 38=>x"8500", 39=>x"8300", 40=>x"8300",
---- 41=>x"8300", 42=>x"8200", 43=>x"8300", 44=>x"8400",
---- 45=>x"8200", 46=>x"8000", 47=>x"8100", 48=>x"7f00",
---- 49=>x"8000", 50=>x"7f00", 51=>x"8000", 52=>x"8000",
---- 53=>x"7d00", 54=>x"7e00", 55=>x"7e00", 56=>x"7d00",
---- 57=>x"7d00", 58=>x"7c00", 59=>x"7c00", 60=>x"7f00",
---- 61=>x"7e00", 62=>x"7d00", 63=>x"7f00", 64=>x"7d00",
---- 65=>x"7b00", 66=>x"7d00", 67=>x"7e00", 68=>x"7d00",
---- 69=>x"8100", 70=>x"7d00", 71=>x"7a00", 72=>x"7c00",
---- 73=>x"7f00", 74=>x"7b00", 75=>x"7900", 76=>x"7d00",
---- 77=>x"7900", 78=>x"7700", 79=>x"7800", 80=>x"7900",
---- 81=>x"7800", 82=>x"7800", 83=>x"7900", 84=>x"7400",
---- 85=>x"7700", 86=>x"7500", 87=>x"7600", 88=>x"8a00",
---- 89=>x"8800", 90=>x"8900", 91=>x"8000", 92=>x"a400",
---- 93=>x"b100", 94=>x"ac00", 95=>x"a800", 96=>x"b000",
---- 97=>x"ac00", 98=>x"ab00", 99=>x"b100", 100=>x"b200",
---- 101=>x"b600", 102=>x"b200", 103=>x"b100", 104=>x"b400",
---- 105=>x"b700", 106=>x"b500", 107=>x"b200", 108=>x"b100",
---- 109=>x"b200", 110=>x"b500", 111=>x"b400", 112=>x"a300",
---- 113=>x"ae00", 114=>x"b500", 115=>x"b300", 116=>x"a600",
---- 117=>x"a300", 118=>x"b000", 119=>x"af00", 120=>x"5900",
---- 121=>x"ac00", 122=>x"a700", 123=>x"a300", 124=>x"a600",
---- 125=>x"a700", 126=>x"a700", 127=>x"ab00", 128=>x"a200",
---- 129=>x"a000", 130=>x"ae00", 131=>x"ad00", 132=>x"ab00",
---- 133=>x"ae00", 134=>x"ab00", 135=>x"a900", 136=>x"a500",
---- 137=>x"ae00", 138=>x"af00", 139=>x"b000", 140=>x"a300",
---- 141=>x"5200", 142=>x"af00", 143=>x"b200", 144=>x"a400",
---- 145=>x"a800", 146=>x"a700", 147=>x"ac00", 148=>x"9f00",
---- 149=>x"a100", 150=>x"a200", 151=>x"a500", 152=>x"9b00",
---- 153=>x"9e00", 154=>x"9f00", 155=>x"ac00", 156=>x"9b00",
---- 157=>x"a100", 158=>x"a700", 159=>x"aa00", 160=>x"a200",
---- 161=>x"9800", 162=>x"a400", 163=>x"b000", 164=>x"9700",
---- 165=>x"a100", 166=>x"a600", 167=>x"a600", 168=>x"9f00",
---- 169=>x"6300", 170=>x"a300", 171=>x"ab00", 172=>x"9b00",
---- 173=>x"9d00", 174=>x"a800", 175=>x"a500", 176=>x"9d00",
---- 177=>x"9800", 178=>x"a300", 179=>x"ab00", 180=>x"9600",
---- 181=>x"9c00", 182=>x"a300", 183=>x"9c00", 184=>x"9400",
---- 185=>x"9800", 186=>x"a200", 187=>x"ac00", 188=>x"9100",
---- 189=>x"9b00", 190=>x"a700", 191=>x"a300", 192=>x"9c00",
---- 193=>x"9b00", 194=>x"a000", 195=>x"5300", 196=>x"9000",
---- 197=>x"9900", 198=>x"ac00", 199=>x"a900", 200=>x"9400",
---- 201=>x"a100", 202=>x"a200", 203=>x"8e00", 204=>x"8700",
---- 205=>x"9000", 206=>x"8600", 207=>x"8c00", 208=>x"8000",
---- 209=>x"8200", 210=>x"6600", 211=>x"b100", 212=>x"8d00",
---- 213=>x"b300", 214=>x"b900", 215=>x"b000", 216=>x"ae00",
---- 217=>x"c300", 218=>x"ba00", 219=>x"b500", 220=>x"b500",
---- 221=>x"b900", 222=>x"c700", 223=>x"bf00", 224=>x"ba00",
---- 225=>x"4000", 226=>x"c200", 227=>x"3d00", 228=>x"b800",
---- 229=>x"b900", 230=>x"b700", 231=>x"b700", 232=>x"b900",
---- 233=>x"ad00", 234=>x"ad00", 235=>x"ae00", 236=>x"b000",
---- 237=>x"b200", 238=>x"ad00", 239=>x"b100", 240=>x"ab00",
---- 241=>x"b100", 242=>x"b900", 243=>x"ae00", 244=>x"bb00",
---- 245=>x"ba00", 246=>x"a900", 247=>x"a800", 248=>x"ac00",
---- 249=>x"a600", 250=>x"ac00", 251=>x"bd00", 252=>x"a900",
---- 253=>x"b300", 254=>x"b200", 255=>x"4b00", 256=>x"ba00",
---- 257=>x"b900", 258=>x"b200", 259=>x"ae00", 260=>x"b400",
---- 261=>x"b700", 262=>x"b300", 263=>x"aa00", 264=>x"b500",
---- 265=>x"ac00", 266=>x"b600", 267=>x"ba00", 268=>x"b500",
---- 269=>x"b900", 270=>x"b400", 271=>x"bf00", 272=>x"af00",
---- 273=>x"b700", 274=>x"b000", 275=>x"ad00", 276=>x"ae00",
---- 277=>x"a600", 278=>x"aa00", 279=>x"ab00", 280=>x"a700",
---- 281=>x"a800", 282=>x"a400", 283=>x"a300", 284=>x"5900",
---- 285=>x"a500", 286=>x"af00", 287=>x"b100", 288=>x"ac00",
---- 289=>x"ab00", 290=>x"a700", 291=>x"b800", 292=>x"b600",
---- 293=>x"b700", 294=>x"ac00", 295=>x"a300", 296=>x"b100",
---- 297=>x"b700", 298=>x"b500", 299=>x"a000", 300=>x"a200",
---- 301=>x"a300", 302=>x"a600", 303=>x"9900", 304=>x"a900",
---- 305=>x"8e00", 306=>x"9300", 307=>x"ad00", 308=>x"9700",
---- 309=>x"9600", 310=>x"a500", 311=>x"b300", 312=>x"9d00",
---- 313=>x"b000", 314=>x"af00", 315=>x"aa00", 316=>x"aa00",
---- 317=>x"ac00", 318=>x"b100", 319=>x"ab00", 320=>x"6000",
---- 321=>x"a800", 322=>x"a500", 323=>x"a300", 324=>x"9e00",
---- 325=>x"9700", 326=>x"9900", 327=>x"9e00", 328=>x"a300",
---- 329=>x"9d00", 330=>x"9600", 331=>x"9f00", 332=>x"9200",
---- 333=>x"9e00", 334=>x"a900", 335=>x"9600", 336=>x"9800",
---- 337=>x"9600", 338=>x"a600", 339=>x"a300", 340=>x"8800",
---- 341=>x"8b00", 342=>x"8700", 343=>x"9200", 344=>x"6c00",
---- 345=>x"6600", 346=>x"6200", 347=>x"6200", 348=>x"8900",
---- 349=>x"7700", 350=>x"7400", 351=>x"6a00", 352=>x"7e00",
---- 353=>x"7a00", 354=>x"7200", 355=>x"6c00", 356=>x"6300",
---- 357=>x"6900", 358=>x"5f00", 359=>x"4c00", 360=>x"6c00",
---- 361=>x"9700", 362=>x"5700", 363=>x"5e00", 364=>x"7b00",
---- 365=>x"6500", 366=>x"7200", 367=>x"8b00", 368=>x"6f00",
---- 369=>x"6c00", 370=>x"7b00", 371=>x"7000", 372=>x"7400",
---- 373=>x"5700", 374=>x"4500", 375=>x"3a00", 376=>x"5000",
---- 377=>x"4700", 378=>x"4700", 379=>x"3c00", 380=>x"5d00",
---- 381=>x"4f00", 382=>x"4600", 383=>x"3500", 384=>x"4200",
---- 385=>x"3700", 386=>x"3600", 387=>x"2f00", 388=>x"2b00",
---- 389=>x"3300", 390=>x"3900", 391=>x"2e00", 392=>x"3400",
---- 393=>x"3f00", 394=>x"2b00", 395=>x"2a00", 396=>x"4a00",
---- 397=>x"3700", 398=>x"2400", 399=>x"2800", 400=>x"4900",
---- 401=>x"2400", 402=>x"2500", 403=>x"2a00", 404=>x"2c00",
---- 405=>x"2600", 406=>x"2700", 407=>x"3400", 408=>x"2000",
---- 409=>x"2800", 410=>x"2900", 411=>x"3900", 412=>x"2300",
---- 413=>x"2b00", 414=>x"2e00", 415=>x"c500", 416=>x"2100",
---- 417=>x"2d00", 418=>x"4f00", 419=>x"4000", 420=>x"2d00",
---- 421=>x"3f00", 422=>x"5300", 423=>x"3000", 424=>x"4d00",
---- 425=>x"4600", 426=>x"2f00", 427=>x"2e00", 428=>x"6800",
---- 429=>x"4600", 430=>x"2a00", 431=>x"2e00", 432=>x"7e00",
---- 433=>x"5700", 434=>x"2700", 435=>x"2c00", 436=>x"7d00",
---- 437=>x"7c00", 438=>x"4300", 439=>x"2b00", 440=>x"5100",
---- 441=>x"8a00", 442=>x"6f00", 443=>x"5700", 444=>x"3600",
---- 445=>x"8600", 446=>x"5e00", 447=>x"3900", 448=>x"3300",
---- 449=>x"8200", 450=>x"5f00", 451=>x"2000", 452=>x"2400",
---- 453=>x"5f00", 454=>x"7600", 455=>x"2700", 456=>x"d300",
---- 457=>x"3f00", 458=>x"7c00", 459=>x"3300", 460=>x"5300",
---- 461=>x"4d00", 462=>x"9400", 463=>x"5e00", 464=>x"3e00",
---- 465=>x"3b00", 466=>x"8a00", 467=>x"5d00", 468=>x"2100",
---- 469=>x"1b00", 470=>x"5500", 471=>x"7a00", 472=>x"1d00",
---- 473=>x"1f00", 474=>x"2e00", 475=>x"6e00", 476=>x"1b00",
---- 477=>x"1f00", 478=>x"1e00", 479=>x"4500", 480=>x"2800",
---- 481=>x"2000", 482=>x"2d00", 483=>x"7200", 484=>x"3400",
---- 485=>x"2200", 486=>x"6300", 487=>x"9700", 488=>x"2100",
---- 489=>x"4c00", 490=>x"9b00", 491=>x"7600", 492=>x"3400",
---- 493=>x"8e00", 494=>x"8300", 495=>x"a500", 496=>x"7300",
---- 497=>x"9600", 498=>x"5b00", 499=>x"8000", 500=>x"a100",
---- 501=>x"7300", 502=>x"7300", 503=>x"b900", 504=>x"9600",
---- 505=>x"7100", 506=>x"a900", 507=>x"b700", 508=>x"6900",
---- 509=>x"9d00", 510=>x"bd00", 511=>x"a500", 512=>x"8000",
---- 513=>x"c000", 514=>x"aa00", 515=>x"a900", 516=>x"b500",
---- 517=>x"b200", 518=>x"aa00", 519=>x"b000", 520=>x"bf00",
---- 521=>x"a500", 522=>x"b000", 523=>x"b400", 524=>x"ac00",
---- 525=>x"a800", 526=>x"b000", 527=>x"b600", 528=>x"a700",
---- 529=>x"b200", 530=>x"b200", 531=>x"b600", 532=>x"b200",
---- 533=>x"b800", 534=>x"b600", 535=>x"c100", 536=>x"a000",
---- 537=>x"b100", 538=>x"bd00", 539=>x"c900", 540=>x"b100",
---- 541=>x"be00", 542=>x"c600", 543=>x"c700", 544=>x"bd00",
---- 545=>x"c600", 546=>x"c800", 547=>x"c400", 548=>x"c200",
---- 549=>x"c900", 550=>x"c500", 551=>x"c500", 552=>x"c900",
---- 553=>x"c700", 554=>x"c800", 555=>x"8f00", 556=>x"c800",
---- 557=>x"cb00", 558=>x"9100", 559=>x"5600", 560=>x"ce00",
---- 561=>x"9600", 562=>x"4c00", 563=>x"5f00", 564=>x"9e00",
---- 565=>x"4b00", 566=>x"5a00", 567=>x"6c00", 568=>x"4900",
---- 569=>x"5400", 570=>x"9500", 571=>x"6f00", 572=>x"4700",
---- 573=>x"6200", 574=>x"7000", 575=>x"7400", 576=>x"5700",
---- 577=>x"6600", 578=>x"7000", 579=>x"7800", 580=>x"5800",
---- 581=>x"6d00", 582=>x"7200", 583=>x"7700", 584=>x"5b00",
---- 585=>x"6f00", 586=>x"7600", 587=>x"7800", 588=>x"6400",
---- 589=>x"7100", 590=>x"7900", 591=>x"8400", 592=>x"6600",
---- 593=>x"7500", 594=>x"7900", 595=>x"7b00", 596=>x"6b00",
---- 597=>x"7500", 598=>x"7700", 599=>x"7d00", 600=>x"6a00",
---- 601=>x"7500", 602=>x"7800", 603=>x"7800", 604=>x"6700",
---- 605=>x"7300", 606=>x"7b00", 607=>x"7a00", 608=>x"6500",
---- 609=>x"6f00", 610=>x"7600", 611=>x"7d00", 612=>x"6200",
---- 613=>x"6c00", 614=>x"7300", 615=>x"7900", 616=>x"6400",
---- 617=>x"6b00", 618=>x"7400", 619=>x"7b00", 620=>x"6200",
---- 621=>x"6c00", 622=>x"7200", 623=>x"7d00", 624=>x"6000",
---- 625=>x"6900", 626=>x"7600", 627=>x"7900", 628=>x"5c00",
---- 629=>x"6900", 630=>x"7200", 631=>x"7600", 632=>x"5900",
---- 633=>x"6b00", 634=>x"7200", 635=>x"7700", 636=>x"5d00",
---- 637=>x"6d00", 638=>x"7400", 639=>x"7a00", 640=>x"6000",
---- 641=>x"6e00", 642=>x"7400", 643=>x"7900", 644=>x"6000",
---- 645=>x"6b00", 646=>x"7400", 647=>x"7900", 648=>x"6300",
---- 649=>x"6900", 650=>x"7200", 651=>x"7700", 652=>x"6800",
---- 653=>x"7000", 654=>x"7200", 655=>x"7700", 656=>x"6b00",
---- 657=>x"7000", 658=>x"7400", 659=>x"7800", 660=>x"6c00",
---- 661=>x"7300", 662=>x"7500", 663=>x"7800", 664=>x"6a00",
---- 665=>x"7000", 666=>x"7700", 667=>x"7900", 668=>x"6b00",
---- 669=>x"7300", 670=>x"7900", 671=>x"7d00", 672=>x"6f00",
---- 673=>x"7100", 674=>x"7800", 675=>x"7d00", 676=>x"6900",
---- 677=>x"7100", 678=>x"7500", 679=>x"7800", 680=>x"6700",
---- 681=>x"7000", 682=>x"7400", 683=>x"7a00", 684=>x"5e00",
---- 685=>x"6c00", 686=>x"7300", 687=>x"7b00", 688=>x"5900",
---- 689=>x"6900", 690=>x"7200", 691=>x"7600", 692=>x"5300",
---- 693=>x"6400", 694=>x"7000", 695=>x"7700", 696=>x"4f00",
---- 697=>x"6300", 698=>x"6c00", 699=>x"7100", 700=>x"4800",
---- 701=>x"5c00", 702=>x"6b00", 703=>x"7500", 704=>x"4d00",
---- 705=>x"5a00", 706=>x"6400", 707=>x"7100", 708=>x"4d00",
---- 709=>x"5800", 710=>x"6400", 711=>x"6e00", 712=>x"4b00",
---- 713=>x"4c00", 714=>x"5e00", 715=>x"6b00", 716=>x"4200",
---- 717=>x"4b00", 718=>x"5a00", 719=>x"6700", 720=>x"3f00",
---- 721=>x"4900", 722=>x"5700", 723=>x"6300", 724=>x"4000",
---- 725=>x"4300", 726=>x"4f00", 727=>x"5c00", 728=>x"4100",
---- 729=>x"4200", 730=>x"4a00", 731=>x"5100", 732=>x"4200",
---- 733=>x"3a00", 734=>x"4900", 735=>x"5000", 736=>x"4700",
---- 737=>x"3700", 738=>x"4700", 739=>x"5100", 740=>x"4500",
---- 741=>x"3700", 742=>x"3b00", 743=>x"4700", 744=>x"4600",
---- 745=>x"3a00", 746=>x"3500", 747=>x"4600", 748=>x"3e00",
---- 749=>x"3800", 750=>x"3200", 751=>x"4900", 752=>x"3e00",
---- 753=>x"3e00", 754=>x"3400", 755=>x"4500", 756=>x"3800",
---- 757=>x"4300", 758=>x"3600", 759=>x"3d00", 760=>x"3900",
---- 761=>x"4400", 762=>x"3700", 763=>x"3900", 764=>x"3c00",
---- 765=>x"3f00", 766=>x"3600", 767=>x"3900", 768=>x"4000",
---- 769=>x"3f00", 770=>x"3b00", 771=>x"3700", 772=>x"4200",
---- 773=>x"4100", 774=>x"3e00", 775=>x"3600", 776=>x"3b00",
---- 777=>x"3b00", 778=>x"3d00", 779=>x"3500", 780=>x"3b00",
---- 781=>x"3a00", 782=>x"3600", 783=>x"3300", 784=>x"3700",
---- 785=>x"3f00", 786=>x"3500", 787=>x"3200", 788=>x"3900",
---- 789=>x"3900", 790=>x"3400", 791=>x"3900", 792=>x"3900",
---- 793=>x"3b00", 794=>x"3b00", 795=>x"3600", 796=>x"3a00",
---- 797=>x"3a00", 798=>x"3a00", 799=>x"3800", 800=>x"3b00",
---- 801=>x"4300", 802=>x"4000", 803=>x"3700", 804=>x"3f00",
---- 805=>x"4800", 806=>x"4400", 807=>x"3900", 808=>x"3c00",
---- 809=>x"4100", 810=>x"5000", 811=>x"4000", 812=>x"4000",
---- 813=>x"3c00", 814=>x"5200", 815=>x"4600", 816=>x"4300",
---- 817=>x"4100", 818=>x"5600", 819=>x"5400", 820=>x"3e00",
---- 821=>x"4600", 822=>x"5a00", 823=>x"6200", 824=>x"3e00",
---- 825=>x"4900", 826=>x"6000", 827=>x"6a00", 828=>x"4000",
---- 829=>x"4b00", 830=>x"6700", 831=>x"6e00", 832=>x"4100",
---- 833=>x"4c00", 834=>x"6d00", 835=>x"7700", 836=>x"3d00",
---- 837=>x"5800", 838=>x"7400", 839=>x"7600", 840=>x"3a00",
---- 841=>x"5d00", 842=>x"7500", 843=>x"7800", 844=>x"4400",
---- 845=>x"6700", 846=>x"7500", 847=>x"7600", 848=>x"4e00",
---- 849=>x"6500", 850=>x"6c00", 851=>x"7200", 852=>x"5600",
---- 853=>x"6a00", 854=>x"6f00", 855=>x"6700", 856=>x"6300",
---- 857=>x"7100", 858=>x"6500", 859=>x"6200", 860=>x"5f00",
---- 861=>x"6300", 862=>x"6300", 863=>x"7300", 864=>x"6200",
---- 865=>x"6c00", 866=>x"7600", 867=>x"7b00", 868=>x"7200",
---- 869=>x"7800", 870=>x"7b00", 871=>x"7d00", 872=>x"7900",
---- 873=>x"7b00", 874=>x"7d00", 875=>x"7a00", 876=>x"7c00",
---- 877=>x"7d00", 878=>x"7b00", 879=>x"7800", 880=>x"7e00",
---- 881=>x"7d00", 882=>x"7b00", 883=>x"7c00", 884=>x"7d00",
---- 885=>x"7c00", 886=>x"7d00", 887=>x"7b00", 888=>x"7c00",
---- 889=>x"7a00", 890=>x"8000", 891=>x"7f00", 892=>x"7c00",
---- 893=>x"8000", 894=>x"8100", 895=>x"8100", 896=>x"8100",
---- 897=>x"7f00", 898=>x"8100", 899=>x"8300", 900=>x"7e00",
---- 901=>x"8100", 902=>x"8100", 903=>x"7e00", 904=>x"7d00",
---- 905=>x"8100", 906=>x"8000", 907=>x"7800", 908=>x"7f00",
---- 909=>x"7d00", 910=>x"7d00", 911=>x"7300", 912=>x"7d00",
---- 913=>x"7c00", 914=>x"7b00", 915=>x"6300", 916=>x"7b00",
---- 917=>x"7b00", 918=>x"7700", 919=>x"4e00", 920=>x"7b00",
---- 921=>x"7d00", 922=>x"6900", 923=>x"3c00", 924=>x"7c00",
---- 925=>x"7a00", 926=>x"5900", 927=>x"3200", 928=>x"7b00",
---- 929=>x"6c00", 930=>x"3800", 931=>x"3100", 932=>x"7700",
---- 933=>x"4d00", 934=>x"2900", 935=>x"4000", 936=>x"6100",
---- 937=>x"3000", 938=>x"2800", 939=>x"4a00", 940=>x"3900",
---- 941=>x"2200", 942=>x"3900", 943=>x"5a00", 944=>x"2700",
---- 945=>x"2a00", 946=>x"4c00", 947=>x"6600", 948=>x"2900",
---- 949=>x"3e00", 950=>x"5d00", 951=>x"7800", 952=>x"2e00",
---- 953=>x"5300", 954=>x"7100", 955=>x"8100", 956=>x"4900",
---- 957=>x"6600", 958=>x"7c00", 959=>x"8100", 960=>x"6400",
---- 961=>x"7a00", 962=>x"7f00", 963=>x"7f00", 964=>x"7200",
---- 965=>x"7b00", 966=>x"7d00", 967=>x"8100", 968=>x"7a00",
---- 969=>x"7c00", 970=>x"7f00", 971=>x"7f00", 972=>x"7a00",
---- 973=>x"7c00", 974=>x"7f00", 975=>x"8300", 976=>x"7d00",
---- 977=>x"7d00", 978=>x"8000", 979=>x"8300", 980=>x"7a00",
---- 981=>x"7d00", 982=>x"8300", 983=>x"8200", 984=>x"8000",
---- 985=>x"7f00", 986=>x"8000", 987=>x"7e00", 988=>x"7f00",
---- 989=>x"8000", 990=>x"8000", 991=>x"8100", 992=>x"8200",
---- 993=>x"8300", 994=>x"7d00", 995=>x"8000", 996=>x"7f00",
---- 997=>x"8100", 998=>x"8000", 999=>x"8000", 1000=>x"8000",
---- 1001=>x"8100", 1002=>x"8000", 1003=>x"8100", 1004=>x"8000",
---- 1005=>x"8100", 1006=>x"8000", 1007=>x"8500", 1008=>x"8000",
---- 1009=>x"8300", 1010=>x"8300", 1011=>x"8300", 1012=>x"8100",
---- 1013=>x"8400", 1014=>x"8300", 1015=>x"8200", 1016=>x"8000",
---- 1017=>x"8200", 1018=>x"8000", 1019=>x"8200", 1020=>x"7e00",
---- 1021=>x"8000", 1022=>x"8100", 1023=>x"8400"),
----
---- 29 => (0=>x"8400", 1=>x"8400", 2=>x"8300", 3=>x"8400", 4=>x"8400",
---- 5=>x"8400", 6=>x"8300", 7=>x"8400", 8=>x"8200",
---- 9=>x"8300", 10=>x"8200", 11=>x"8300", 12=>x"8100",
---- 13=>x"8000", 14=>x"7e00", 15=>x"8400", 16=>x"8200",
---- 17=>x"8000", 18=>x"8100", 19=>x"8400", 20=>x"8000",
---- 21=>x"8100", 22=>x"8200", 23=>x"8100", 24=>x"8100",
---- 25=>x"8000", 26=>x"8200", 27=>x"8300", 28=>x"8000",
---- 29=>x"7f00", 30=>x"8300", 31=>x"8200", 32=>x"8100",
---- 33=>x"8100", 34=>x"8200", 35=>x"8300", 36=>x"8100",
---- 37=>x"7f00", 38=>x"8100", 39=>x"8400", 40=>x"8000",
---- 41=>x"7f00", 42=>x"8000", 43=>x"8200", 44=>x"8000",
---- 45=>x"7f00", 46=>x"8000", 47=>x"8000", 48=>x"8000",
---- 49=>x"7e00", 50=>x"7d00", 51=>x"8000", 52=>x"8000",
---- 53=>x"7d00", 54=>x"7c00", 55=>x"7e00", 56=>x"8300",
---- 57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7c00",
---- 61=>x"7b00", 62=>x"7e00", 63=>x"7f00", 64=>x"7e00",
---- 65=>x"7e00", 66=>x"7c00", 67=>x"7c00", 68=>x"7a00",
---- 69=>x"7c00", 70=>x"7a00", 71=>x"7c00", 72=>x"7a00",
---- 73=>x"7700", 74=>x"7700", 75=>x"7c00", 76=>x"7800",
---- 77=>x"7600", 78=>x"7900", 79=>x"7900", 80=>x"7900",
---- 81=>x"7700", 82=>x"7900", 83=>x"7800", 84=>x"7400",
---- 85=>x"7700", 86=>x"7500", 87=>x"7500", 88=>x"7d00",
---- 89=>x"7b00", 90=>x"7400", 91=>x"7200", 92=>x"aa00",
---- 93=>x"ab00", 94=>x"a300", 95=>x"9f00", 96=>x"b700",
---- 97=>x"b800", 98=>x"bc00", 99=>x"bc00", 100=>x"b000",
---- 101=>x"b800", 102=>x"b100", 103=>x"b400", 104=>x"b300",
---- 105=>x"ae00", 106=>x"a700", 107=>x"aa00", 108=>x"b000",
---- 109=>x"ac00", 110=>x"ac00", 111=>x"ac00", 112=>x"b000",
---- 113=>x"b300", 114=>x"b100", 115=>x"af00", 116=>x"a700",
---- 117=>x"af00", 118=>x"4b00", 119=>x"b100", 120=>x"aa00",
---- 121=>x"b200", 122=>x"b400", 123=>x"b100", 124=>x"af00",
---- 125=>x"b500", 126=>x"b400", 127=>x"b200", 128=>x"ac00",
---- 129=>x"b000", 130=>x"b600", 131=>x"bd00", 132=>x"ae00",
---- 133=>x"b100", 134=>x"b800", 135=>x"ba00", 136=>x"5000",
---- 137=>x"b200", 138=>x"b400", 139=>x"b400", 140=>x"ae00",
---- 141=>x"af00", 142=>x"b500", 143=>x"ae00", 144=>x"ab00",
---- 145=>x"ae00", 146=>x"b300", 147=>x"b600", 148=>x"a800",
---- 149=>x"af00", 150=>x"b600", 151=>x"b500", 152=>x"ac00",
---- 153=>x"b300", 154=>x"b500", 155=>x"b300", 156=>x"ae00",
---- 157=>x"4900", 158=>x"b600", 159=>x"b900", 160=>x"b000",
---- 161=>x"b500", 162=>x"be00", 163=>x"bc00", 164=>x"b300",
---- 165=>x"be00", 166=>x"b300", 167=>x"b400", 168=>x"ac00",
---- 169=>x"b600", 170=>x"ba00", 171=>x"ba00", 172=>x"b000",
---- 173=>x"bc00", 174=>x"af00", 175=>x"b200", 176=>x"a700",
---- 177=>x"ad00", 178=>x"b700", 179=>x"b600", 180=>x"ab00",
---- 181=>x"b700", 182=>x"b100", 183=>x"b000", 184=>x"ae00",
---- 185=>x"4f00", 186=>x"b500", 187=>x"b200", 188=>x"af00",
---- 189=>x"af00", 190=>x"ab00", 191=>x"9a00", 192=>x"b200",
---- 193=>x"9b00", 194=>x"8800", 195=>x"9300", 196=>x"9100",
---- 197=>x"7e00", 198=>x"9800", 199=>x"ba00", 200=>x"8500",
---- 201=>x"a500", 202=>x"c700", 203=>x"c100", 204=>x"b200",
---- 205=>x"c600", 206=>x"c700", 207=>x"3a00", 208=>x"c200",
---- 209=>x"be00", 210=>x"c600", 211=>x"c600", 212=>x"b500",
---- 213=>x"c500", 214=>x"c500", 215=>x"ca00", 216=>x"bc00",
---- 217=>x"c000", 218=>x"c300", 219=>x"c100", 220=>x"bf00",
---- 221=>x"b700", 222=>x"bb00", 223=>x"b900", 224=>x"b500",
---- 225=>x"b900", 226=>x"b400", 227=>x"bd00", 228=>x"bd00",
---- 229=>x"bb00", 230=>x"c100", 231=>x"b800", 232=>x"be00",
---- 233=>x"c400", 234=>x"bf00", 235=>x"af00", 236=>x"b700",
---- 237=>x"b100", 238=>x"ad00", 239=>x"b800", 240=>x"a000",
---- 241=>x"a300", 242=>x"b900", 243=>x"bd00", 244=>x"b100",
---- 245=>x"b700", 246=>x"b000", 247=>x"b400", 248=>x"bb00",
---- 249=>x"b200", 250=>x"ae00", 251=>x"a800", 252=>x"b800",
---- 253=>x"b200", 254=>x"af00", 255=>x"b500", 256=>x"ae00",
---- 257=>x"b400", 258=>x"be00", 259=>x"bd00", 260=>x"b300",
---- 261=>x"ba00", 262=>x"bd00", 263=>x"b900", 264=>x"b400",
---- 265=>x"b100", 266=>x"b500", 267=>x"bd00", 268=>x"b300",
---- 269=>x"a900", 270=>x"af00", 271=>x"b200", 272=>x"b500",
---- 273=>x"b200", 274=>x"a800", 275=>x"b400", 276=>x"a800",
---- 277=>x"b900", 278=>x"bb00", 279=>x"b000", 280=>x"b400",
---- 281=>x"b700", 282=>x"bc00", 283=>x"bb00", 284=>x"a500",
---- 285=>x"b700", 286=>x"b200", 287=>x"af00", 288=>x"ac00",
---- 289=>x"9f00", 290=>x"a400", 291=>x"9600", 292=>x"b200",
---- 293=>x"9a00", 294=>x"6300", 295=>x"ac00", 296=>x"9700",
---- 297=>x"9b00", 298=>x"ad00", 299=>x"ba00", 300=>x"a400",
---- 301=>x"b100", 302=>x"a600", 303=>x"ae00", 304=>x"b500",
---- 305=>x"b300", 306=>x"ae00", 307=>x"a100", 308=>x"b200",
---- 309=>x"b000", 310=>x"ab00", 311=>x"a700", 312=>x"a700",
---- 313=>x"a500", 314=>x"aa00", 315=>x"a900", 316=>x"a500",
---- 317=>x"a200", 318=>x"a500", 319=>x"a900", 320=>x"ab00",
---- 321=>x"a800", 322=>x"a200", 323=>x"a700", 324=>x"a200",
---- 325=>x"b100", 326=>x"ac00", 327=>x"9e00", 328=>x"a200",
---- 329=>x"a200", 330=>x"a900", 331=>x"9d00", 332=>x"9900",
---- 333=>x"9b00", 334=>x"9300", 335=>x"9100", 336=>x"9c00",
---- 337=>x"9d00", 338=>x"9400", 339=>x"8c00", 340=>x"9a00",
---- 341=>x"9900", 342=>x"9300", 343=>x"8500", 344=>x"6c00",
---- 345=>x"8700", 346=>x"9700", 347=>x"7400", 348=>x"6300",
---- 349=>x"5900", 350=>x"6700", 351=>x"6200", 352=>x"6b00",
---- 353=>x"5d00", 354=>x"4500", 355=>x"5300", 356=>x"4300",
---- 357=>x"4800", 358=>x"3f00", 359=>x"4a00", 360=>x"6600",
---- 361=>x"5200", 362=>x"5000", 363=>x"6700", 364=>x"7e00",
---- 365=>x"6700", 366=>x"5100", 367=>x"5e00", 368=>x"5d00",
---- 369=>x"4500", 370=>x"4500", 371=>x"4e00", 372=>x"3900",
---- 373=>x"3900", 374=>x"3700", 375=>x"3a00", 376=>x"3600",
---- 377=>x"3c00", 378=>x"3b00", 379=>x"3b00", 380=>x"3300",
---- 381=>x"3500", 382=>x"3300", 383=>x"5200", 384=>x"3700",
---- 385=>x"2d00", 386=>x"3e00", 387=>x"7a00", 388=>x"3400",
---- 389=>x"2b00", 390=>x"5700", 391=>x"7c00", 392=>x"3100",
---- 393=>x"3a00", 394=>x"7c00", 395=>x"6500", 396=>x"3700",
---- 397=>x"5c00", 398=>x"8d00", 399=>x"4000", 400=>x"4a00",
---- 401=>x"5b00", 402=>x"5900", 403=>x"2f00", 404=>x"5d00",
---- 405=>x"5000", 406=>x"4500", 407=>x"2700", 408=>x"6100",
---- 409=>x"4b00", 410=>x"3900", 411=>x"2c00", 412=>x"5300",
---- 413=>x"4b00", 414=>x"3b00", 415=>x"2a00", 416=>x"3400",
---- 417=>x"3900", 418=>x"3900", 419=>x"3b00", 420=>x"2e00",
---- 421=>x"3200", 422=>x"3200", 423=>x"3800", 424=>x"2f00",
---- 425=>x"2f00", 426=>x"2f00", 427=>x"3100", 428=>x"3200",
---- 429=>x"2e00", 430=>x"3000", 431=>x"3100", 432=>x"3200",
---- 433=>x"3100", 434=>x"3000", 435=>x"2c00", 436=>x"2900",
---- 437=>x"2e00", 438=>x"2d00", 439=>x"2a00", 440=>x"5700",
---- 441=>x"3c00", 442=>x"2400", 443=>x"2700", 444=>x"4d00",
---- 445=>x"3e00", 446=>x"2700", 447=>x"2400", 448=>x"2500",
---- 449=>x"2400", 450=>x"2300", 451=>x"2200", 452=>x"2700",
---- 453=>x"2300", 454=>x"2300", 455=>x"1d00", 456=>x"1f00",
---- 457=>x"2100", 458=>x"2000", 459=>x"3600", 460=>x"1e00",
---- 461=>x"1c00", 462=>x"2e00", 463=>x"7f00", 464=>x"1700",
---- 465=>x"2500", 466=>x"7000", 467=>x"9e00", 468=>x"2200",
---- 469=>x"5d00", 470=>x"9c00", 471=>x"7e00", 472=>x"6400",
---- 473=>x"9500", 474=>x"8900", 475=>x"9400", 476=>x"8c00",
---- 477=>x"8800", 478=>x"6c00", 479=>x"8700", 480=>x"7700",
---- 481=>x"5a00", 482=>x"7a00", 483=>x"b100", 484=>x"5d00",
---- 485=>x"6a00", 486=>x"b300", 487=>x"ae00", 488=>x"5d00",
---- 489=>x"a900", 490=>x"bb00", 491=>x"a300", 492=>x"9200",
---- 493=>x"bc00", 494=>x"a700", 495=>x"ac00", 496=>x"b600",
---- 497=>x"a800", 498=>x"ad00", 499=>x"b400", 500=>x"ab00",
---- 501=>x"a700", 502=>x"b400", 503=>x"4200", 504=>x"a400",
---- 505=>x"af00", 506=>x"b700", 507=>x"c400", 508=>x"ac00",
---- 509=>x"b600", 510=>x"bf00", 511=>x"c700", 512=>x"b400",
---- 513=>x"c000", 514=>x"c900", 515=>x"c700", 516=>x"bb00",
---- 517=>x"c700", 518=>x"ca00", 519=>x"c100", 520=>x"bc00",
---- 521=>x"c900", 522=>x"c500", 523=>x"bf00", 524=>x"c100",
---- 525=>x"cc00", 526=>x"c500", 527=>x"be00", 528=>x"c700",
---- 529=>x"ca00", 530=>x"c300", 531=>x"c500", 532=>x"cd00",
---- 533=>x"c700", 534=>x"c700", 535=>x"cc00", 536=>x"c800",
---- 537=>x"c300", 538=>x"cc00", 539=>x"9300", 540=>x"c300",
---- 541=>x"ca00", 542=>x"9600", 543=>x"6500", 544=>x"c600",
---- 545=>x"9700", 546=>x"6900", 547=>x"7800", 548=>x"7100",
---- 549=>x"6200", 550=>x"7a00", 551=>x"7e00", 552=>x"5b00",
---- 553=>x"7200", 554=>x"7e00", 555=>x"7f00", 556=>x"6b00",
---- 557=>x"7a00", 558=>x"8200", 559=>x"8700", 560=>x"7200",
---- 561=>x"7e00", 562=>x"8300", 563=>x"8800", 564=>x"7700",
---- 565=>x"7f00", 566=>x"8600", 567=>x"8c00", 568=>x"7600",
---- 569=>x"8000", 570=>x"8600", 571=>x"8b00", 572=>x"7900",
---- 573=>x"8400", 574=>x"8700", 575=>x"8900", 576=>x"7c00",
---- 577=>x"7d00", 578=>x"8900", 579=>x"8b00", 580=>x"7d00",
---- 581=>x"8100", 582=>x"8400", 583=>x"8b00", 584=>x"7e00",
---- 585=>x"8000", 586=>x"8400", 587=>x"8c00", 588=>x"7d00",
---- 589=>x"8000", 590=>x"8500", 591=>x"8a00", 592=>x"7c00",
---- 593=>x"7c00", 594=>x"8300", 595=>x"8b00", 596=>x"8000",
---- 597=>x"7d00", 598=>x"8400", 599=>x"8600", 600=>x"8000",
---- 601=>x"8500", 602=>x"8500", 603=>x"8300", 604=>x"7d00",
---- 605=>x"8300", 606=>x"8400", 607=>x"8800", 608=>x"8000",
---- 609=>x"8000", 610=>x"8400", 611=>x"8800", 612=>x"8100",
---- 613=>x"8100", 614=>x"8500", 615=>x"7a00", 616=>x"7e00",
---- 617=>x"7e00", 618=>x"8200", 619=>x"8300", 620=>x"7c00",
---- 621=>x"7f00", 622=>x"8300", 623=>x"8300", 624=>x"7d00",
---- 625=>x"8100", 626=>x"8100", 627=>x"8500", 628=>x"7e00",
---- 629=>x"8000", 630=>x"8200", 631=>x"8500", 632=>x"7c00",
---- 633=>x"7e00", 634=>x"8000", 635=>x"8300", 636=>x"7c00",
---- 637=>x"8000", 638=>x"8000", 639=>x"8200", 640=>x"7e00",
---- 641=>x"8000", 642=>x"8200", 643=>x"8000", 644=>x"7b00",
---- 645=>x"7c00", 646=>x"8100", 647=>x"8000", 648=>x"7800",
---- 649=>x"7c00", 650=>x"8000", 651=>x"8200", 652=>x"7c00",
---- 653=>x"7a00", 654=>x"7f00", 655=>x"8200", 656=>x"7d00",
---- 657=>x"7c00", 658=>x"7d00", 659=>x"8300", 660=>x"7b00",
---- 661=>x"7d00", 662=>x"7f00", 663=>x"8200", 664=>x"7b00",
---- 665=>x"7c00", 666=>x"7a00", 667=>x"7f00", 668=>x"7d00",
---- 669=>x"7e00", 670=>x"7f00", 671=>x"8100", 672=>x"7d00",
---- 673=>x"7f00", 674=>x"8000", 675=>x"7f00", 676=>x"7d00",
---- 677=>x"7e00", 678=>x"8200", 679=>x"8200", 680=>x"7d00",
---- 681=>x"8100", 682=>x"8100", 683=>x"8200", 684=>x"7c00",
---- 685=>x"8000", 686=>x"7d00", 687=>x"8000", 688=>x"7b00",
---- 689=>x"7f00", 690=>x"7f00", 691=>x"8200", 692=>x"7c00",
---- 693=>x"7d00", 694=>x"8200", 695=>x"8200", 696=>x"7900",
---- 697=>x"8000", 698=>x"8300", 699=>x"8100", 700=>x"7700",
---- 701=>x"7e00", 702=>x"8500", 703=>x"8100", 704=>x"7900",
---- 705=>x"7b00", 706=>x"7f00", 707=>x"7f00", 708=>x"7500",
---- 709=>x"7800", 710=>x"7d00", 711=>x"7c00", 712=>x"7300",
---- 713=>x"7300", 714=>x"7700", 715=>x"7a00", 716=>x"6e00",
---- 717=>x"7100", 718=>x"7400", 719=>x"7500", 720=>x"6b00",
---- 721=>x"6f00", 722=>x"7400", 723=>x"8c00", 724=>x"6800",
---- 725=>x"6900", 726=>x"6a00", 727=>x"6e00", 728=>x"5f00",
---- 729=>x"6900", 730=>x"6900", 731=>x"6900", 732=>x"5600",
---- 733=>x"9d00", 734=>x"6700", 735=>x"6600", 736=>x"5400",
---- 737=>x"5900", 738=>x"5d00", 739=>x"6600", 740=>x"4600",
---- 741=>x"5600", 742=>x"5900", 743=>x"6100", 744=>x"4000",
---- 745=>x"4700", 746=>x"5300", 747=>x"5b00", 748=>x"4600",
---- 749=>x"3300", 750=>x"3f00", 751=>x"5000", 752=>x"4b00",
---- 753=>x"3500", 754=>x"3000", 755=>x"3d00", 756=>x"4c00",
---- 757=>x"3d00", 758=>x"2e00", 759=>x"2e00", 760=>x"4800",
---- 761=>x"4500", 762=>x"3500", 763=>x"2d00", 764=>x"4a00",
---- 765=>x"4a00", 766=>x"4200", 767=>x"3300", 768=>x"bb00",
---- 769=>x"4900", 770=>x"4800", 771=>x"3d00", 772=>x"3d00",
---- 773=>x"4600", 774=>x"5100", 775=>x"5000", 776=>x"3400",
---- 777=>x"4000", 778=>x"b300", 779=>x"5000", 780=>x"2e00",
---- 781=>x"3900", 782=>x"4600", 783=>x"4e00", 784=>x"3200",
---- 785=>x"3400", 786=>x"4900", 787=>x"5100", 788=>x"3400",
---- 789=>x"3500", 790=>x"4900", 791=>x"5500", 792=>x"3600",
---- 793=>x"3200", 794=>x"4300", 795=>x"5300", 796=>x"3800",
---- 797=>x"2f00", 798=>x"3f00", 799=>x"5200", 800=>x"3600",
---- 801=>x"2e00", 802=>x"3800", 803=>x"4d00", 804=>x"3900",
---- 805=>x"3200", 806=>x"3800", 807=>x"4900", 808=>x"3900",
---- 809=>x"3300", 810=>x"3800", 811=>x"4d00", 812=>x"3400",
---- 813=>x"3900", 814=>x"3600", 815=>x"4e00", 816=>x"3800",
---- 817=>x"3300", 818=>x"3400", 819=>x"5000", 820=>x"4400",
---- 821=>x"2e00", 822=>x"2b00", 823=>x"4800", 824=>x"5400",
---- 825=>x"3400", 826=>x"2d00", 827=>x"3d00", 828=>x"5c00",
---- 829=>x"3800", 830=>x"2b00", 831=>x"3d00", 832=>x"6700",
---- 833=>x"3f00", 834=>x"2900", 835=>x"3600", 836=>x"6b00",
---- 837=>x"4800", 838=>x"2a00", 839=>x"3600", 840=>x"6f00",
---- 841=>x"5000", 842=>x"2800", 843=>x"2f00", 844=>x"6e00",
---- 845=>x"4e00", 846=>x"2900", 847=>x"2b00", 848=>x"9200",
---- 849=>x"5000", 850=>x"2b00", 851=>x"2d00", 852=>x"9b00",
---- 853=>x"5a00", 854=>x"3200", 855=>x"2f00", 856=>x"7000",
---- 857=>x"6000", 858=>x"3200", 859=>x"2f00", 860=>x"7b00",
---- 861=>x"6000", 862=>x"3400", 863=>x"3000", 864=>x"7800",
---- 865=>x"6400", 866=>x"3200", 867=>x"3200", 868=>x"7800",
---- 869=>x"6800", 870=>x"3100", 871=>x"3900", 872=>x"7a00",
---- 873=>x"6000", 874=>x"3200", 875=>x"4200", 876=>x"7600",
---- 877=>x"5700", 878=>x"2d00", 879=>x"4800", 880=>x"7700",
---- 881=>x"4f00", 882=>x"2d00", 883=>x"4b00", 884=>x"7a00",
---- 885=>x"4900", 886=>x"2e00", 887=>x"4e00", 888=>x"7300",
---- 889=>x"4a00", 890=>x"3400", 891=>x"5500", 892=>x"6e00",
---- 893=>x"4300", 894=>x"3a00", 895=>x"5a00", 896=>x"6800",
---- 897=>x"3a00", 898=>x"4200", 899=>x"5f00", 900=>x"5d00",
---- 901=>x"3700", 902=>x"4b00", 903=>x"6500", 904=>x"4f00",
---- 905=>x"3400", 906=>x"5100", 907=>x"6500", 908=>x"4200",
---- 909=>x"3a00", 910=>x"5a00", 911=>x"6500", 912=>x"3700",
---- 913=>x"4200", 914=>x"6000", 915=>x"6b00", 916=>x"3200",
---- 917=>x"5300", 918=>x"6100", 919=>x"7400", 920=>x"3700",
---- 921=>x"5700", 922=>x"6700", 923=>x"7e00", 924=>x"4100",
---- 925=>x"5a00", 926=>x"7000", 927=>x"8800", 928=>x"5100",
---- 929=>x"6000", 930=>x"7c00", 931=>x"8300", 932=>x"5a00",
---- 933=>x"6c00", 934=>x"8100", 935=>x"8500", 936=>x"6800",
---- 937=>x"7700", 938=>x"8400", 939=>x"8700", 940=>x"6f00",
---- 941=>x"8100", 942=>x"8600", 943=>x"8700", 944=>x"7b00",
---- 945=>x"8300", 946=>x"8400", 947=>x"8900", 948=>x"8200",
---- 949=>x"8100", 950=>x"8600", 951=>x"8a00", 952=>x"8100",
---- 953=>x"8200", 954=>x"8900", 955=>x"8600", 956=>x"8100",
---- 957=>x"8500", 958=>x"8800", 959=>x"8600", 960=>x"8300",
---- 961=>x"8400", 962=>x"8600", 963=>x"8800", 964=>x"8400",
---- 965=>x"8100", 966=>x"8700", 967=>x"8700", 968=>x"8300",
---- 969=>x"8300", 970=>x"8700", 971=>x"8800", 972=>x"8400",
---- 973=>x"8500", 974=>x"8600", 975=>x"8900", 976=>x"8200",
---- 977=>x"8400", 978=>x"8800", 979=>x"8700", 980=>x"8400",
---- 981=>x"8100", 982=>x"8600", 983=>x"8800", 984=>x"8200",
---- 985=>x"8300", 986=>x"8500", 987=>x"8600", 988=>x"8200",
---- 989=>x"7f00", 990=>x"8200", 991=>x"8600", 992=>x"7e00",
---- 993=>x"7f00", 994=>x"8200", 995=>x"8700", 996=>x"8000",
---- 997=>x"8000", 998=>x"8700", 999=>x"8400", 1000=>x"8100",
---- 1001=>x"8100", 1002=>x"8700", 1003=>x"8400", 1004=>x"8500",
---- 1005=>x"8100", 1006=>x"8300", 1007=>x"8300", 1008=>x"8500",
---- 1009=>x"8300", 1010=>x"8200", 1011=>x"8400", 1012=>x"8400",
---- 1013=>x"8500", 1014=>x"8100", 1015=>x"8100", 1016=>x"8400",
---- 1017=>x"8300", 1018=>x"8200", 1019=>x"8200", 1020=>x"8300",
---- 1021=>x"8500", 1022=>x"8400", 1023=>x"8200"),
----
---- 30 => (0=>x"8600", 1=>x"8500", 2=>x"8500", 3=>x"8700", 4=>x"8600",
---- 5=>x"8400", 6=>x"8600", 7=>x"8800", 8=>x"8700",
---- 9=>x"8500", 10=>x"8500", 11=>x"8700", 12=>x"8400",
---- 13=>x"8500", 14=>x"8600", 15=>x"8200", 16=>x"8300",
---- 17=>x"8400", 18=>x"8300", 19=>x"8300", 20=>x"8200",
---- 21=>x"8100", 22=>x"8400", 23=>x"8400", 24=>x"8500",
---- 25=>x"8700", 26=>x"8800", 27=>x"8500", 28=>x"8400",
---- 29=>x"8600", 30=>x"8600", 31=>x"8600", 32=>x"8400",
---- 33=>x"8800", 34=>x"8500", 35=>x"8900", 36=>x"8600",
---- 37=>x"8800", 38=>x"8700", 39=>x"8800", 40=>x"8200",
---- 41=>x"8400", 42=>x"8700", 43=>x"8900", 44=>x"8300",
---- 45=>x"8300", 46=>x"8500", 47=>x"8600", 48=>x"8400",
---- 49=>x"8200", 50=>x"8200", 51=>x"8200", 52=>x"7c00",
---- 53=>x"8000", 54=>x"8000", 55=>x"8200", 56=>x"7f00",
---- 57=>x"8200", 58=>x"8100", 59=>x"7e00", 60=>x"7f00",
---- 61=>x"8200", 62=>x"8400", 63=>x"8100", 64=>x"7d00",
---- 65=>x"7e00", 66=>x"8300", 67=>x"8000", 68=>x"7b00",
---- 69=>x"7e00", 70=>x"8100", 71=>x"8000", 72=>x"7c00",
---- 73=>x"7c00", 74=>x"8200", 75=>x"8100", 76=>x"7d00",
---- 77=>x"7d00", 78=>x"7d00", 79=>x"7f00", 80=>x"7a00",
---- 81=>x"7900", 82=>x"7d00", 83=>x"8000", 84=>x"7800",
---- 85=>x"7800", 86=>x"7c00", 87=>x"7d00", 88=>x"7500",
---- 89=>x"7400", 90=>x"7900", 91=>x"7c00", 92=>x"8b00",
---- 93=>x"8300", 94=>x"7500", 95=>x"7300", 96=>x"bd00",
---- 97=>x"b100", 98=>x"a100", 99=>x"9900", 100=>x"b200",
---- 101=>x"b600", 102=>x"c300", 103=>x"c200", 104=>x"b100",
---- 105=>x"b700", 106=>x"b400", 107=>x"ba00", 108=>x"5000",
---- 109=>x"b600", 110=>x"b400", 111=>x"b600", 112=>x"b200",
---- 113=>x"b400", 114=>x"b400", 115=>x"b400", 116=>x"ad00",
---- 117=>x"b500", 118=>x"b700", 119=>x"ba00", 120=>x"5200",
---- 121=>x"b700", 122=>x"ba00", 123=>x"bb00", 124=>x"b700",
---- 125=>x"b900", 126=>x"b800", 127=>x"bc00", 128=>x"be00",
---- 129=>x"ba00", 130=>x"b600", 131=>x"b700", 132=>x"b300",
---- 133=>x"b900", 134=>x"bb00", 135=>x"b800", 136=>x"b500",
---- 137=>x"b900", 138=>x"bb00", 139=>x"b600", 140=>x"b000",
---- 141=>x"ba00", 142=>x"b400", 143=>x"b200", 144=>x"b900",
---- 145=>x"b500", 146=>x"b500", 147=>x"bc00", 148=>x"b700",
---- 149=>x"b700", 150=>x"bb00", 151=>x"bc00", 152=>x"b800",
---- 153=>x"b800", 154=>x"bc00", 155=>x"b900", 156=>x"bd00",
---- 157=>x"be00", 158=>x"b300", 159=>x"bc00", 160=>x"b600",
---- 161=>x"ba00", 162=>x"bb00", 163=>x"b700", 164=>x"bc00",
---- 165=>x"bb00", 166=>x"b400", 167=>x"bc00", 168=>x"bb00",
---- 169=>x"b800", 170=>x"3c00", 171=>x"c100", 172=>x"4400",
---- 173=>x"ba00", 174=>x"bb00", 175=>x"c000", 176=>x"af00",
---- 177=>x"b700", 178=>x"bc00", 179=>x"b300", 180=>x"b600",
---- 181=>x"bd00", 182=>x"a000", 183=>x"9700", 184=>x"a700",
---- 185=>x"9d00", 186=>x"9900", 187=>x"b700", 188=>x"8d00",
---- 189=>x"9d00", 190=>x"bf00", 191=>x"d200", 192=>x"aa00",
---- 193=>x"c700", 194=>x"cb00", 195=>x"cb00", 196=>x"c400",
---- 197=>x"c400", 198=>x"cb00", 199=>x"c900", 200=>x"c000",
---- 201=>x"c200", 202=>x"c100", 203=>x"cc00", 204=>x"bf00",
---- 205=>x"c200", 206=>x"c700", 207=>x"c000", 208=>x"c800",
---- 209=>x"be00", 210=>x"c300", 211=>x"c200", 212=>x"c100",
---- 213=>x"c200", 214=>x"bb00", 215=>x"c300", 216=>x"be00",
---- 217=>x"bf00", 218=>x"c300", 219=>x"b900", 220=>x"c000",
---- 221=>x"c200", 222=>x"c200", 223=>x"c100", 224=>x"c100",
---- 225=>x"be00", 226=>x"b500", 227=>x"ac00", 228=>x"af00",
---- 229=>x"a700", 230=>x"b200", 231=>x"bc00", 232=>x"a800",
---- 233=>x"b800", 234=>x"ba00", 235=>x"bf00", 236=>x"c100",
---- 237=>x"be00", 238=>x"bc00", 239=>x"b700", 240=>x"bd00",
---- 241=>x"b600", 242=>x"b900", 243=>x"bc00", 244=>x"b600",
---- 245=>x"bc00", 246=>x"bf00", 247=>x"bc00", 248=>x"bc00",
---- 249=>x"bf00", 250=>x"c200", 251=>x"bd00", 252=>x"b800",
---- 253=>x"c500", 254=>x"bc00", 255=>x"c300", 256=>x"ba00",
---- 257=>x"b700", 258=>x"bd00", 259=>x"b700", 260=>x"b800",
---- 261=>x"b800", 262=>x"b500", 263=>x"b800", 264=>x"b900",
---- 265=>x"b600", 266=>x"b500", 267=>x"b300", 268=>x"b900",
---- 269=>x"b300", 270=>x"b400", 271=>x"b700", 272=>x"b300",
---- 273=>x"ba00", 274=>x"ba00", 275=>x"ab00", 276=>x"b300",
---- 277=>x"b100", 278=>x"ad00", 279=>x"a100", 280=>x"a800",
---- 281=>x"9b00", 282=>x"9f00", 283=>x"b800", 284=>x"9900",
---- 285=>x"9c00", 286=>x"b400", 287=>x"b500", 288=>x"a800",
---- 289=>x"b200", 290=>x"ad00", 291=>x"af00", 292=>x"b100",
---- 293=>x"b300", 294=>x"ae00", 295=>x"a600", 296=>x"b100",
---- 297=>x"a800", 298=>x"ae00", 299=>x"b000", 300=>x"b000",
---- 301=>x"a800", 302=>x"a800", 303=>x"af00", 304=>x"a100",
---- 305=>x"b000", 306=>x"ae00", 307=>x"ac00", 308=>x"a100",
---- 309=>x"a500", 310=>x"4d00", 311=>x"b100", 312=>x"a800",
---- 313=>x"a300", 314=>x"a100", 315=>x"aa00", 316=>x"a900",
---- 317=>x"ac00", 318=>x"a700", 319=>x"9f00", 320=>x"ac00",
---- 321=>x"a900", 322=>x"ab00", 323=>x"a200", 324=>x"a400",
---- 325=>x"9f00", 326=>x"9f00", 327=>x"a400", 328=>x"9b00",
---- 329=>x"6000", 330=>x"a000", 331=>x"a200", 332=>x"9700",
---- 333=>x"a600", 334=>x"a700", 335=>x"aa00", 336=>x"8300",
---- 337=>x"8300", 338=>x"8700", 339=>x"8400", 340=>x"8400",
---- 341=>x"8a00", 342=>x"8100", 343=>x"6700", 344=>x"8c00",
---- 345=>x"9600", 346=>x"9800", 347=>x"9100", 348=>x"8d00",
---- 349=>x"a200", 350=>x"a600", 351=>x"a200", 352=>x"9900",
---- 353=>x"ab00", 354=>x"a500", 355=>x"a700", 356=>x"9000",
---- 357=>x"9c00", 358=>x"a400", 359=>x"9e00", 360=>x"8200",
---- 361=>x"8a00", 362=>x"8d00", 363=>x"8a00", 364=>x"6b00",
---- 365=>x"5800", 366=>x"7400", 367=>x"8400", 368=>x"4b00",
---- 369=>x"5000", 370=>x"7300", 371=>x"6400", 372=>x"4200",
---- 373=>x"5e00", 374=>x"6400", 375=>x"7900", 376=>x"5b00",
---- 377=>x"6800", 378=>x"7300", 379=>x"7500", 380=>x"7b00",
---- 381=>x"6800", 382=>x"7400", 383=>x"5700", 384=>x"7c00",
---- 385=>x"7400", 386=>x"6100", 387=>x"3400", 388=>x"7000",
---- 389=>x"5f00", 390=>x"3600", 391=>x"3200", 392=>x"4c00",
---- 393=>x"4400", 394=>x"2b00", 395=>x"3200", 396=>x"3a00",
---- 397=>x"3700", 398=>x"3100", 399=>x"4600", 400=>x"3400",
---- 401=>x"3500", 402=>x"3700", 403=>x"6a00", 404=>x"2e00",
---- 405=>x"3800", 406=>x"3f00", 407=>x"5100", 408=>x"3b00",
---- 409=>x"3d00", 410=>x"3c00", 411=>x"3600", 412=>x"3e00",
---- 413=>x"2f00", 414=>x"3000", 415=>x"3400", 416=>x"4e00",
---- 417=>x"5500", 418=>x"4f00", 419=>x"5400", 420=>x"3d00",
---- 421=>x"4400", 422=>x"4a00", 423=>x"4300", 424=>x"3100",
---- 425=>x"2e00", 426=>x"2f00", 427=>x"2800", 428=>x"3600",
---- 429=>x"3100", 430=>x"2c00", 431=>x"2e00", 432=>x"2f00",
---- 433=>x"2f00", 434=>x"2600", 435=>x"2500", 436=>x"2800",
---- 437=>x"2400", 438=>x"2300", 439=>x"2500", 440=>x"2300",
---- 441=>x"2400", 442=>x"2100", 443=>x"a600", 444=>x"2100",
---- 445=>x"e200", 446=>x"5400", 447=>x"9d00", 448=>x"1900",
---- 449=>x"4200", 450=>x"a000", 451=>x"8e00", 452=>x"3b00",
---- 453=>x"9500", 454=>x"9400", 455=>x"6900", 456=>x"8a00",
---- 457=>x"9b00", 458=>x"7600", 459=>x"7e00", 460=>x"9a00",
---- 461=>x"7700", 462=>x"7800", 463=>x"af00", 464=>x"7800",
---- 465=>x"7300", 466=>x"a000", 467=>x"b400", 468=>x"7500",
---- 469=>x"9800", 470=>x"ac00", 471=>x"5c00", 472=>x"8e00",
---- 473=>x"b000", 474=>x"9f00", 475=>x"a200", 476=>x"b300",
---- 477=>x"a100", 478=>x"a000", 479=>x"a000", 480=>x"a500",
---- 481=>x"a100", 482=>x"a400", 483=>x"a100", 484=>x"a400",
---- 485=>x"ac00", 486=>x"ac00", 487=>x"a300", 488=>x"ad00",
---- 489=>x"b500", 490=>x"af00", 491=>x"9e00", 492=>x"b500",
---- 493=>x"c000", 494=>x"ac00", 495=>x"6600", 496=>x"bf00",
---- 497=>x"c100", 498=>x"a500", 499=>x"9700", 500=>x"c600",
---- 501=>x"b600", 502=>x"9800", 503=>x"9b00", 504=>x"c400",
---- 505=>x"a800", 506=>x"9700", 507=>x"a500", 508=>x"ba00",
---- 509=>x"a500", 510=>x"a200", 511=>x"b000", 512=>x"b800",
---- 513=>x"ac00", 514=>x"ae00", 515=>x"c300", 516=>x"b900",
---- 517=>x"b400", 518=>x"c100", 519=>x"c000", 520=>x"ba00",
---- 521=>x"be00", 522=>x"c100", 523=>x"6600", 524=>x"c200",
---- 525=>x"c200", 526=>x"6800", 527=>x"4400", 528=>x"c300",
---- 529=>x"7300", 530=>x"4900", 531=>x"5400", 532=>x"8200",
---- 533=>x"5300", 534=>x"5b00", 535=>x"4800", 536=>x"5e00",
---- 537=>x"7100", 538=>x"6900", 539=>x"5700", 540=>x"7200",
---- 541=>x"7d00", 542=>x"7d00", 543=>x"7400", 544=>x"7700",
---- 545=>x"7c00", 546=>x"8500", 547=>x"8900", 548=>x"7e00",
---- 549=>x"7d00", 550=>x"8500", 551=>x"9200", 552=>x"8600",
---- 553=>x"8300", 554=>x"8700", 555=>x"9100", 556=>x"8b00",
---- 557=>x"8b00", 558=>x"8c00", 559=>x"9000", 560=>x"9100",
---- 561=>x"8f00", 562=>x"9000", 563=>x"9400", 564=>x"9300",
---- 565=>x"6800", 566=>x"9900", 567=>x"9600", 568=>x"9600",
---- 569=>x"9900", 570=>x"9900", 571=>x"9700", 572=>x"9400",
---- 573=>x"9600", 574=>x"9a00", 575=>x"9d00", 576=>x"9100",
---- 577=>x"9600", 578=>x"9a00", 579=>x"9e00", 580=>x"8f00",
---- 581=>x"9700", 582=>x"9900", 583=>x"9d00", 584=>x"9000",
---- 585=>x"9600", 586=>x"9700", 587=>x"9b00", 588=>x"9100",
---- 589=>x"9400", 590=>x"9600", 591=>x"9b00", 592=>x"8f00",
---- 593=>x"9200", 594=>x"9800", 595=>x"9900", 596=>x"8800",
---- 597=>x"9100", 598=>x"9500", 599=>x"9300", 600=>x"8a00",
---- 601=>x"9100", 602=>x"9000", 603=>x"9200", 604=>x"8b00",
---- 605=>x"8f00", 606=>x"9300", 607=>x"9600", 608=>x"8c00",
---- 609=>x"8e00", 610=>x"9300", 611=>x"9700", 612=>x"8800",
---- 613=>x"8c00", 614=>x"9000", 615=>x"9400", 616=>x"8700",
---- 617=>x"8b00", 618=>x"8d00", 619=>x"9300", 620=>x"8a00",
---- 621=>x"8800", 622=>x"8b00", 623=>x"9500", 624=>x"8500",
---- 625=>x"8a00", 626=>x"8f00", 627=>x"8f00", 628=>x"8700",
---- 629=>x"8500", 630=>x"8a00", 631=>x"8c00", 632=>x"8700",
---- 633=>x"8a00", 634=>x"8b00", 635=>x"8f00", 636=>x"8400",
---- 637=>x"8800", 638=>x"8b00", 639=>x"8f00", 640=>x"8400",
---- 641=>x"8500", 642=>x"8d00", 643=>x"8b00", 644=>x"8400",
---- 645=>x"8900", 646=>x"8b00", 647=>x"8a00", 648=>x"8200",
---- 649=>x"8700", 650=>x"8800", 651=>x"8b00", 652=>x"8300",
---- 653=>x"8700", 654=>x"8800", 655=>x"8d00", 656=>x"8200",
---- 657=>x"8500", 658=>x"8800", 659=>x"8900", 660=>x"7f00",
---- 661=>x"8400", 662=>x"8600", 663=>x"8900", 664=>x"8200",
---- 665=>x"8200", 666=>x"8600", 667=>x"8800", 668=>x"8200",
---- 669=>x"8600", 670=>x"8b00", 671=>x"8b00", 672=>x"8200",
---- 673=>x"8500", 674=>x"8800", 675=>x"8a00", 676=>x"8100",
---- 677=>x"8400", 678=>x"8900", 679=>x"8800", 680=>x"8000",
---- 681=>x"8400", 682=>x"8800", 683=>x"8700", 684=>x"8100",
---- 685=>x"8600", 686=>x"8900", 687=>x"8900", 688=>x"8300",
---- 689=>x"8300", 690=>x"8800", 691=>x"8900", 692=>x"7f00",
---- 693=>x"8300", 694=>x"8600", 695=>x"8700", 696=>x"7c00",
---- 697=>x"8100", 698=>x"8300", 699=>x"8500", 700=>x"7d00",
---- 701=>x"7f00", 702=>x"8100", 703=>x"8200", 704=>x"7d00",
---- 705=>x"7d00", 706=>x"8100", 707=>x"8300", 708=>x"8600",
---- 709=>x"7e00", 710=>x"7f00", 711=>x"8000", 712=>x"7800",
---- 713=>x"7c00", 714=>x"7d00", 715=>x"7f00", 716=>x"7700",
---- 717=>x"7a00", 718=>x"7a00", 719=>x"7b00", 720=>x"7300",
---- 721=>x"7700", 722=>x"7800", 723=>x"7c00", 724=>x"7400",
---- 725=>x"7600", 726=>x"7800", 727=>x"7c00", 728=>x"6f00",
---- 729=>x"7300", 730=>x"7700", 731=>x"7700", 732=>x"6b00",
---- 733=>x"6900", 734=>x"7200", 735=>x"7400", 736=>x"6900",
---- 737=>x"6c00", 738=>x"6e00", 739=>x"7500", 740=>x"6800",
---- 741=>x"6a00", 742=>x"6f00", 743=>x"7100", 744=>x"6300",
---- 745=>x"6600", 746=>x"6b00", 747=>x"6e00", 748=>x"5600",
---- 749=>x"5c00", 750=>x"6600", 751=>x"6800", 752=>x"4800",
---- 753=>x"5300", 754=>x"5e00", 755=>x"5e00", 756=>x"3500",
---- 757=>x"4300", 758=>x"5100", 759=>x"5800", 760=>x"2c00",
---- 761=>x"3600", 762=>x"3f00", 763=>x"4c00", 764=>x"3000",
---- 765=>x"2c00", 766=>x"3200", 767=>x"3a00", 768=>x"3700",
---- 769=>x"3600", 770=>x"3100", 771=>x"3800", 772=>x"3f00",
---- 773=>x"3c00", 774=>x"3d00", 775=>x"4500", 776=>x"4900",
---- 777=>x"4b00", 778=>x"5400", 779=>x"6600", 780=>x"5400",
---- 781=>x"5a00", 782=>x"6a00", 783=>x"6e00", 784=>x"5400",
---- 785=>x"6300", 786=>x"6f00", 787=>x"8900", 788=>x"5700",
---- 789=>x"6600", 790=>x"7500", 791=>x"7b00", 792=>x"5b00",
---- 793=>x"6b00", 794=>x"7300", 795=>x"7900", 796=>x"5900",
---- 797=>x"6b00", 798=>x"7900", 799=>x"7900", 800=>x"5a00",
---- 801=>x"6700", 802=>x"7300", 803=>x"7400", 804=>x"5e00",
---- 805=>x"6700", 806=>x"6f00", 807=>x"7000", 808=>x"5900",
---- 809=>x"6500", 810=>x"7100", 811=>x"7400", 812=>x"5a00",
---- 813=>x"6500", 814=>x"7100", 815=>x"7500", 816=>x"5500",
---- 817=>x"6800", 818=>x"7100", 819=>x"7400", 820=>x"5300",
---- 821=>x"6b00", 822=>x"7400", 823=>x"7200", 824=>x"5200",
---- 825=>x"6e00", 826=>x"7900", 827=>x"7800", 828=>x"5200",
---- 829=>x"7000", 830=>x"7b00", 831=>x"7b00", 832=>x"5200",
---- 833=>x"6800", 834=>x"7b00", 835=>x"7100", 836=>x"5200",
---- 837=>x"6200", 838=>x"6f00", 839=>x"6c00", 840=>x"4d00",
---- 841=>x"6000", 842=>x"6d00", 843=>x"7900", 844=>x"4a00",
---- 845=>x"6500", 846=>x"7300", 847=>x"7600", 848=>x"4f00",
---- 849=>x"6600", 850=>x"7200", 851=>x"7600", 852=>x"5000",
---- 853=>x"6600", 854=>x"7700", 855=>x"7900", 856=>x"5300",
---- 857=>x"6000", 858=>x"7200", 859=>x"7c00", 860=>x"5800",
---- 861=>x"6300", 862=>x"7200", 863=>x"8000", 864=>x"5800",
---- 865=>x"6700", 866=>x"7200", 867=>x"8000", 868=>x"5b00",
---- 869=>x"6600", 870=>x"7300", 871=>x"8000", 872=>x"5d00",
---- 873=>x"6800", 874=>x"7700", 875=>x"7d00", 876=>x"5e00",
---- 877=>x"6700", 878=>x"7900", 879=>x"7c00", 880=>x"5e00",
---- 881=>x"6700", 882=>x"7a00", 883=>x"8400", 884=>x"6300",
---- 885=>x"6e00", 886=>x"7b00", 887=>x"7f00", 888=>x"6500",
---- 889=>x"7000", 890=>x"7e00", 891=>x"7e00", 892=>x"6400",
---- 893=>x"7300", 894=>x"8500", 895=>x"8200", 896=>x"6400",
---- 897=>x"7b00", 898=>x"8700", 899=>x"8300", 900=>x"6c00",
---- 901=>x"8100", 902=>x"8400", 903=>x"8300", 904=>x"7100",
---- 905=>x"8100", 906=>x"8300", 907=>x"8400", 908=>x"7800",
---- 909=>x"8200", 910=>x"8600", 911=>x"8800", 912=>x"7d00",
---- 913=>x"8500", 914=>x"8700", 915=>x"8900", 916=>x"8200",
---- 917=>x"8500", 918=>x"8700", 919=>x"8800", 920=>x"8200",
---- 921=>x"8800", 922=>x"8700", 923=>x"8800", 924=>x"8600",
---- 925=>x"8600", 926=>x"8600", 927=>x"8700", 928=>x"8600",
---- 929=>x"8400", 930=>x"8700", 931=>x"8900", 932=>x"8300",
---- 933=>x"8900", 934=>x"8700", 935=>x"8500", 936=>x"8600",
---- 937=>x"8600", 938=>x"8500", 939=>x"8800", 940=>x"8a00",
---- 941=>x"8600", 942=>x"8700", 943=>x"8900", 944=>x"8a00",
---- 945=>x"8700", 946=>x"8800", 947=>x"8b00", 948=>x"8800",
---- 949=>x"8900", 950=>x"8900", 951=>x"8900", 952=>x"8500",
---- 953=>x"8900", 954=>x"8c00", 955=>x"8b00", 956=>x"8600",
---- 957=>x"8800", 958=>x"8c00", 959=>x"8c00", 960=>x"8800",
---- 961=>x"8900", 962=>x"8b00", 963=>x"8b00", 964=>x"8700",
---- 965=>x"8b00", 966=>x"8a00", 967=>x"8c00", 968=>x"8600",
---- 969=>x"8c00", 970=>x"8b00", 971=>x"8c00", 972=>x"8800",
---- 973=>x"8800", 974=>x"8a00", 975=>x"8a00", 976=>x"8700",
---- 977=>x"8800", 978=>x"8900", 979=>x"8700", 980=>x"8800",
---- 981=>x"8b00", 982=>x"8800", 983=>x"8a00", 984=>x"8200",
---- 985=>x"8a00", 986=>x"8700", 987=>x"8800", 988=>x"8100",
---- 989=>x"8600", 990=>x"8700", 991=>x"8b00", 992=>x"8600",
---- 993=>x"8600", 994=>x"8700", 995=>x"8800", 996=>x"8500",
---- 997=>x"8b00", 998=>x"8a00", 999=>x"8900", 1000=>x"8600",
---- 1001=>x"8800", 1002=>x"8700", 1003=>x"8700", 1004=>x"8400",
---- 1005=>x"8600", 1006=>x"8500", 1007=>x"8700", 1008=>x"8100",
---- 1009=>x"8700", 1010=>x"8500", 1011=>x"8500", 1012=>x"8700",
---- 1013=>x"8700", 1014=>x"8b00", 1015=>x"8900", 1016=>x"8500",
---- 1017=>x"8600", 1018=>x"8800", 1019=>x"8900", 1020=>x"8200",
---- 1021=>x"8400", 1022=>x"8800", 1023=>x"8a00"),
----
---- 31 => (0=>x"8500", 1=>x"8400", 2=>x"8200", 3=>x"8500", 4=>x"8500",
---- 5=>x"8400", 6=>x"8100", 7=>x"8500", 8=>x"8500",
---- 9=>x"8400", 10=>x"8200", 11=>x"8500", 12=>x"8400",
---- 13=>x"8300", 14=>x"8300", 15=>x"8400", 16=>x"8000",
---- 17=>x"8200", 18=>x"8300", 19=>x"8400", 20=>x"8200",
---- 21=>x"8200", 22=>x"8000", 23=>x"7f00", 24=>x"8400",
---- 25=>x"8300", 26=>x"8300", 27=>x"8100", 28=>x"8500",
---- 29=>x"8100", 30=>x"8400", 31=>x"8400", 32=>x"8700",
---- 33=>x"8100", 34=>x"8600", 35=>x"8200", 36=>x"8700",
---- 37=>x"8400", 38=>x"8400", 39=>x"8300", 40=>x"8c00",
---- 41=>x"8700", 42=>x"8400", 43=>x"8300", 44=>x"8800",
---- 45=>x"8300", 46=>x"8400", 47=>x"8200", 48=>x"8300",
---- 49=>x"8500", 50=>x"8300", 51=>x"8200", 52=>x"8400",
---- 53=>x"8300", 54=>x"8400", 55=>x"8200", 56=>x"8200",
---- 57=>x"8200", 58=>x"8200", 59=>x"8400", 60=>x"8000",
---- 61=>x"8000", 62=>x"8000", 63=>x"8300", 64=>x"8100",
---- 65=>x"8100", 66=>x"8000", 67=>x"7f00", 68=>x"8100",
---- 69=>x"8300", 70=>x"8100", 71=>x"8000", 72=>x"7f00",
---- 73=>x"8100", 74=>x"8400", 75=>x"8200", 76=>x"8000",
---- 77=>x"7e00", 78=>x"8100", 79=>x"8100", 80=>x"7e00",
---- 81=>x"7f00", 82=>x"8500", 83=>x"8100", 84=>x"7d00",
---- 85=>x"8000", 86=>x"8100", 87=>x"8100", 88=>x"7900",
---- 89=>x"7900", 90=>x"7d00", 91=>x"7f00", 92=>x"7300",
---- 93=>x"7500", 94=>x"7700", 95=>x"7800", 96=>x"8400",
---- 97=>x"7900", 98=>x"7200", 99=>x"7300", 100=>x"ba00",
---- 101=>x"aa00", 102=>x"9500", 103=>x"8400", 104=>x"ba00",
---- 105=>x"c200", 106=>x"c500", 107=>x"b700", 108=>x"b800",
---- 109=>x"be00", 110=>x"bb00", 111=>x"c300", 112=>x"b400",
---- 113=>x"ba00", 114=>x"bf00", 115=>x"bd00", 116=>x"bc00",
---- 117=>x"b900", 118=>x"c000", 119=>x"bf00", 120=>x"bb00",
---- 121=>x"bd00", 122=>x"bf00", 123=>x"4000", 124=>x"4800",
---- 125=>x"b700", 126=>x"bf00", 127=>x"bc00", 128=>x"b700",
---- 129=>x"bd00", 130=>x"c000", 131=>x"bb00", 132=>x"bb00",
---- 133=>x"be00", 134=>x"bd00", 135=>x"b800", 136=>x"bd00",
---- 137=>x"bb00", 138=>x"bb00", 139=>x"bf00", 140=>x"b800",
---- 141=>x"bf00", 142=>x"be00", 143=>x"3f00", 144=>x"c000",
---- 145=>x"bf00", 146=>x"bf00", 147=>x"c400", 148=>x"c000",
---- 149=>x"c100", 150=>x"bf00", 151=>x"bd00", 152=>x"ba00",
---- 153=>x"c000", 154=>x"c000", 155=>x"be00", 156=>x"be00",
---- 157=>x"b700", 158=>x"be00", 159=>x"be00", 160=>x"b900",
---- 161=>x"be00", 162=>x"be00", 163=>x"c000", 164=>x"be00",
---- 165=>x"b800", 166=>x"b900", 167=>x"c100", 168=>x"b800",
---- 169=>x"bd00", 170=>x"bd00", 171=>x"b800", 172=>x"c200",
---- 173=>x"ac00", 174=>x"a300", 175=>x"a800", 176=>x"aa00",
---- 177=>x"9d00", 178=>x"ac00", 179=>x"c200", 180=>x"a400",
---- 181=>x"b800", 182=>x"ce00", 183=>x"d000", 184=>x"ca00",
---- 185=>x"cd00", 186=>x"cb00", 187=>x"d000", 188=>x"cf00",
---- 189=>x"d000", 190=>x"cb00", 191=>x"c600", 192=>x"ca00",
---- 193=>x"ca00", 194=>x"cb00", 195=>x"c800", 196=>x"c300",
---- 197=>x"cb00", 198=>x"d000", 199=>x"d100", 200=>x"ca00",
---- 201=>x"c500", 202=>x"cf00", 203=>x"ce00", 204=>x"c600",
---- 205=>x"c300", 206=>x"c300", 207=>x"c400", 208=>x"bb00",
---- 209=>x"c100", 210=>x"c100", 211=>x"be00", 212=>x"c100",
---- 213=>x"b800", 214=>x"c400", 215=>x"c300", 216=>x"c000",
---- 217=>x"c200", 218=>x"b800", 219=>x"b800", 220=>x"b100",
---- 221=>x"ba00", 222=>x"be00", 223=>x"c200", 224=>x"b700",
---- 225=>x"c400", 226=>x"ca00", 227=>x"c200", 228=>x"c200",
---- 229=>x"c300", 230=>x"c500", 231=>x"c800", 232=>x"bc00",
---- 233=>x"c200", 234=>x"c200", 235=>x"3b00", 236=>x"bd00",
---- 237=>x"c300", 238=>x"c600", 239=>x"c100", 240=>x"b700",
---- 241=>x"c000", 242=>x"c400", 243=>x"bf00", 244=>x"bf00",
---- 245=>x"bf00", 246=>x"c200", 247=>x"bb00", 248=>x"b900",
---- 249=>x"bf00", 250=>x"ba00", 251=>x"c100", 252=>x"ba00",
---- 253=>x"b600", 254=>x"4700", 255=>x"b900", 256=>x"c100",
---- 257=>x"ba00", 258=>x"bc00", 259=>x"b700", 260=>x"b600",
---- 261=>x"bd00", 262=>x"ba00", 263=>x"b200", 264=>x"bb00",
---- 265=>x"b400", 266=>x"aa00", 267=>x"a300", 268=>x"b100",
---- 269=>x"a100", 270=>x"a600", 271=>x"b700", 272=>x"9c00",
---- 273=>x"a400", 274=>x"be00", 275=>x"bd00", 276=>x"ae00",
---- 277=>x"b600", 278=>x"b200", 279=>x"ba00", 280=>x"b600",
---- 281=>x"b100", 282=>x"af00", 283=>x"ad00", 284=>x"ae00",
---- 285=>x"ac00", 286=>x"ad00", 287=>x"b000", 288=>x"b200",
---- 289=>x"b200", 290=>x"b200", 291=>x"ae00", 292=>x"af00",
---- 293=>x"b500", 294=>x"b300", 295=>x"ad00", 296=>x"a800",
---- 297=>x"ab00", 298=>x"b200", 299=>x"5100", 300=>x"b400",
---- 301=>x"5300", 302=>x"a500", 303=>x"b000", 304=>x"b100",
---- 305=>x"b800", 306=>x"ae00", 307=>x"a700", 308=>x"ad00",
---- 309=>x"b000", 310=>x"b600", 311=>x"ae00", 312=>x"b100",
---- 313=>x"aa00", 314=>x"a500", 315=>x"a800", 316=>x"a400",
---- 317=>x"ae00", 318=>x"a400", 319=>x"9d00", 320=>x"9c00",
---- 321=>x"9d00", 322=>x"b100", 323=>x"a800", 324=>x"a500",
---- 325=>x"9f00", 326=>x"9f00", 327=>x"ac00", 328=>x"a400",
---- 329=>x"ae00", 330=>x"a600", 331=>x"9b00", 332=>x"aa00",
---- 333=>x"a500", 334=>x"9d00", 335=>x"9000", 336=>x"8900",
---- 337=>x"9300", 338=>x"9c00", 339=>x"9e00", 340=>x"4a00",
---- 341=>x"8500", 342=>x"ae00", 343=>x"9e00", 344=>x"6100",
---- 345=>x"6a00", 346=>x"9c00", 347=>x"9c00", 348=>x"9000",
---- 349=>x"7100", 350=>x"6c00", 351=>x"6c00", 352=>x"9600",
---- 353=>x"7f00", 354=>x"8200", 355=>x"7700", 356=>x"8500",
---- 357=>x"8300", 358=>x"8300", 359=>x"7a00", 360=>x"8900",
---- 361=>x"7900", 362=>x"5900", 363=>x"4600", 364=>x"5f00",
---- 365=>x"4e00", 366=>x"5100", 367=>x"3d00", 368=>x"6400",
---- 369=>x"5500", 370=>x"4c00", 371=>x"4800", 372=>x"6d00",
---- 373=>x"6a00", 374=>x"6300", 375=>x"7b00", 376=>x"5a00",
---- 377=>x"4d00", 378=>x"4e00", 379=>x"6500", 380=>x"3b00",
---- 381=>x"3000", 382=>x"3800", 383=>x"6000", 384=>x"2a00",
---- 385=>x"2800", 386=>x"4f00", 387=>x"7600", 388=>x"2c00",
---- 389=>x"4800", 390=>x"8200", 391=>x"4e00", 392=>x"5000",
---- 393=>x"8300", 394=>x"6b00", 395=>x"4c00", 396=>x"7600",
---- 397=>x"5800", 398=>x"6200", 399=>x"7900", 400=>x"5300",
---- 401=>x"4d00", 402=>x"7000", 403=>x"5e00", 404=>x"3d00",
---- 405=>x"4000", 406=>x"6100", 407=>x"4400", 408=>x"2a00",
---- 409=>x"4200", 410=>x"6d00", 411=>x"2e00", 412=>x"2500",
---- 413=>x"4900", 414=>x"6900", 415=>x"2800", 416=>x"3c00",
---- 417=>x"5b00", 418=>x"6100", 419=>x"3b00", 420=>x"3e00",
---- 421=>x"5700", 422=>x"5200", 423=>x"4400", 424=>x"2300",
---- 425=>x"c100", 426=>x"4400", 427=>x"4e00", 428=>x"2700",
---- 429=>x"3d00", 430=>x"6100", 431=>x"7000", 432=>x"2d00",
---- 433=>x"5400", 434=>x"7f00", 435=>x"a200", 436=>x"5c00",
---- 437=>x"7c00", 438=>x"6d00", 439=>x"5100", 440=>x"9c00",
---- 441=>x"7500", 442=>x"5700", 443=>x"7b00", 444=>x"8b00",
---- 445=>x"6600", 446=>x"7e00", 447=>x"b500", 448=>x"6700",
---- 449=>x"8600", 450=>x"b700", 451=>x"b200", 452=>x"8100",
---- 453=>x"b200", 454=>x"b100", 455=>x"a600", 456=>x"4d00",
---- 457=>x"b100", 458=>x"af00", 459=>x"af00", 460=>x"b500",
---- 461=>x"ac00", 462=>x"b900", 463=>x"b400", 464=>x"a800",
---- 465=>x"b000", 466=>x"bb00", 467=>x"bc00", 468=>x"ae00",
---- 469=>x"af00", 470=>x"bc00", 471=>x"bd00", 472=>x"a700",
---- 473=>x"b300", 474=>x"bc00", 475=>x"b900", 476=>x"a200",
---- 477=>x"5400", 478=>x"ba00", 479=>x"bc00", 480=>x"9f00",
---- 481=>x"a600", 482=>x"ba00", 483=>x"c000", 484=>x"9d00",
---- 485=>x"a800", 486=>x"bc00", 487=>x"bf00", 488=>x"9800",
---- 489=>x"5900", 490=>x"bb00", 491=>x"c100", 492=>x"9800",
---- 493=>x"ac00", 494=>x"be00", 495=>x"c100", 496=>x"a000",
---- 497=>x"b600", 498=>x"bc00", 499=>x"c000", 500=>x"ac00",
---- 501=>x"ba00", 502=>x"c100", 503=>x"c800", 504=>x"b800",
---- 505=>x"c500", 506=>x"c800", 507=>x"9a00", 508=>x"c400",
---- 509=>x"c800", 510=>x"8800", 511=>x"6200", 512=>x"c400",
---- 513=>x"7400", 514=>x"5200", 515=>x"6100", 516=>x"6700",
---- 517=>x"4700", 518=>x"5100", 519=>x"4b00", 520=>x"3900",
---- 521=>x"4600", 522=>x"3a00", 523=>x"c900", 524=>x"4600",
---- 525=>x"3b00", 526=>x"3000", 527=>x"3000", 528=>x"4500",
---- 529=>x"3300", 530=>x"2900", 531=>x"2f00", 532=>x"3500",
---- 533=>x"3000", 534=>x"2c00", 535=>x"3800", 536=>x"4a00",
---- 537=>x"3a00", 538=>x"2c00", 539=>x"4000", 540=>x"7100",
---- 541=>x"5c00", 542=>x"3400", 543=>x"3400", 544=>x"8600",
---- 545=>x"7600", 546=>x"5100", 547=>x"4200", 548=>x"8d00",
---- 549=>x"8a00", 550=>x"7a00", 551=>x"6b00", 552=>x"9000",
---- 553=>x"9000", 554=>x"8d00", 555=>x"7b00", 556=>x"9000",
---- 557=>x"9000", 558=>x"9200", 559=>x"8d00", 560=>x"9500",
---- 561=>x"9100", 562=>x"8d00", 563=>x"9000", 564=>x"9700",
---- 565=>x"9700", 566=>x"9700", 567=>x"9400", 568=>x"9d00",
---- 569=>x"a000", 570=>x"a200", 571=>x"a000", 572=>x"a300",
---- 573=>x"a700", 574=>x"a400", 575=>x"a300", 576=>x"a100",
---- 577=>x"aa00", 578=>x"a400", 579=>x"a400", 580=>x"a100",
---- 581=>x"a600", 582=>x"aa00", 583=>x"a700", 584=>x"a100",
---- 585=>x"a400", 586=>x"ad00", 587=>x"ab00", 588=>x"9f00",
---- 589=>x"a600", 590=>x"a800", 591=>x"ab00", 592=>x"9d00",
---- 593=>x"a200", 594=>x"a900", 595=>x"ae00", 596=>x"9900",
---- 597=>x"a000", 598=>x"a800", 599=>x"ab00", 600=>x"6700",
---- 601=>x"9c00", 602=>x"9e00", 603=>x"a300", 604=>x"9900",
---- 605=>x"9800", 606=>x"9b00", 607=>x"a100", 608=>x"9800",
---- 609=>x"9b00", 610=>x"9d00", 611=>x"a000", 612=>x"9700",
---- 613=>x"9b00", 614=>x"9e00", 615=>x"a000", 616=>x"9800",
---- 617=>x"9c00", 618=>x"9b00", 619=>x"9f00", 620=>x"6d00",
---- 621=>x"9800", 622=>x"9800", 623=>x"9d00", 624=>x"9200",
---- 625=>x"9600", 626=>x"9600", 627=>x"9800", 628=>x"9300",
---- 629=>x"9400", 630=>x"9600", 631=>x"9700", 632=>x"9200",
---- 633=>x"9100", 634=>x"9a00", 635=>x"9800", 636=>x"8f00",
---- 637=>x"8f00", 638=>x"6c00", 639=>x"9600", 640=>x"8f00",
---- 641=>x"9000", 642=>x"9200", 643=>x"9600", 644=>x"8f00",
---- 645=>x"8f00", 646=>x"9600", 647=>x"9600", 648=>x"6e00",
---- 649=>x"9100", 650=>x"9300", 651=>x"9700", 652=>x"9100",
---- 653=>x"9100", 654=>x"9100", 655=>x"9400", 656=>x"8d00",
---- 657=>x"9300", 658=>x"9100", 659=>x"9400", 660=>x"8a00",
---- 661=>x"8f00", 662=>x"9000", 663=>x"9000", 664=>x"8900",
---- 665=>x"8e00", 666=>x"9100", 667=>x"8f00", 668=>x"8d00",
---- 669=>x"8d00", 670=>x"8b00", 671=>x"8d00", 672=>x"8d00",
---- 673=>x"8d00", 674=>x"8d00", 675=>x"8a00", 676=>x"8c00",
---- 677=>x"8b00", 678=>x"8d00", 679=>x"8b00", 680=>x"8b00",
---- 681=>x"8e00", 682=>x"8c00", 683=>x"8900", 684=>x"7500",
---- 685=>x"8f00", 686=>x"8b00", 687=>x"8e00", 688=>x"8b00",
---- 689=>x"8a00", 690=>x"8d00", 691=>x"8a00", 692=>x"8600",
---- 693=>x"8a00", 694=>x"8d00", 695=>x"8d00", 696=>x"8600",
---- 697=>x"8500", 698=>x"8b00", 699=>x"9100", 700=>x"8700",
---- 701=>x"8a00", 702=>x"8b00", 703=>x"8d00", 704=>x"8700",
---- 705=>x"8b00", 706=>x"8800", 707=>x"8b00", 708=>x"8400",
---- 709=>x"8800", 710=>x"8800", 711=>x"8700", 712=>x"8100",
---- 713=>x"8200", 714=>x"8600", 715=>x"8800", 716=>x"7f00",
---- 717=>x"8200", 718=>x"7e00", 719=>x"8500", 720=>x"7d00",
---- 721=>x"8100", 722=>x"8000", 723=>x"8200", 724=>x"7c00",
---- 725=>x"8200", 726=>x"8400", 727=>x"8400", 728=>x"7800",
---- 729=>x"7f00", 730=>x"8300", 731=>x"8100", 732=>x"7800",
---- 733=>x"7c00", 734=>x"8100", 735=>x"8100", 736=>x"7a00",
---- 737=>x"7e00", 738=>x"8000", 739=>x"7f00", 740=>x"7700",
---- 741=>x"7e00", 742=>x"7e00", 743=>x"7f00", 744=>x"7100",
---- 745=>x"7c00", 746=>x"7f00", 747=>x"7f00", 748=>x"6f00",
---- 749=>x"7600", 750=>x"7c00", 751=>x"8300", 752=>x"6800",
---- 753=>x"7000", 754=>x"7600", 755=>x"7f00", 756=>x"5c00",
---- 757=>x"9600", 758=>x"7500", 759=>x"7800", 760=>x"5200",
---- 761=>x"6000", 762=>x"6f00", 763=>x"7600", 764=>x"4a00",
---- 765=>x"5400", 766=>x"6000", 767=>x"6800", 768=>x"3b00",
---- 769=>x"4000", 770=>x"4300", 771=>x"4500", 772=>x"4500",
---- 773=>x"4600", 774=>x"4800", 775=>x"4d00", 776=>x"6c00",
---- 777=>x"6d00", 778=>x"7500", 779=>x"7c00", 780=>x"7700",
---- 781=>x"7b00", 782=>x"8200", 783=>x"8300", 784=>x"8000",
---- 785=>x"8200", 786=>x"8100", 787=>x"7e00", 788=>x"7f00",
---- 789=>x"8000", 790=>x"7e00", 791=>x"7c00", 792=>x"7c00",
---- 793=>x"7d00", 794=>x"7e00", 795=>x"7c00", 796=>x"7500",
---- 797=>x"7c00", 798=>x"7e00", 799=>x"7d00", 800=>x"7a00",
---- 801=>x"7c00", 802=>x"7a00", 803=>x"7b00", 804=>x"7200",
---- 805=>x"7a00", 806=>x"7b00", 807=>x"7c00", 808=>x"7400",
---- 809=>x"7700", 810=>x"7b00", 811=>x"7e00", 812=>x"8800",
---- 813=>x"7600", 814=>x"7b00", 815=>x"8100", 816=>x"7800",
---- 817=>x"7d00", 818=>x"7e00", 819=>x"7e00", 820=>x"7900",
---- 821=>x"8300", 822=>x"7e00", 823=>x"7200", 824=>x"7700",
---- 825=>x"7c00", 826=>x"7100", 827=>x"6f00", 828=>x"7300",
---- 829=>x"7000", 830=>x"7700", 831=>x"8100", 832=>x"6c00",
---- 833=>x"7900", 834=>x"8800", 835=>x"8300", 836=>x"7a00",
---- 837=>x"8500", 838=>x"8a00", 839=>x"8200", 840=>x"7c00",
---- 841=>x"8300", 842=>x"8700", 843=>x"8300", 844=>x"7f00",
---- 845=>x"8500", 846=>x"8500", 847=>x"8300", 848=>x"8000",
---- 849=>x"8300", 850=>x"8000", 851=>x"8000", 852=>x"8000",
---- 853=>x"8200", 854=>x"7e00", 855=>x"7d00", 856=>x"8500",
---- 857=>x"8400", 858=>x"8100", 859=>x"8100", 860=>x"8300",
---- 861=>x"8000", 862=>x"8000", 863=>x"8200", 864=>x"8400",
---- 865=>x"8300", 866=>x"8400", 867=>x"8600", 868=>x"8400",
---- 869=>x"8500", 870=>x"8800", 871=>x"8600", 872=>x"8200",
---- 873=>x"8100", 874=>x"8700", 875=>x"8a00", 876=>x"7f00",
---- 877=>x"8400", 878=>x"8500", 879=>x"8800", 880=>x"8200",
---- 881=>x"8500", 882=>x"8300", 883=>x"8500", 884=>x"8400",
---- 885=>x"8500", 886=>x"8300", 887=>x"8700", 888=>x"8500",
---- 889=>x"8600", 890=>x"8600", 891=>x"8400", 892=>x"8400",
---- 893=>x"8700", 894=>x"8600", 895=>x"8700", 896=>x"8600",
---- 897=>x"8500", 898=>x"8a00", 899=>x"8a00", 900=>x"7800",
---- 901=>x"7500", 902=>x"8a00", 903=>x"8a00", 904=>x"8a00",
---- 905=>x"8c00", 906=>x"8900", 907=>x"8c00", 908=>x"8c00",
---- 909=>x"8d00", 910=>x"8c00", 911=>x"8b00", 912=>x"8900",
---- 913=>x"8e00", 914=>x"8e00", 915=>x"8a00", 916=>x"8c00",
---- 917=>x"8800", 918=>x"8c00", 919=>x"8e00", 920=>x"8b00",
---- 921=>x"8a00", 922=>x"8a00", 923=>x"8b00", 924=>x"8a00",
---- 925=>x"8c00", 926=>x"8b00", 927=>x"8e00", 928=>x"8b00",
---- 929=>x"8d00", 930=>x"8f00", 931=>x"8f00", 932=>x"8800",
---- 933=>x"8d00", 934=>x"8d00", 935=>x"8e00", 936=>x"8800",
---- 937=>x"8900", 938=>x"8d00", 939=>x"8b00", 940=>x"8a00",
---- 941=>x"8c00", 942=>x"8d00", 943=>x"8c00", 944=>x"8b00",
---- 945=>x"8b00", 946=>x"8b00", 947=>x"8b00", 948=>x"8900",
---- 949=>x"8900", 950=>x"8b00", 951=>x"8b00", 952=>x"8b00",
---- 953=>x"8b00", 954=>x"8b00", 955=>x"8b00", 956=>x"8a00",
---- 957=>x"8a00", 958=>x"8900", 959=>x"8c00", 960=>x"8b00",
---- 961=>x"8a00", 962=>x"8a00", 963=>x"8c00", 964=>x"8c00",
---- 965=>x"8b00", 966=>x"8900", 967=>x"8a00", 968=>x"8b00",
---- 969=>x"8900", 970=>x"8c00", 971=>x"7500", 972=>x"8900",
---- 973=>x"8c00", 974=>x"8f00", 975=>x"8b00", 976=>x"8900",
---- 977=>x"8e00", 978=>x"8c00", 979=>x"8d00", 980=>x"8a00",
---- 981=>x"8b00", 982=>x"8c00", 983=>x"8a00", 984=>x"8b00",
---- 985=>x"8c00", 986=>x"8b00", 987=>x"8900", 988=>x"8a00",
---- 989=>x"8800", 990=>x"8700", 991=>x"8800", 992=>x"8700",
---- 993=>x"8600", 994=>x"8800", 995=>x"8c00", 996=>x"8700",
---- 997=>x"8900", 998=>x"8800", 999=>x"8b00", 1000=>x"8600",
---- 1001=>x"8b00", 1002=>x"8900", 1003=>x"8a00", 1004=>x"8a00",
---- 1005=>x"8a00", 1006=>x"8900", 1007=>x"8900", 1008=>x"8a00",
---- 1009=>x"8900", 1010=>x"8700", 1011=>x"8700", 1012=>x"8800",
---- 1013=>x"8500", 1014=>x"8500", 1015=>x"8700", 1016=>x"8a00",
---- 1017=>x"8900", 1018=>x"8400", 1019=>x"8600", 1020=>x"8b00",
---- 1021=>x"8800", 1022=>x"8500", 1023=>x"8500"),
----
---- 32 => (0=>x"8c00", 1=>x"8800", 2=>x"8200", 3=>x"8000", 4=>x"8c00",
---- 5=>x"8600", 6=>x"8200", 7=>x"8000", 8=>x"8a00",
---- 9=>x"8800", 10=>x"8300", 11=>x"7f00", 12=>x"8300",
---- 13=>x"8600", 14=>x"8400", 15=>x"8000", 16=>x"8300",
---- 17=>x"8500", 18=>x"8200", 19=>x"8200", 20=>x"8100",
---- 21=>x"8300", 22=>x"8200", 23=>x"8400", 24=>x"8100",
---- 25=>x"8200", 26=>x"8200", 27=>x"8300", 28=>x"8100",
---- 29=>x"8300", 30=>x"8200", 31=>x"8200", 32=>x"8200",
---- 33=>x"8100", 34=>x"8300", 35=>x"8200", 36=>x"8300",
---- 37=>x"8300", 38=>x"8300", 39=>x"8400", 40=>x"8400",
---- 41=>x"8300", 42=>x"8200", 43=>x"8000", 44=>x"8200",
---- 45=>x"8200", 46=>x"8200", 47=>x"8100", 48=>x"8100",
---- 49=>x"8100", 50=>x"8300", 51=>x"8300", 52=>x"8300",
---- 53=>x"8400", 54=>x"8300", 55=>x"8400", 56=>x"8200",
---- 57=>x"8400", 58=>x"8500", 59=>x"8400", 60=>x"8500",
---- 61=>x"8100", 62=>x"8400", 63=>x"8200", 64=>x"8500",
---- 65=>x"8300", 66=>x"8300", 67=>x"8100", 68=>x"8300",
---- 69=>x"8500", 70=>x"8300", 71=>x"8100", 72=>x"8300",
---- 73=>x"8400", 74=>x"8400", 75=>x"8000", 76=>x"8600",
---- 77=>x"8200", 78=>x"8200", 79=>x"8200", 80=>x"8300",
---- 81=>x"8200", 82=>x"7f00", 83=>x"7e00", 84=>x"8000",
---- 85=>x"8400", 86=>x"8000", 87=>x"8000", 88=>x"7c00",
---- 89=>x"7d00", 90=>x"7c00", 91=>x"7e00", 92=>x"7800",
---- 93=>x"7d00", 94=>x"7b00", 95=>x"7c00", 96=>x"7600",
---- 97=>x"7800", 98=>x"7a00", 99=>x"7c00", 100=>x"7400",
---- 101=>x"7100", 102=>x"7100", 103=>x"7900", 104=>x"a700",
---- 105=>x"8f00", 106=>x"7700", 107=>x"6f00", 108=>x"c400",
---- 109=>x"c000", 110=>x"b100", 111=>x"8900", 112=>x"c200",
---- 113=>x"c600", 114=>x"c800", 115=>x"c200", 116=>x"c100",
---- 117=>x"c400", 118=>x"c200", 119=>x"c500", 120=>x"c100",
---- 121=>x"c400", 122=>x"c000", 123=>x"c100", 124=>x"bc00",
---- 125=>x"c200", 126=>x"c200", 127=>x"c100", 128=>x"bd00",
---- 129=>x"bb00", 130=>x"bf00", 131=>x"c100", 132=>x"b800",
---- 133=>x"bf00", 134=>x"c200", 135=>x"c100", 136=>x"bd00",
---- 137=>x"bd00", 138=>x"c000", 139=>x"c300", 140=>x"c100",
---- 141=>x"be00", 142=>x"bd00", 143=>x"c300", 144=>x"bf00",
---- 145=>x"bf00", 146=>x"c400", 147=>x"c300", 148=>x"c100",
---- 149=>x"3d00", 150=>x"c100", 151=>x"c700", 152=>x"be00",
---- 153=>x"c100", 154=>x"c400", 155=>x"c500", 156=>x"c400",
---- 157=>x"b900", 158=>x"c300", 159=>x"c500", 160=>x"c000",
---- 161=>x"c000", 162=>x"c400", 163=>x"bc00", 164=>x"c100",
---- 165=>x"bc00", 166=>x"b000", 167=>x"b100", 168=>x"ab00",
---- 169=>x"ab00", 170=>x"b100", 171=>x"be00", 172=>x"b400",
---- 173=>x"c500", 174=>x"cf00", 175=>x"d700", 176=>x"d100",
---- 177=>x"d500", 178=>x"d500", 179=>x"d500", 180=>x"d200",
---- 181=>x"d600", 182=>x"ce00", 183=>x"cb00", 184=>x"ca00",
---- 185=>x"cb00", 186=>x"c900", 187=>x"ce00", 188=>x"c800",
---- 189=>x"c900", 190=>x"cf00", 191=>x"d700", 192=>x"c900",
---- 193=>x"d200", 194=>x"ca00", 195=>x"ce00", 196=>x"cb00",
---- 197=>x"c600", 198=>x"ca00", 199=>x"c700", 200=>x"ca00",
---- 201=>x"c300", 202=>x"3a00", 203=>x"ca00", 204=>x"c500",
---- 205=>x"3a00", 206=>x"c600", 207=>x"c900", 208=>x"c300",
---- 209=>x"c600", 210=>x"3b00", 211=>x"c100", 212=>x"b700",
---- 213=>x"bc00", 214=>x"bc00", 215=>x"c400", 216=>x"b700",
---- 217=>x"c100", 218=>x"c900", 219=>x"3800", 220=>x"c700",
---- 221=>x"c300", 222=>x"c400", 223=>x"ca00", 224=>x"c400",
---- 225=>x"c500", 226=>x"c000", 227=>x"c200", 228=>x"c200",
---- 229=>x"c500", 230=>x"ca00", 231=>x"c100", 232=>x"c900",
---- 233=>x"c200", 234=>x"c500", 235=>x"c700", 236=>x"c400",
---- 237=>x"c400", 238=>x"bd00", 239=>x"c800", 240=>x"c300",
---- 241=>x"c400", 242=>x"c400", 243=>x"4200", 244=>x"bf00",
---- 245=>x"c500", 246=>x"c200", 247=>x"c300", 248=>x"ba00",
---- 249=>x"c000", 250=>x"c600", 251=>x"c200", 252=>x"c200",
---- 253=>x"bc00", 254=>x"b600", 255=>x"b300", 256=>x"b600",
---- 257=>x"b300", 258=>x"ad00", 259=>x"bd00", 260=>x"a400",
---- 261=>x"ac00", 262=>x"c000", 263=>x"c000", 264=>x"b100",
---- 265=>x"c000", 266=>x"bf00", 267=>x"bc00", 268=>x"b500",
---- 269=>x"b300", 270=>x"be00", 271=>x"bf00", 272=>x"b700",
---- 273=>x"b100", 274=>x"b500", 275=>x"bf00", 276=>x"bb00",
---- 277=>x"b500", 278=>x"b600", 279=>x"b500", 280=>x"b900",
---- 281=>x"bb00", 282=>x"b200", 283=>x"b400", 284=>x"b000",
---- 285=>x"b500", 286=>x"b500", 287=>x"ac00", 288=>x"af00",
---- 289=>x"b000", 290=>x"ae00", 291=>x"b400", 292=>x"ad00",
---- 293=>x"b200", 294=>x"a900", 295=>x"ad00", 296=>x"b000",
---- 297=>x"ad00", 298=>x"a900", 299=>x"5800", 300=>x"b200",
---- 301=>x"ad00", 302=>x"ae00", 303=>x"aa00", 304=>x"b200",
---- 305=>x"b200", 306=>x"ae00", 307=>x"aa00", 308=>x"a400",
---- 309=>x"a100", 310=>x"a700", 311=>x"b100", 312=>x"a500",
---- 313=>x"9f00", 314=>x"9d00", 315=>x"a500", 316=>x"a900",
---- 317=>x"a700", 318=>x"a600", 319=>x"a500", 320=>x"a000",
---- 321=>x"a800", 322=>x"ac00", 323=>x"aa00", 324=>x"ad00",
---- 325=>x"9b00", 326=>x"9800", 327=>x"9a00", 328=>x"9e00",
---- 329=>x"8800", 330=>x"9800", 331=>x"ab00", 332=>x"9800",
---- 333=>x"a000", 334=>x"5e00", 335=>x"a600", 336=>x"a700",
---- 337=>x"a700", 338=>x"a300", 339=>x"a200", 340=>x"a100",
---- 341=>x"a200", 342=>x"9e00", 343=>x"9d00", 344=>x"a200",
---- 345=>x"a700", 346=>x"a600", 347=>x"a200", 348=>x"7b00",
---- 349=>x"8100", 350=>x"8400", 351=>x"a400", 352=>x"7900",
---- 353=>x"7400", 354=>x"6500", 355=>x"6000", 356=>x"7a00",
---- 357=>x"6e00", 358=>x"5900", 359=>x"4900", 360=>x"4600",
---- 361=>x"3f00", 362=>x"3f00", 363=>x"6d00", 364=>x"3400",
---- 365=>x"4f00", 366=>x"7300", 367=>x"5c00", 368=>x"6100",
---- 369=>x"6500", 370=>x"4d00", 371=>x"4900", 372=>x"6a00",
---- 373=>x"5800", 374=>x"7100", 375=>x"4700", 376=>x"5500",
---- 377=>x"7e00", 378=>x"5c00", 379=>x"4100", 380=>x"5f00",
---- 381=>x"4f00", 382=>x"5500", 383=>x"6200", 384=>x"3f00",
---- 385=>x"5100", 386=>x"7100", 387=>x"4200", 388=>x"4500",
---- 389=>x"6200", 390=>x"4a00", 391=>x"2200", 392=>x"6100",
---- 393=>x"4700", 394=>x"1f00", 395=>x"3600", 396=>x"5d00",
---- 397=>x"2000", 398=>x"3700", 399=>x"6b00", 400=>x"2f00",
---- 401=>x"3100", 402=>x"7d00", 403=>x"a900", 404=>x"2000",
---- 405=>x"6a00", 406=>x"9500", 407=>x"2800", 408=>x"2200",
---- 409=>x"7e00", 410=>x"6800", 411=>x"3700", 412=>x"3f00",
---- 413=>x"8100", 414=>x"6b00", 415=>x"8800", 416=>x"5b00",
---- 417=>x"7500", 418=>x"7200", 419=>x"8e00", 420=>x"4f00",
---- 421=>x"6800", 422=>x"5700", 423=>x"8500", 424=>x"5700",
---- 425=>x"5000", 426=>x"5100", 427=>x"7a00", 428=>x"5b00",
---- 429=>x"4c00", 430=>x"5e00", 431=>x"8600", 432=>x"ae00",
---- 433=>x"6400", 434=>x"8800", 435=>x"9c00", 436=>x"7900",
---- 437=>x"9900", 438=>x"8c00", 439=>x"9e00", 440=>x"af00",
---- 441=>x"a400", 442=>x"7b00", 443=>x"9900", 444=>x"a800",
---- 445=>x"a100", 446=>x"8300", 447=>x"8700", 448=>x"a200",
---- 449=>x"a600", 450=>x"8e00", 451=>x"8700", 452=>x"a500",
---- 453=>x"a800", 454=>x"9200", 455=>x"8f00", 456=>x"a500",
---- 457=>x"ac00", 458=>x"9500", 459=>x"6d00", 460=>x"af00",
---- 461=>x"b200", 462=>x"9e00", 463=>x"9200", 464=>x"b500",
---- 465=>x"b400", 466=>x"9c00", 467=>x"6f00", 468=>x"ba00",
---- 469=>x"b700", 470=>x"9700", 471=>x"8300", 472=>x"bb00",
---- 473=>x"b900", 474=>x"5900", 475=>x"7f00", 476=>x"ba00",
---- 477=>x"ba00", 478=>x"b500", 479=>x"9500", 480=>x"b700",
---- 481=>x"4500", 482=>x"b600", 483=>x"aa00", 484=>x"ba00",
---- 485=>x"bd00", 486=>x"b600", 487=>x"b300", 488=>x"c000",
---- 489=>x"bf00", 490=>x"be00", 491=>x"bb00", 492=>x"c200",
---- 493=>x"c500", 494=>x"b800", 495=>x"8000", 496=>x"c600",
---- 497=>x"b300", 498=>x"8200", 499=>x"7400", 500=>x"a800",
---- 501=>x"7a00", 502=>x"7f00", 503=>x"9100", 504=>x"7000",
---- 505=>x"7d00", 506=>x"8300", 507=>x"8c00", 508=>x"7100",
---- 509=>x"7300", 510=>x"7100", 511=>x"7800", 512=>x"5f00",
---- 513=>x"6000", 514=>x"5100", 515=>x"4b00", 516=>x"3a00",
---- 517=>x"3e00", 518=>x"3b00", 519=>x"3600", 520=>x"3300",
---- 521=>x"3300", 522=>x"3500", 523=>x"3200", 524=>x"2f00",
---- 525=>x"3100", 526=>x"3200", 527=>x"3000", 528=>x"4100",
---- 529=>x"3d00", 530=>x"3300", 531=>x"3b00", 532=>x"5e00",
---- 533=>x"5500", 534=>x"3f00", 535=>x"5d00", 536=>x"6000",
---- 537=>x"7500", 538=>x"4500", 539=>x"4f00", 540=>x"5d00",
---- 541=>x"7800", 542=>x"6c00", 543=>x"4300", 544=>x"6100",
---- 545=>x"7100", 546=>x"8000", 547=>x"7a00", 548=>x"5f00",
---- 549=>x"5f00", 550=>x"7c00", 551=>x"8700", 552=>x"7b00",
---- 553=>x"7e00", 554=>x"6d00", 555=>x"7100", 556=>x"9000",
---- 557=>x"8800", 558=>x"8d00", 559=>x"7b00", 560=>x"9700",
---- 561=>x"8e00", 562=>x"8500", 563=>x"8a00", 564=>x"6c00",
---- 565=>x"9100", 566=>x"9000", 567=>x"9200", 568=>x"9c00",
---- 569=>x"9600", 570=>x"9500", 571=>x"9800", 572=>x"aa00",
---- 573=>x"aa00", 574=>x"a300", 575=>x"a400", 576=>x"ac00",
---- 577=>x"b000", 578=>x"ab00", 579=>x"a600", 580=>x"ac00",
---- 581=>x"af00", 582=>x"ab00", 583=>x"b000", 584=>x"ac00",
---- 585=>x"b400", 586=>x"af00", 587=>x"ab00", 588=>x"ad00",
---- 589=>x"b100", 590=>x"b300", 591=>x"b000", 592=>x"ae00",
---- 593=>x"b300", 594=>x"b300", 595=>x"b300", 596=>x"ae00",
---- 597=>x"b200", 598=>x"b200", 599=>x"b200", 600=>x"a700",
---- 601=>x"ad00", 602=>x"b200", 603=>x"b300", 604=>x"a600",
---- 605=>x"a800", 606=>x"ac00", 607=>x"af00", 608=>x"a700",
---- 609=>x"a900", 610=>x"ad00", 611=>x"af00", 612=>x"9f00",
---- 613=>x"a300", 614=>x"a900", 615=>x"ae00", 616=>x"a200",
---- 617=>x"9f00", 618=>x"a100", 619=>x"a900", 620=>x"a100",
---- 621=>x"9f00", 622=>x"9d00", 623=>x"a100", 624=>x"9a00",
---- 625=>x"9d00", 626=>x"9c00", 627=>x"9b00", 628=>x"6900",
---- 629=>x"9800", 630=>x"9a00", 631=>x"9c00", 632=>x"9700",
---- 633=>x"9800", 634=>x"9900", 635=>x"9c00", 636=>x"9700",
---- 637=>x"9700", 638=>x"9e00", 639=>x"9c00", 640=>x"9700",
---- 641=>x"9600", 642=>x"9600", 643=>x"9800", 644=>x"9600",
---- 645=>x"9800", 646=>x"9900", 647=>x"9700", 648=>x"9700",
---- 649=>x"9700", 650=>x"9900", 651=>x"9500", 652=>x"9700",
---- 653=>x"9300", 654=>x"9600", 655=>x"9800", 656=>x"9400",
---- 657=>x"9000", 658=>x"9500", 659=>x"9300", 660=>x"9000",
---- 661=>x"9200", 662=>x"9700", 663=>x"9400", 664=>x"9000",
---- 665=>x"9000", 666=>x"9000", 667=>x"9400", 668=>x"8f00",
---- 669=>x"9000", 670=>x"9400", 671=>x"9800", 672=>x"8a00",
---- 673=>x"8c00", 674=>x"9000", 675=>x"9300", 676=>x"8e00",
---- 677=>x"8d00", 678=>x"8e00", 679=>x"8e00", 680=>x"8f00",
---- 681=>x"8c00", 682=>x"8d00", 683=>x"8e00", 684=>x"8c00",
---- 685=>x"8800", 686=>x"8a00", 687=>x"8b00", 688=>x"8a00",
---- 689=>x"8700", 690=>x"8900", 691=>x"8c00", 692=>x"8c00",
---- 693=>x"8700", 694=>x"8800", 695=>x"8d00", 696=>x"8e00",
---- 697=>x"8c00", 698=>x"8c00", 699=>x"9200", 700=>x"8f00",
---- 701=>x"9000", 702=>x"8f00", 703=>x"9200", 704=>x"9000",
---- 705=>x"9400", 706=>x"9100", 707=>x"9100", 708=>x"9100",
---- 709=>x"9300", 710=>x"9200", 711=>x"9100", 712=>x"8f00",
---- 713=>x"9300", 714=>x"9100", 715=>x"8f00", 716=>x"8a00",
---- 717=>x"8e00", 718=>x"8f00", 719=>x"9300", 720=>x"8700",
---- 721=>x"8c00", 722=>x"8d00", 723=>x"9000", 724=>x"8800",
---- 725=>x"8900", 726=>x"8a00", 727=>x"8b00", 728=>x"8600",
---- 729=>x"8900", 730=>x"8a00", 731=>x"8c00", 732=>x"8300",
---- 733=>x"7900", 734=>x"8a00", 735=>x"8900", 736=>x"8400",
---- 737=>x"8500", 738=>x"8700", 739=>x"8a00", 740=>x"8600",
---- 741=>x"8400", 742=>x"8800", 743=>x"7600", 744=>x"8300",
---- 745=>x"8700", 746=>x"8800", 747=>x"8900", 748=>x"8400",
---- 749=>x"8400", 750=>x"8400", 751=>x"8900", 752=>x"8100",
---- 753=>x"8200", 754=>x"8400", 755=>x"8600", 756=>x"7d00",
---- 757=>x"8100", 758=>x"8400", 759=>x"8700", 760=>x"7900",
---- 761=>x"7c00", 762=>x"7f00", 763=>x"8400", 764=>x"6900",
---- 765=>x"7000", 766=>x"7b00", 767=>x"7c00", 768=>x"4600",
---- 769=>x"4f00", 770=>x"5c00", 771=>x"6200", 772=>x"5900",
---- 773=>x"5d00", 774=>x"6200", 775=>x"6400", 776=>x"7f00",
---- 777=>x"8400", 778=>x"8900", 779=>x"8b00", 780=>x"8300",
---- 781=>x"8600", 782=>x"8c00", 783=>x"8d00", 784=>x"7d00",
---- 785=>x"8000", 786=>x"8400", 787=>x"8500", 788=>x"7e00",
---- 789=>x"8000", 790=>x"8400", 791=>x"8400", 792=>x"7c00",
---- 793=>x"7e00", 794=>x"8100", 795=>x"8300", 796=>x"7d00",
---- 797=>x"8100", 798=>x"7d00", 799=>x"8200", 800=>x"7c00",
---- 801=>x"7f00", 802=>x"8000", 803=>x"8200", 804=>x"7e00",
---- 805=>x"8100", 806=>x"8300", 807=>x"7e00", 808=>x"7c00",
---- 809=>x"8200", 810=>x"7b00", 811=>x"7c00", 812=>x"7f00",
---- 813=>x"7b00", 814=>x"7c00", 815=>x"8400", 816=>x"7a00",
---- 817=>x"7800", 818=>x"8400", 819=>x"8800", 820=>x"7200",
---- 821=>x"8000", 822=>x"8800", 823=>x"8b00", 824=>x"7c00",
---- 825=>x"8700", 826=>x"8500", 827=>x"8b00", 828=>x"8400",
---- 829=>x"8600", 830=>x"8800", 831=>x"8b00", 832=>x"7f00",
---- 833=>x"8800", 834=>x"8a00", 835=>x"8b00", 836=>x"8000",
---- 837=>x"8600", 838=>x"8900", 839=>x"8800", 840=>x"8500",
---- 841=>x"8300", 842=>x"8600", 843=>x"8900", 844=>x"8500",
---- 845=>x"8500", 846=>x"8600", 847=>x"8700", 848=>x"8800",
---- 849=>x"8800", 850=>x"8300", 851=>x"8300", 852=>x"8600",
---- 853=>x"8600", 854=>x"8600", 855=>x"8700", 856=>x"8400",
---- 857=>x"8900", 858=>x"8a00", 859=>x"8a00", 860=>x"8800",
---- 861=>x"8900", 862=>x"8800", 863=>x"8a00", 864=>x"8800",
---- 865=>x"8900", 866=>x"8700", 867=>x"8900", 868=>x"8600",
---- 869=>x"8a00", 870=>x"8a00", 871=>x"8800", 872=>x"8900",
---- 873=>x"8800", 874=>x"8c00", 875=>x"8900", 876=>x"8900",
---- 877=>x"8b00", 878=>x"8a00", 879=>x"8a00", 880=>x"8a00",
---- 881=>x"8a00", 882=>x"8c00", 883=>x"8c00", 884=>x"8a00",
---- 885=>x"8b00", 886=>x"9000", 887=>x"8f00", 888=>x"8900",
---- 889=>x"8c00", 890=>x"8e00", 891=>x"8d00", 892=>x"8b00",
---- 893=>x"8900", 894=>x"8d00", 895=>x"8b00", 896=>x"8b00",
---- 897=>x"8c00", 898=>x"8900", 899=>x"8b00", 900=>x"8a00",
---- 901=>x"8c00", 902=>x"8c00", 903=>x"8c00", 904=>x"8a00",
---- 905=>x"8a00", 906=>x"8d00", 907=>x"8f00", 908=>x"8c00",
---- 909=>x"9000", 910=>x"8d00", 911=>x"8a00", 912=>x"8d00",
---- 913=>x"9200", 914=>x"9000", 915=>x"8b00", 916=>x"8c00",
---- 917=>x"8f00", 918=>x"9500", 919=>x"8f00", 920=>x"8d00",
---- 921=>x"9000", 922=>x"8f00", 923=>x"9000", 924=>x"8f00",
---- 925=>x"8f00", 926=>x"8f00", 927=>x"9100", 928=>x"8e00",
---- 929=>x"9200", 930=>x"8f00", 931=>x"8b00", 932=>x"8e00",
---- 933=>x"9200", 934=>x"9000", 935=>x"8a00", 936=>x"8d00",
---- 937=>x"9000", 938=>x"8e00", 939=>x"8b00", 940=>x"8e00",
---- 941=>x"8c00", 942=>x"8d00", 943=>x"8e00", 944=>x"8900",
---- 945=>x"8c00", 946=>x"8d00", 947=>x"8e00", 948=>x"8a00",
---- 949=>x"8d00", 950=>x"8b00", 951=>x"9000", 952=>x"8b00",
---- 953=>x"8d00", 954=>x"8a00", 955=>x"9000", 956=>x"8b00",
---- 957=>x"8c00", 958=>x"8a00", 959=>x"9100", 960=>x"8c00",
---- 961=>x"8c00", 962=>x"8c00", 963=>x"8e00", 964=>x"8c00",
---- 965=>x"8900", 966=>x"8900", 967=>x"8a00", 968=>x"8c00",
---- 969=>x"8b00", 970=>x"8c00", 971=>x"8c00", 972=>x"8b00",
---- 973=>x"8c00", 974=>x"8d00", 975=>x"8e00", 976=>x"8b00",
---- 977=>x"8b00", 978=>x"8e00", 979=>x"8f00", 980=>x"8800",
---- 981=>x"8b00", 982=>x"9000", 983=>x"8e00", 984=>x"8a00",
---- 985=>x"8c00", 986=>x"8c00", 987=>x"8a00", 988=>x"8c00",
---- 989=>x"8d00", 990=>x"8e00", 991=>x"8d00", 992=>x"8e00",
---- 993=>x"8d00", 994=>x"8c00", 995=>x"8d00", 996=>x"8d00",
---- 997=>x"8c00", 998=>x"8b00", 999=>x"8c00", 1000=>x"8b00",
---- 1001=>x"8900", 1002=>x"8800", 1003=>x"8c00", 1004=>x"8800",
---- 1005=>x"8a00", 1006=>x"8c00", 1007=>x"8c00", 1008=>x"8b00",
---- 1009=>x"7200", 1010=>x"8b00", 1011=>x"8a00", 1012=>x"8d00",
---- 1013=>x"8d00", 1014=>x"8a00", 1015=>x"8d00", 1016=>x"8800",
---- 1017=>x"8800", 1018=>x"8b00", 1019=>x"8c00", 1020=>x"8700",
---- 1021=>x"8600", 1022=>x"8900", 1023=>x"8b00"),
----
---- 33 => (0=>x"8400", 1=>x"8200", 2=>x"8500", 3=>x"8300", 4=>x"8500",
---- 5=>x"8200", 6=>x"8500", 7=>x"8300", 8=>x"8300",
---- 9=>x"8400", 10=>x"8300", 11=>x"8200", 12=>x"8000",
---- 13=>x"7f00", 14=>x"7e00", 15=>x"8300", 16=>x"8000",
---- 17=>x"7f00", 18=>x"8100", 19=>x"8000", 20=>x"8200",
---- 21=>x"8100", 22=>x"7e00", 23=>x"7f00", 24=>x"8300",
---- 25=>x"8400", 26=>x"8100", 27=>x"8100", 28=>x"8100",
---- 29=>x"8200", 30=>x"8200", 31=>x"7f00", 32=>x"8300",
---- 33=>x"8300", 34=>x"8200", 35=>x"7e00", 36=>x"8600",
---- 37=>x"8100", 38=>x"8100", 39=>x"7f00", 40=>x"8900",
---- 41=>x"8000", 42=>x"8100", 43=>x"7e00", 44=>x"8200",
---- 45=>x"8200", 46=>x"8100", 47=>x"8100", 48=>x"8100",
---- 49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7f00",
---- 53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"8100",
---- 57=>x"7e00", 58=>x"7f00", 59=>x"7f00", 60=>x"7f00",
---- 61=>x"7d00", 62=>x"8000", 63=>x"7f00", 64=>x"8000",
---- 65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"7f00",
---- 69=>x"8100", 70=>x"8000", 71=>x"8000", 72=>x"7f00",
---- 73=>x"8000", 74=>x"8100", 75=>x"8000", 76=>x"7e00",
---- 77=>x"8100", 78=>x"7f00", 79=>x"7f00", 80=>x"7d00",
---- 81=>x"8100", 82=>x"7f00", 83=>x"7c00", 84=>x"8300",
---- 85=>x"8000", 86=>x"7e00", 87=>x"7f00", 88=>x"7f00",
---- 89=>x"7f00", 90=>x"7e00", 91=>x"8000", 92=>x"7d00",
---- 93=>x"7d00", 94=>x"7c00", 95=>x"7f00", 96=>x"7c00",
---- 97=>x"7c00", 98=>x"7d00", 99=>x"7d00", 100=>x"7900",
---- 101=>x"7a00", 102=>x"7c00", 103=>x"7a00", 104=>x"7500",
---- 105=>x"7600", 106=>x"7900", 107=>x"7800", 108=>x"7200",
---- 109=>x"7000", 110=>x"7700", 111=>x"7800", 112=>x"a500",
---- 113=>x"7c00", 114=>x"6f00", 115=>x"7300", 116=>x"c600",
---- 117=>x"bb00", 118=>x"8e00", 119=>x"9100", 120=>x"c300",
---- 121=>x"cb00", 122=>x"c400", 123=>x"a200", 124=>x"c600",
---- 125=>x"c500", 126=>x"ca00", 127=>x"c800", 128=>x"c500",
---- 129=>x"c400", 130=>x"c400", 131=>x"c200", 132=>x"c500",
---- 133=>x"c300", 134=>x"c400", 135=>x"c500", 136=>x"c400",
---- 137=>x"c300", 138=>x"c700", 139=>x"c500", 140=>x"c300",
---- 141=>x"c600", 142=>x"c500", 143=>x"c400", 144=>x"c400",
---- 145=>x"c400", 146=>x"c400", 147=>x"c400", 148=>x"c400",
---- 149=>x"c400", 150=>x"c400", 151=>x"c000", 152=>x"c300",
---- 153=>x"c300", 154=>x"c500", 155=>x"c000", 156=>x"c300",
---- 157=>x"c000", 158=>x"c000", 159=>x"bc00", 160=>x"ba00",
---- 161=>x"b900", 162=>x"b900", 163=>x"b900", 164=>x"b800",
---- 165=>x"bc00", 166=>x"cb00", 167=>x"d300", 168=>x"ce00",
---- 169=>x"d400", 170=>x"d300", 171=>x"d500", 172=>x"d500",
---- 173=>x"d200", 174=>x"cd00", 175=>x"cd00", 176=>x"d200",
---- 177=>x"ce00", 178=>x"c800", 179=>x"3500", 180=>x"cb00",
---- 181=>x"cd00", 182=>x"d000", 183=>x"c900", 184=>x"d500",
---- 185=>x"d000", 186=>x"cd00", 187=>x"cb00", 188=>x"d000",
---- 189=>x"d000", 190=>x"cc00", 191=>x"c900", 192=>x"cc00",
---- 193=>x"c500", 194=>x"c500", 195=>x"c400", 196=>x"c300",
---- 197=>x"c200", 198=>x"c300", 199=>x"c700", 200=>x"c400",
---- 201=>x"cb00", 202=>x"c600", 203=>x"c200", 204=>x"ca00",
---- 205=>x"c000", 206=>x"c400", 207=>x"c500", 208=>x"c400",
---- 209=>x"c800", 210=>x"cc00", 211=>x"cb00", 212=>x"cc00",
---- 213=>x"cd00", 214=>x"ce00", 215=>x"cc00", 216=>x"c900",
---- 217=>x"cd00", 218=>x"cc00", 219=>x"ce00", 220=>x"c500",
---- 221=>x"c900", 222=>x"cc00", 223=>x"cb00", 224=>x"c700",
---- 225=>x"c600", 226=>x"cd00", 227=>x"ce00", 228=>x"c300",
---- 229=>x"cc00", 230=>x"c700", 231=>x"3100", 232=>x"c400",
---- 233=>x"c600", 234=>x"c500", 235=>x"c400", 236=>x"c400",
---- 237=>x"c000", 238=>x"c600", 239=>x"c600", 240=>x"c400",
---- 241=>x"c100", 242=>x"c000", 243=>x"c200", 244=>x"be00",
---- 245=>x"be00", 246=>x"bb00", 247=>x"b700", 248=>x"ba00",
---- 249=>x"b100", 250=>x"c100", 251=>x"c300", 252=>x"b400",
---- 253=>x"c600", 254=>x"c900", 255=>x"ca00", 256=>x"c000",
---- 257=>x"c400", 258=>x"c800", 259=>x"c700", 260=>x"bc00",
---- 261=>x"be00", 262=>x"c500", 263=>x"c800", 264=>x"b500",
---- 265=>x"bc00", 266=>x"c100", 267=>x"c300", 268=>x"b800",
---- 269=>x"b400", 270=>x"bc00", 271=>x"bf00", 272=>x"c100",
---- 273=>x"b900", 274=>x"b800", 275=>x"c000", 276=>x"b200",
---- 277=>x"bd00", 278=>x"bd00", 279=>x"b500", 280=>x"af00",
---- 281=>x"ae00", 282=>x"b400", 283=>x"ba00", 284=>x"b700",
---- 285=>x"b500", 286=>x"a700", 287=>x"b500", 288=>x"af00",
---- 289=>x"b700", 290=>x"b500", 291=>x"af00", 292=>x"b800",
---- 293=>x"ac00", 294=>x"b900", 295=>x"c300", 296=>x"ac00",
---- 297=>x"b500", 298=>x"4900", 299=>x"bc00", 300=>x"a800",
---- 301=>x"ac00", 302=>x"b200", 303=>x"ae00", 304=>x"a900",
---- 305=>x"a800", 306=>x"a900", 307=>x"ad00", 308=>x"a800",
---- 309=>x"a000", 310=>x"a800", 311=>x"ae00", 312=>x"ac00",
---- 313=>x"ac00", 314=>x"aa00", 315=>x"a800", 316=>x"a400",
---- 317=>x"ac00", 318=>x"a100", 319=>x"9500", 320=>x"9900",
---- 321=>x"9800", 322=>x"a100", 323=>x"a300", 324=>x"a600",
---- 325=>x"a100", 326=>x"a300", 327=>x"a600", 328=>x"a800",
---- 329=>x"a700", 330=>x"5c00", 331=>x"a800", 332=>x"aa00",
---- 333=>x"9d00", 334=>x"a500", 335=>x"a900", 336=>x"a100",
---- 337=>x"a200", 338=>x"a000", 339=>x"9e00", 340=>x"9d00",
---- 341=>x"a300", 342=>x"a400", 343=>x"a300", 344=>x"8f00",
---- 345=>x"8900", 346=>x"9300", 347=>x"9900", 348=>x"a700",
---- 349=>x"9900", 350=>x"6300", 351=>x"9100", 352=>x"7500",
---- 353=>x"8700", 354=>x"9100", 355=>x"9700", 356=>x"5600",
---- 357=>x"5d00", 358=>x"4a00", 359=>x"4f00", 360=>x"7800",
---- 361=>x"4000", 362=>x"be00", 363=>x"4900", 364=>x"4700",
---- 365=>x"3f00", 366=>x"4600", 367=>x"5400", 368=>x"4f00",
---- 369=>x"4400", 370=>x"4800", 371=>x"4f00", 372=>x"3900",
---- 373=>x"3000", 374=>x"4900", 375=>x"6400", 376=>x"5700",
---- 377=>x"3800", 378=>x"4400", 379=>x"6d00", 380=>x"4900",
---- 381=>x"2500", 382=>x"4000", 383=>x"5b00", 384=>x"2700",
---- 385=>x"2100", 386=>x"4e00", 387=>x"6100", 388=>x"2b00",
---- 389=>x"2500", 390=>x"5d00", 391=>x"5a00", 392=>x"2f00",
---- 393=>x"2600", 394=>x"6400", 395=>x"4100", 396=>x"1d00",
---- 397=>x"2b00", 398=>x"7d00", 399=>x"7000", 400=>x"1400",
---- 401=>x"5200", 402=>x"a700", 403=>x"a700", 404=>x"2600",
---- 405=>x"8900", 406=>x"6a00", 407=>x"7400", 408=>x"6d00",
---- 409=>x"8000", 410=>x"6a00", 411=>x"6a00", 412=>x"8d00",
---- 413=>x"5400", 414=>x"6600", 415=>x"8a00", 416=>x"7d00",
---- 417=>x"6000", 418=>x"9800", 419=>x"a800", 420=>x"7900",
---- 421=>x"9300", 422=>x"b100", 423=>x"a900", 424=>x"7700",
---- 425=>x"8f00", 426=>x"9500", 427=>x"a800", 428=>x"8a00",
---- 429=>x"9f00", 430=>x"a500", 431=>x"b000", 432=>x"a000",
---- 433=>x"bb00", 434=>x"b000", 435=>x"b500", 436=>x"ac00",
---- 437=>x"b800", 438=>x"b600", 439=>x"b600", 440=>x"bb00",
---- 441=>x"b300", 442=>x"b400", 443=>x"bb00", 444=>x"b700",
---- 445=>x"b600", 446=>x"ab00", 447=>x"bc00", 448=>x"a600",
---- 449=>x"a900", 450=>x"a700", 451=>x"be00", 452=>x"b000",
---- 453=>x"a100", 454=>x"ac00", 455=>x"bf00", 456=>x"b100",
---- 457=>x"ad00", 458=>x"b400", 459=>x"bf00", 460=>x"a500",
---- 461=>x"a600", 462=>x"b900", 463=>x"c300", 464=>x"a000",
---- 465=>x"a600", 466=>x"ba00", 467=>x"c900", 468=>x"a100",
---- 469=>x"b300", 470=>x"c000", 471=>x"c000", 472=>x"9d00",
---- 473=>x"bc00", 474=>x"c000", 475=>x"5200", 476=>x"a700",
---- 477=>x"4500", 478=>x"ab00", 479=>x"a800", 480=>x"b400",
---- 481=>x"b100", 482=>x"a900", 483=>x"a200", 484=>x"b900",
---- 485=>x"a900", 486=>x"8a00", 487=>x"8400", 488=>x"9100",
---- 489=>x"5600", 490=>x"5300", 491=>x"9200", 492=>x"5200",
---- 493=>x"5800", 494=>x"6300", 495=>x"6300", 496=>x"8800",
---- 497=>x"8e00", 498=>x"8a00", 499=>x"8000", 500=>x"9a00",
---- 501=>x"9700", 502=>x"9500", 503=>x"9f00", 504=>x"9100",
---- 505=>x"8f00", 506=>x"7900", 507=>x"8e00", 508=>x"7700",
---- 509=>x"7d00", 510=>x"5000", 511=>x"5800", 512=>x"4d00",
---- 513=>x"4c00", 514=>x"3200", 515=>x"3800", 516=>x"3300",
---- 517=>x"3100", 518=>x"3100", 519=>x"3300", 520=>x"3000",
---- 521=>x"2e00", 522=>x"2d00", 523=>x"3400", 524=>x"2c00",
---- 525=>x"3000", 526=>x"3400", 527=>x"4c00", 528=>x"2300",
---- 529=>x"3000", 530=>x"4c00", 531=>x"5000", 532=>x"3200",
---- 533=>x"3000", 534=>x"6000", 535=>x"3300", 536=>x"5900",
---- 537=>x"5600", 538=>x"4600", 539=>x"4c00", 540=>x"3e00",
---- 541=>x"4000", 542=>x"4d00", 543=>x"9c00", 544=>x"6100",
---- 545=>x"6e00", 546=>x"a200", 547=>x"c600", 548=>x"9400",
---- 549=>x"9d00", 550=>x"a900", 551=>x"b400", 552=>x"7100",
---- 553=>x"7900", 554=>x"8c00", 555=>x"8d00", 556=>x"6700",
---- 557=>x"7200", 558=>x"8800", 559=>x"7e00", 560=>x"7e00",
---- 561=>x"8300", 562=>x"8800", 563=>x"8a00", 564=>x"8d00",
---- 565=>x"8d00", 566=>x"8d00", 567=>x"9400", 568=>x"9600",
---- 569=>x"9900", 570=>x"9c00", 571=>x"a100", 572=>x"a400",
---- 573=>x"a300", 574=>x"ab00", 575=>x"ad00", 576=>x"a700",
---- 577=>x"a700", 578=>x"ac00", 579=>x"af00", 580=>x"b000",
---- 581=>x"ad00", 582=>x"ad00", 583=>x"ab00", 584=>x"b200",
---- 585=>x"b100", 586=>x"b200", 587=>x"af00", 588=>x"b000",
---- 589=>x"b200", 590=>x"b100", 591=>x"b000", 592=>x"b300",
---- 593=>x"b000", 594=>x"ae00", 595=>x"af00", 596=>x"b700",
---- 597=>x"b800", 598=>x"af00", 599=>x"ac00", 600=>x"af00",
---- 601=>x"b400", 602=>x"b100", 603=>x"ad00", 604=>x"af00",
---- 605=>x"b300", 606=>x"b100", 607=>x"ab00", 608=>x"ad00",
---- 609=>x"af00", 610=>x"b000", 611=>x"5500", 612=>x"a800",
---- 613=>x"aa00", 614=>x"ac00", 615=>x"ac00", 616=>x"a700",
---- 617=>x"a800", 618=>x"a800", 619=>x"a900", 620=>x"a400",
---- 621=>x"a600", 622=>x"a500", 623=>x"a800", 624=>x"9e00",
---- 625=>x"a300", 626=>x"a500", 627=>x"a400", 628=>x"9f00",
---- 629=>x"a100", 630=>x"a300", 631=>x"a000", 632=>x"9d00",
---- 633=>x"9e00", 634=>x"9f00", 635=>x"a000", 636=>x"9d00",
---- 637=>x"9d00", 638=>x"9f00", 639=>x"a100", 640=>x"9c00",
---- 641=>x"9b00", 642=>x"9c00", 643=>x"a000", 644=>x"9a00",
---- 645=>x"9b00", 646=>x"9d00", 647=>x"9e00", 648=>x"9b00",
---- 649=>x"9b00", 650=>x"9f00", 651=>x"9d00", 652=>x"9b00",
---- 653=>x"9900", 654=>x"9c00", 655=>x"9c00", 656=>x"9b00",
---- 657=>x"9600", 658=>x"9700", 659=>x"6200", 660=>x"9b00",
---- 661=>x"9900", 662=>x"9b00", 663=>x"9b00", 664=>x"9a00",
---- 665=>x"9a00", 666=>x"9b00", 667=>x"9c00", 668=>x"9900",
---- 669=>x"9900", 670=>x"9a00", 671=>x"9c00", 672=>x"9700",
---- 673=>x"9700", 674=>x"9800", 675=>x"6600", 676=>x"9200",
---- 677=>x"9600", 678=>x"9500", 679=>x"9700", 680=>x"8c00",
---- 681=>x"9100", 682=>x"9400", 683=>x"9500", 684=>x"8c00",
---- 685=>x"8e00", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
---- 689=>x"8e00", 690=>x"8900", 691=>x"8c00", 692=>x"8a00",
---- 693=>x"8a00", 694=>x"8700", 695=>x"8400", 696=>x"8800",
---- 697=>x"6d00", 698=>x"6300", 699=>x"8f00", 700=>x"8200",
---- 701=>x"5c00", 702=>x"5000", 703=>x"5100", 704=>x"8300",
---- 705=>x"7600", 706=>x"7a00", 707=>x"7400", 708=>x"8e00",
---- 709=>x"8b00", 710=>x"8100", 711=>x"8100", 712=>x"9600",
---- 713=>x"8f00", 714=>x"8500", 715=>x"8100", 716=>x"9300",
---- 717=>x"9000", 718=>x"8a00", 719=>x"8800", 720=>x"9300",
---- 721=>x"9000", 722=>x"8c00", 723=>x"8800", 724=>x"8c00",
---- 725=>x"8e00", 726=>x"8e00", 727=>x"8900", 728=>x"8b00",
---- 729=>x"8f00", 730=>x"8d00", 731=>x"8b00", 732=>x"8c00",
---- 733=>x"8e00", 734=>x"8c00", 735=>x"8b00", 736=>x"8900",
---- 737=>x"8d00", 738=>x"8900", 739=>x"8900", 740=>x"8800",
---- 741=>x"8b00", 742=>x"8900", 743=>x"8a00", 744=>x"8a00",
---- 745=>x"8b00", 746=>x"8b00", 747=>x"7100", 748=>x"8a00",
---- 749=>x"8a00", 750=>x"8e00", 751=>x"8d00", 752=>x"8900",
---- 753=>x"8b00", 754=>x"9100", 755=>x"9200", 756=>x"8600",
---- 757=>x"8c00", 758=>x"9100", 759=>x"9100", 760=>x"8700",
---- 761=>x"8900", 762=>x"8b00", 763=>x"9200", 764=>x"8100",
---- 765=>x"8000", 766=>x"8800", 767=>x"8a00", 768=>x"6b00",
---- 769=>x"7100", 770=>x"7800", 771=>x"7c00", 772=>x"6600",
---- 773=>x"7200", 774=>x"7900", 775=>x"7900", 776=>x"8500",
---- 777=>x"8400", 778=>x"8700", 779=>x"8900", 780=>x"8a00",
---- 781=>x"8900", 782=>x"8800", 783=>x"8e00", 784=>x"8600",
---- 785=>x"8400", 786=>x"8600", 787=>x"8800", 788=>x"8500",
---- 789=>x"8500", 790=>x"8a00", 791=>x"8a00", 792=>x"8500",
---- 793=>x"8900", 794=>x"8a00", 795=>x"8b00", 796=>x"8a00",
---- 797=>x"8900", 798=>x"8800", 799=>x"8800", 800=>x"8700",
---- 801=>x"8700", 802=>x"8700", 803=>x"8800", 804=>x"8100",
---- 805=>x"8700", 806=>x"8600", 807=>x"8b00", 808=>x"8400",
---- 809=>x"8800", 810=>x"8b00", 811=>x"8d00", 812=>x"8700",
---- 813=>x"8900", 814=>x"8d00", 815=>x"8f00", 816=>x"8800",
---- 817=>x"8800", 818=>x"8c00", 819=>x"8d00", 820=>x"8b00",
---- 821=>x"8700", 822=>x"8700", 823=>x"8a00", 824=>x"8b00",
---- 825=>x"8800", 826=>x"8a00", 827=>x"8d00", 828=>x"8a00",
---- 829=>x"8a00", 830=>x"8c00", 831=>x"8c00", 832=>x"8a00",
---- 833=>x"8a00", 834=>x"8c00", 835=>x"8a00", 836=>x"8d00",
---- 837=>x"8a00", 838=>x"8d00", 839=>x"8a00", 840=>x"8a00",
---- 841=>x"8d00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
---- 845=>x"8b00", 846=>x"8d00", 847=>x"8b00", 848=>x"8a00",
---- 849=>x"8700", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
---- 853=>x"8800", 854=>x"7400", 855=>x"8d00", 856=>x"8c00",
---- 857=>x"8900", 858=>x"8900", 859=>x"8b00", 860=>x"8b00",
---- 861=>x"8b00", 862=>x"8400", 863=>x"8900", 864=>x"7500",
---- 865=>x"8a00", 866=>x"8900", 867=>x"8700", 868=>x"8800",
---- 869=>x"8700", 870=>x"8800", 871=>x"8b00", 872=>x"8800",
---- 873=>x"8800", 874=>x"8700", 875=>x"8900", 876=>x"8a00",
---- 877=>x"8900", 878=>x"8700", 879=>x"8900", 880=>x"8900",
---- 881=>x"8800", 882=>x"8800", 883=>x"8900", 884=>x"8a00",
---- 885=>x"8800", 886=>x"8900", 887=>x"8800", 888=>x"8a00",
---- 889=>x"8b00", 890=>x"8b00", 891=>x"8900", 892=>x"8a00",
---- 893=>x"8800", 894=>x"8a00", 895=>x"8b00", 896=>x"8c00",
---- 897=>x"8b00", 898=>x"8c00", 899=>x"8800", 900=>x"8f00",
---- 901=>x"8d00", 902=>x"8900", 903=>x"8700", 904=>x"8d00",
---- 905=>x"8c00", 906=>x"8d00", 907=>x"8a00", 908=>x"8a00",
---- 909=>x"8a00", 910=>x"8a00", 911=>x"7600", 912=>x"8b00",
---- 913=>x"8a00", 914=>x"8a00", 915=>x"8a00", 916=>x"8b00",
---- 917=>x"8a00", 918=>x"8c00", 919=>x"8d00", 920=>x"8c00",
---- 921=>x"8c00", 922=>x"8d00", 923=>x"7100", 924=>x"8f00",
---- 925=>x"8d00", 926=>x"8c00", 927=>x"8e00", 928=>x"8b00",
---- 929=>x"8e00", 930=>x"8f00", 931=>x"8d00", 932=>x"8c00",
---- 933=>x"8f00", 934=>x"8d00", 935=>x"8900", 936=>x"8c00",
---- 937=>x"8e00", 938=>x"8e00", 939=>x"8c00", 940=>x"8f00",
---- 941=>x"8f00", 942=>x"9000", 943=>x"8b00", 944=>x"8e00",
---- 945=>x"9000", 946=>x"8e00", 947=>x"8d00", 948=>x"9000",
---- 949=>x"9000", 950=>x"9000", 951=>x"8e00", 952=>x"8f00",
---- 953=>x"9100", 954=>x"9000", 955=>x"8e00", 956=>x"8f00",
---- 957=>x"8e00", 958=>x"8f00", 959=>x"8f00", 960=>x"8f00",
---- 961=>x"8e00", 962=>x"8e00", 963=>x"8d00", 964=>x"9000",
---- 965=>x"9100", 966=>x"8d00", 967=>x"8b00", 968=>x"9100",
---- 969=>x"9000", 970=>x"8d00", 971=>x"8c00", 972=>x"8e00",
---- 973=>x"8e00", 974=>x"8f00", 975=>x"9100", 976=>x"8f00",
---- 977=>x"8f00", 978=>x"9000", 979=>x"9100", 980=>x"8d00",
---- 981=>x"8f00", 982=>x"8f00", 983=>x"8f00", 984=>x"8c00",
---- 985=>x"8d00", 986=>x"9200", 987=>x"8f00", 988=>x"8e00",
---- 989=>x"8d00", 990=>x"9100", 991=>x"8f00", 992=>x"8f00",
---- 993=>x"8d00", 994=>x"8b00", 995=>x"8e00", 996=>x"8f00",
---- 997=>x"8c00", 998=>x"8d00", 999=>x"8d00", 1000=>x"8d00",
---- 1001=>x"8d00", 1002=>x"8e00", 1003=>x"8d00", 1004=>x"8c00",
---- 1005=>x"8b00", 1006=>x"8d00", 1007=>x"8a00", 1008=>x"8d00",
---- 1009=>x"8b00", 1010=>x"8d00", 1011=>x"8c00", 1012=>x"7100",
---- 1013=>x"8a00", 1014=>x"8c00", 1015=>x"8f00", 1016=>x"8c00",
---- 1017=>x"8d00", 1018=>x"8b00", 1019=>x"8e00", 1020=>x"8b00",
---- 1021=>x"8d00", 1022=>x"8d00", 1023=>x"8b00"),
----
---- 34 => (0=>x"8000", 1=>x"8200", 2=>x"8100", 3=>x"8600", 4=>x"8000",
---- 5=>x"8200", 6=>x"8100", 7=>x"8600", 8=>x"8000",
---- 9=>x"8200", 10=>x"8000", 11=>x"8600", 12=>x"7f00",
---- 13=>x"8000", 14=>x"8000", 15=>x"8000", 16=>x"7f00",
---- 17=>x"7f00", 18=>x"7f00", 19=>x"8000", 20=>x"8000",
---- 21=>x"8000", 22=>x"8000", 23=>x"8000", 24=>x"8000",
---- 25=>x"8100", 26=>x"8200", 27=>x"8100", 28=>x"8000",
---- 29=>x"8100", 30=>x"7f00", 31=>x"7f00", 32=>x"8200",
---- 33=>x"8100", 34=>x"7f00", 35=>x"7f00", 36=>x"7f00",
---- 37=>x"8300", 38=>x"8200", 39=>x"8200", 40=>x"8100",
---- 41=>x"8000", 42=>x"8000", 43=>x"8200", 44=>x"8000",
---- 45=>x"8200", 46=>x"7e00", 47=>x"7c00", 48=>x"7f00",
---- 49=>x"8200", 50=>x"8000", 51=>x"7f00", 52=>x"7d00",
---- 53=>x"7f00", 54=>x"8000", 55=>x"7e00", 56=>x"8000",
---- 57=>x"8000", 58=>x"8000", 59=>x"8000", 60=>x"7d00",
---- 61=>x"8200", 62=>x"7f00", 63=>x"8000", 64=>x"7c00",
---- 65=>x"8200", 66=>x"8000", 67=>x"7d00", 68=>x"8000",
---- 69=>x"8300", 70=>x"7e00", 71=>x"7e00", 72=>x"8000",
---- 73=>x"7f00", 74=>x"8000", 75=>x"7e00", 76=>x"8000",
---- 77=>x"8200", 78=>x"8100", 79=>x"7f00", 80=>x"7f00",
---- 81=>x"8000", 82=>x"7f00", 83=>x"7f00", 84=>x"7b00",
---- 85=>x"7e00", 86=>x"8200", 87=>x"7a00", 88=>x"7e00",
---- 89=>x"8100", 90=>x"8100", 91=>x"8200", 92=>x"7f00",
---- 93=>x"8100", 94=>x"8200", 95=>x"8100", 96=>x"7f00",
---- 97=>x"8200", 98=>x"8200", 99=>x"8100", 100=>x"7e00",
---- 101=>x"8200", 102=>x"8300", 103=>x"8200", 104=>x"7d00",
---- 105=>x"7d00", 106=>x"7f00", 107=>x"7f00", 108=>x"7800",
---- 109=>x"7b00", 110=>x"7c00", 111=>x"7e00", 112=>x"7500",
---- 113=>x"7600", 114=>x"7e00", 115=>x"7c00", 116=>x"6c00",
---- 117=>x"7600", 118=>x"7c00", 119=>x"7900", 120=>x"7800",
---- 121=>x"6c00", 122=>x"8800", 123=>x"7300", 124=>x"b800",
---- 125=>x"8f00", 126=>x"7000", 127=>x"6d00", 128=>x"c900",
---- 129=>x"c400", 130=>x"9f00", 131=>x"7400", 132=>x"c300",
---- 133=>x"c100", 134=>x"c500", 135=>x"b500", 136=>x"c100",
---- 137=>x"c300", 138=>x"c200", 139=>x"c900", 140=>x"c300",
---- 141=>x"c500", 142=>x"c600", 143=>x"c900", 144=>x"c300",
---- 145=>x"c300", 146=>x"c500", 147=>x"ca00", 148=>x"c300",
---- 149=>x"c600", 150=>x"c800", 151=>x"c600", 152=>x"c100",
---- 153=>x"c100", 154=>x"bc00", 155=>x"b800", 156=>x"b800",
---- 157=>x"bc00", 158=>x"be00", 159=>x"cb00", 160=>x"c500",
---- 161=>x"d100", 162=>x"d400", 163=>x"d400", 164=>x"d800",
---- 165=>x"d300", 166=>x"d300", 167=>x"d200", 168=>x"d300",
---- 169=>x"cf00", 170=>x"cf00", 171=>x"d300", 172=>x"ce00",
---- 173=>x"d000", 174=>x"d100", 175=>x"cf00", 176=>x"d000",
---- 177=>x"ce00", 178=>x"cf00", 179=>x"d000", 180=>x"ce00",
---- 181=>x"d100", 182=>x"ce00", 183=>x"cf00", 184=>x"c900",
---- 185=>x"cf00", 186=>x"ce00", 187=>x"cb00", 188=>x"c500",
---- 189=>x"c100", 190=>x"c400", 191=>x"cb00", 192=>x"ca00",
---- 193=>x"c700", 194=>x"c700", 195=>x"cf00", 196=>x"2e00",
---- 197=>x"d100", 198=>x"c900", 199=>x"c700", 200=>x"c700",
---- 201=>x"c800", 202=>x"c900", 203=>x"ca00", 204=>x"cd00",
---- 205=>x"c400", 206=>x"cb00", 207=>x"d300", 208=>x"ce00",
---- 209=>x"d100", 210=>x"c500", 211=>x"cd00", 212=>x"c500",
---- 213=>x"ce00", 214=>x"d100", 215=>x"c800", 216=>x"cd00",
---- 217=>x"c800", 218=>x"d400", 219=>x"ce00", 220=>x"cf00",
---- 221=>x"ca00", 222=>x"c900", 223=>x"d100", 224=>x"cd00",
---- 225=>x"cc00", 226=>x"c600", 227=>x"3300", 228=>x"cd00",
---- 229=>x"ca00", 230=>x"c800", 231=>x"cc00", 232=>x"ca00",
---- 233=>x"ce00", 234=>x"c700", 235=>x"c500", 236=>x"c700",
---- 237=>x"c800", 238=>x"bf00", 239=>x"be00", 240=>x"bf00",
---- 241=>x"bb00", 242=>x"c200", 243=>x"cb00", 244=>x"be00",
---- 245=>x"c700", 246=>x"c900", 247=>x"cb00", 248=>x"c400",
---- 249=>x"c900", 250=>x"c800", 251=>x"c300", 252=>x"c400",
---- 253=>x"c400", 254=>x"c600", 255=>x"c500", 256=>x"c900",
---- 257=>x"c200", 258=>x"c000", 259=>x"c800", 260=>x"c800",
---- 261=>x"c500", 262=>x"bd00", 263=>x"c100", 264=>x"c300",
---- 265=>x"c600", 266=>x"c600", 267=>x"c300", 268=>x"c000",
---- 269=>x"c600", 270=>x"c500", 271=>x"c100", 272=>x"c100",
---- 273=>x"bc00", 274=>x"c200", 275=>x"be00", 276=>x"b600",
---- 277=>x"c000", 278=>x"be00", 279=>x"c000", 280=>x"ac00",
---- 281=>x"b400", 282=>x"c100", 283=>x"c600", 284=>x"ba00",
---- 285=>x"b400", 286=>x"bd00", 287=>x"b900", 288=>x"bf00",
---- 289=>x"bc00", 290=>x"c100", 291=>x"b000", 292=>x"c100",
---- 293=>x"bc00", 294=>x"b400", 295=>x"af00", 296=>x"b700",
---- 297=>x"b000", 298=>x"b200", 299=>x"b800", 300=>x"af00",
---- 301=>x"b900", 302=>x"bc00", 303=>x"b700", 304=>x"b300",
---- 305=>x"b600", 306=>x"ba00", 307=>x"b800", 308=>x"b200",
---- 309=>x"b300", 310=>x"a900", 311=>x"a800", 312=>x"a400",
---- 313=>x"a100", 314=>x"ab00", 315=>x"aa00", 316=>x"a100",
---- 317=>x"a900", 318=>x"af00", 319=>x"af00", 320=>x"a900",
---- 321=>x"a900", 322=>x"a800", 323=>x"af00", 324=>x"a500",
---- 325=>x"aa00", 326=>x"aa00", 327=>x"a700", 328=>x"a300",
---- 329=>x"9f00", 330=>x"aa00", 331=>x"aa00", 332=>x"ab00",
---- 333=>x"a400", 334=>x"a100", 335=>x"a700", 336=>x"a400",
---- 337=>x"a900", 338=>x"a500", 339=>x"9d00", 340=>x"a100",
---- 341=>x"a400", 342=>x"a600", 343=>x"9c00", 344=>x"9b00",
---- 345=>x"a500", 346=>x"a300", 347=>x"a300", 348=>x"7400",
---- 349=>x"8d00", 350=>x"9300", 351=>x"9500", 352=>x"7e00",
---- 353=>x"6a00", 354=>x"6b00", 355=>x"5200", 356=>x"5000",
---- 357=>x"4d00", 358=>x"4a00", 359=>x"3800", 360=>x"3500",
---- 361=>x"3300", 362=>x"3400", 363=>x"3000", 364=>x"3400",
---- 365=>x"2b00", 366=>x"2900", 367=>x"2200", 368=>x"3800",
---- 369=>x"3300", 370=>x"2800", 371=>x"2200", 372=>x"2b00",
---- 373=>x"2a00", 374=>x"2c00", 375=>x"2300", 376=>x"2300",
---- 377=>x"2100", 378=>x"2100", 379=>x"2d00", 380=>x"1e00",
---- 381=>x"1f00", 382=>x"1e00", 383=>x"5c00", 384=>x"2c00",
---- 385=>x"2200", 386=>x"9b00", 387=>x"ae00", 388=>x"4000",
---- 389=>x"7300", 390=>x"b200", 391=>x"9b00", 392=>x"8100",
---- 393=>x"b100", 394=>x"9500", 395=>x"7500", 396=>x"a900",
---- 397=>x"8800", 398=>x"7500", 399=>x"8f00", 400=>x"7b00",
---- 401=>x"7000", 402=>x"9100", 403=>x"bb00", 404=>x"7700",
---- 405=>x"9a00", 406=>x"bd00", 407=>x"c400", 408=>x"a400",
---- 409=>x"c200", 410=>x"c600", 411=>x"c200", 412=>x"c100",
---- 413=>x"bf00", 414=>x"c300", 415=>x"c100", 416=>x"bb00",
---- 417=>x"be00", 418=>x"bd00", 419=>x"ba00", 420=>x"ba00",
---- 421=>x"b700", 422=>x"b300", 423=>x"b800", 424=>x"b600",
---- 425=>x"ae00", 426=>x"5000", 427=>x"b500", 428=>x"b200",
---- 429=>x"b000", 430=>x"b600", 431=>x"b900", 432=>x"b400",
---- 433=>x"b900", 434=>x"bd00", 435=>x"b900", 436=>x"ba00",
---- 437=>x"bc00", 438=>x"bb00", 439=>x"b400", 440=>x"bf00",
---- 441=>x"c300", 442=>x"bb00", 443=>x"af00", 444=>x"bf00",
---- 445=>x"bc00", 446=>x"b300", 447=>x"a800", 448=>x"b500",
---- 449=>x"b200", 450=>x"b100", 451=>x"a900", 452=>x"ba00",
---- 453=>x"b600", 454=>x"ab00", 455=>x"aa00", 456=>x"c200",
---- 457=>x"b500", 458=>x"a800", 459=>x"a900", 460=>x"c500",
---- 461=>x"b100", 462=>x"a700", 463=>x"ac00", 464=>x"bc00",
---- 465=>x"a900", 466=>x"a400", 467=>x"a400", 468=>x"ae00",
---- 469=>x"a200", 470=>x"9d00", 471=>x"a400", 472=>x"a200",
---- 473=>x"9b00", 474=>x"9800", 475=>x"9c00", 476=>x"9e00",
---- 477=>x"9a00", 478=>x"9c00", 479=>x"a300", 480=>x"9a00",
---- 481=>x"9e00", 482=>x"a600", 483=>x"a600", 484=>x"9200",
---- 485=>x"9a00", 486=>x"9d00", 487=>x"a300", 488=>x"7600",
---- 489=>x"8200", 490=>x"8e00", 491=>x"9400", 492=>x"5f00",
---- 493=>x"6600", 494=>x"6100", 495=>x"6500", 496=>x"7400",
---- 497=>x"6c00", 498=>x"5900", 499=>x"4400", 500=>x"9a00",
---- 501=>x"8d00", 502=>x"7800", 503=>x"6300", 504=>x"a500",
---- 505=>x"9b00", 506=>x"8400", 507=>x"7800", 508=>x"9a00",
---- 509=>x"8800", 510=>x"6800", 511=>x"7400", 512=>x"6300",
---- 513=>x"4d00", 514=>x"cb00", 515=>x"4400", 516=>x"2e00",
---- 517=>x"2d00", 518=>x"2c00", 519=>x"2700", 520=>x"4500",
---- 521=>x"4c00", 522=>x"3300", 523=>x"2a00", 524=>x"8800",
---- 525=>x"9e00", 526=>x"6b00", 527=>x"3900", 528=>x"a800",
---- 529=>x"cf00", 530=>x"b300", 531=>x"8d00", 532=>x"9400",
---- 533=>x"d200", 534=>x"c700", 535=>x"c500", 536=>x"ba00",
---- 537=>x"d400", 538=>x"cf00", 539=>x"cc00", 540=>x"d100",
---- 541=>x"ce00", 542=>x"ce00", 543=>x"c900", 544=>x"c900",
---- 545=>x"ce00", 546=>x"cf00", 547=>x"be00", 548=>x"be00",
---- 549=>x"c500", 550=>x"be00", 551=>x"b200", 552=>x"9200",
---- 553=>x"9400", 554=>x"9600", 555=>x"ae00", 556=>x"6f00",
---- 557=>x"7200", 558=>x"8100", 559=>x"9d00", 560=>x"8100",
---- 561=>x"9000", 562=>x"9400", 563=>x"9b00", 564=>x"9800",
---- 565=>x"9a00", 566=>x"a100", 567=>x"a200", 568=>x"a200",
---- 569=>x"a800", 570=>x"a800", 571=>x"a600", 572=>x"ab00",
---- 573=>x"ad00", 574=>x"a400", 575=>x"aa00", 576=>x"aa00",
---- 577=>x"a600", 578=>x"a900", 579=>x"a900", 580=>x"a700",
---- 581=>x"af00", 582=>x"b000", 583=>x"af00", 584=>x"ad00",
---- 585=>x"af00", 586=>x"b100", 587=>x"ad00", 588=>x"b100",
---- 589=>x"b200", 590=>x"b000", 591=>x"aa00", 592=>x"af00",
---- 593=>x"b000", 594=>x"aa00", 595=>x"a900", 596=>x"ab00",
---- 597=>x"ac00", 598=>x"ab00", 599=>x"a700", 600=>x"ad00",
---- 601=>x"ae00", 602=>x"a800", 603=>x"a400", 604=>x"aa00",
---- 605=>x"ab00", 606=>x"a800", 607=>x"a300", 608=>x"aa00",
---- 609=>x"a900", 610=>x"a600", 611=>x"a300", 612=>x"aa00",
---- 613=>x"a800", 614=>x"a400", 615=>x"a300", 616=>x"a900",
---- 617=>x"a600", 618=>x"a300", 619=>x"a000", 620=>x"a500",
---- 621=>x"a400", 622=>x"5b00", 623=>x"a100", 624=>x"a000",
---- 625=>x"a300", 626=>x"a100", 627=>x"9e00", 628=>x"5b00",
---- 629=>x"a200", 630=>x"9d00", 631=>x"6600", 632=>x"a100",
---- 633=>x"a100", 634=>x"9c00", 635=>x"9800", 636=>x"9e00",
---- 637=>x"9e00", 638=>x"9e00", 639=>x"9400", 640=>x"9f00",
---- 641=>x"9f00", 642=>x"9c00", 643=>x"9700", 644=>x"9e00",
---- 645=>x"9c00", 646=>x"9d00", 647=>x"9a00", 648=>x"9e00",
---- 649=>x"9d00", 650=>x"9f00", 651=>x"9800", 652=>x"9f00",
---- 653=>x"9c00", 654=>x"9d00", 655=>x"9c00", 656=>x"9e00",
---- 657=>x"6000", 658=>x"9d00", 659=>x"9d00", 660=>x"9b00",
---- 661=>x"9f00", 662=>x"9f00", 663=>x"9c00", 664=>x"a000",
---- 665=>x"9f00", 666=>x"9d00", 667=>x"9e00", 668=>x"9d00",
---- 669=>x"9f00", 670=>x"9d00", 671=>x"9d00", 672=>x"9600",
---- 673=>x"9a00", 674=>x"9a00", 675=>x"9c00", 676=>x"9400",
---- 677=>x"9900", 678=>x"9800", 679=>x"9a00", 680=>x"9400",
---- 681=>x"9400", 682=>x"9400", 683=>x"9a00", 684=>x"9100",
---- 685=>x"9100", 686=>x"8f00", 687=>x"9400", 688=>x"9000",
---- 689=>x"8f00", 690=>x"8c00", 691=>x"8f00", 692=>x"8700",
---- 693=>x"8700", 694=>x"8900", 695=>x"8e00", 696=>x"7a00",
---- 697=>x"7f00", 698=>x"8400", 699=>x"8900", 700=>x"5200",
---- 701=>x"5900", 702=>x"6300", 703=>x"6800", 704=>x"6700",
---- 705=>x"5e00", 706=>x"5b00", 707=>x"6000", 708=>x"7f00",
---- 709=>x"7d00", 710=>x"7c00", 711=>x"7900", 712=>x"7c00",
---- 713=>x"7f00", 714=>x"7f00", 715=>x"8100", 716=>x"8000",
---- 717=>x"7d00", 718=>x"8600", 719=>x"8000", 720=>x"8500",
---- 721=>x"8400", 722=>x"7c00", 723=>x"7a00", 724=>x"8600",
---- 725=>x"8400", 726=>x"8300", 727=>x"7e00", 728=>x"8700",
---- 729=>x"8500", 730=>x"8500", 731=>x"8200", 732=>x"8900",
---- 733=>x"8700", 734=>x"8500", 735=>x"8100", 736=>x"8800",
---- 737=>x"8900", 738=>x"8700", 739=>x"8800", 740=>x"8b00",
---- 741=>x"8c00", 742=>x"8900", 743=>x"8b00", 744=>x"8b00",
---- 745=>x"8e00", 746=>x"9300", 747=>x"9700", 748=>x"8d00",
---- 749=>x"9300", 750=>x"9500", 751=>x"9c00", 752=>x"9000",
---- 753=>x"9600", 754=>x"9800", 755=>x"a000", 756=>x"9100",
---- 757=>x"9400", 758=>x"9a00", 759=>x"9c00", 760=>x"9100",
---- 761=>x"9300", 762=>x"9600", 763=>x"9600", 764=>x"8e00",
---- 765=>x"9200", 766=>x"9300", 767=>x"9400", 768=>x"8400",
---- 769=>x"7700", 770=>x"8d00", 771=>x"9400", 772=>x"8000",
---- 773=>x"8700", 774=>x"8700", 775=>x"9000", 776=>x"8700",
---- 777=>x"9200", 778=>x"8e00", 779=>x"9d00", 780=>x"8c00",
---- 781=>x"8d00", 782=>x"9100", 783=>x"9900", 784=>x"8d00",
---- 785=>x"8e00", 786=>x"9300", 787=>x"9600", 788=>x"8a00",
---- 789=>x"8c00", 790=>x"9100", 791=>x"9300", 792=>x"8a00",
---- 793=>x"8c00", 794=>x"8e00", 795=>x"6b00", 796=>x"7300",
---- 797=>x"8b00", 798=>x"8d00", 799=>x"8e00", 800=>x"8700",
---- 801=>x"8b00", 802=>x"8d00", 803=>x"8b00", 804=>x"8a00",
---- 805=>x"8d00", 806=>x"8c00", 807=>x"8b00", 808=>x"8d00",
---- 809=>x"8f00", 810=>x"8c00", 811=>x"7500", 812=>x"8e00",
---- 813=>x"8c00", 814=>x"8d00", 815=>x"8800", 816=>x"8c00",
---- 817=>x"8d00", 818=>x"8e00", 819=>x"8900", 820=>x"8900",
---- 821=>x"8d00", 822=>x"8d00", 823=>x"8900", 824=>x"8e00",
---- 825=>x"8c00", 826=>x"8900", 827=>x"8d00", 828=>x"9000",
---- 829=>x"8a00", 830=>x"7100", 831=>x"8c00", 832=>x"8900",
---- 833=>x"8b00", 834=>x"8c00", 835=>x"8b00", 836=>x"8b00",
---- 837=>x"8b00", 838=>x"8a00", 839=>x"8f00", 840=>x"8d00",
---- 841=>x"8d00", 842=>x"8c00", 843=>x"8c00", 844=>x"8c00",
---- 845=>x"8d00", 846=>x"8d00", 847=>x"8f00", 848=>x"7100",
---- 849=>x"8e00", 850=>x"8d00", 851=>x"8d00", 852=>x"8b00",
---- 853=>x"8c00", 854=>x"8d00", 855=>x"8e00", 856=>x"8b00",
---- 857=>x"8d00", 858=>x"8d00", 859=>x"8e00", 860=>x"8a00",
---- 861=>x"8c00", 862=>x"8a00", 863=>x"8d00", 864=>x"8800",
---- 865=>x"8a00", 866=>x"8800", 867=>x"8c00", 868=>x"8800",
---- 869=>x"8700", 870=>x"8900", 871=>x"8b00", 872=>x"8800",
---- 873=>x"8a00", 874=>x"8a00", 875=>x"8a00", 876=>x"8a00",
---- 877=>x"8c00", 878=>x"8c00", 879=>x"7700", 880=>x"8900",
---- 881=>x"8800", 882=>x"8a00", 883=>x"8a00", 884=>x"8100",
---- 885=>x"8700", 886=>x"8700", 887=>x"8900", 888=>x"8400",
---- 889=>x"8600", 890=>x"8600", 891=>x"8900", 892=>x"8700",
---- 893=>x"8600", 894=>x"8500", 895=>x"8700", 896=>x"8500",
---- 897=>x"8600", 898=>x"8600", 899=>x"8800", 900=>x"8700",
---- 901=>x"8800", 902=>x"8700", 903=>x"8900", 904=>x"8700",
---- 905=>x"8a00", 906=>x"8500", 907=>x"8800", 908=>x"8b00",
---- 909=>x"8800", 910=>x"8900", 911=>x"8800", 912=>x"8a00",
---- 913=>x"8600", 914=>x"8900", 915=>x"8700", 916=>x"8c00",
---- 917=>x"7500", 918=>x"8900", 919=>x"8600", 920=>x"8e00",
---- 921=>x"8c00", 922=>x"8900", 923=>x"8700", 924=>x"8c00",
---- 925=>x"8c00", 926=>x"8700", 927=>x"8a00", 928=>x"8e00",
---- 929=>x"8c00", 930=>x"8700", 931=>x"8700", 932=>x"8c00",
---- 933=>x"7300", 934=>x"8800", 935=>x"8a00", 936=>x"8b00",
---- 937=>x"8e00", 938=>x"8900", 939=>x"8700", 940=>x"8d00",
---- 941=>x"8900", 942=>x"8b00", 943=>x"8c00", 944=>x"9200",
---- 945=>x"8d00", 946=>x"8b00", 947=>x"8d00", 948=>x"8e00",
---- 949=>x"8d00", 950=>x"7400", 951=>x"8c00", 952=>x"8e00",
---- 953=>x"8e00", 954=>x"8e00", 955=>x"7300", 956=>x"8e00",
---- 957=>x"9000", 958=>x"8e00", 959=>x"8b00", 960=>x"9000",
---- 961=>x"9000", 962=>x"8c00", 963=>x"8c00", 964=>x"8f00",
---- 965=>x"9200", 966=>x"8d00", 967=>x"8d00", 968=>x"8d00",
---- 969=>x"9000", 970=>x"9000", 971=>x"8e00", 972=>x"8f00",
---- 973=>x"9100", 974=>x"9100", 975=>x"8f00", 976=>x"9100",
---- 977=>x"9300", 978=>x"6d00", 979=>x"9100", 980=>x"9200",
---- 981=>x"9100", 982=>x"9000", 983=>x"9400", 984=>x"8f00",
---- 985=>x"9100", 986=>x"9100", 987=>x"9200", 988=>x"9100",
---- 989=>x"9300", 990=>x"9200", 991=>x"9500", 992=>x"9100",
---- 993=>x"6d00", 994=>x"9100", 995=>x"9200", 996=>x"8e00",
---- 997=>x"9200", 998=>x"9000", 999=>x"9100", 1000=>x"8f00",
---- 1001=>x"9100", 1002=>x"9200", 1003=>x"6e00", 1004=>x"8f00",
---- 1005=>x"9200", 1006=>x"8e00", 1007=>x"8f00", 1008=>x"8f00",
---- 1009=>x"9000", 1010=>x"8f00", 1011=>x"9200", 1012=>x"8f00",
---- 1013=>x"9100", 1014=>x"9000", 1015=>x"9400", 1016=>x"9100",
---- 1017=>x"9000", 1018=>x"9200", 1019=>x"9100", 1020=>x"8f00",
---- 1021=>x"9100", 1022=>x"9100", 1023=>x"8f00"),
----
---- 35 => (0=>x"8200", 1=>x"7f00", 2=>x"8200", 3=>x"8300", 4=>x"8200",
---- 5=>x"7f00", 6=>x"8200", 7=>x"8300", 8=>x"8100",
---- 9=>x"7e00", 10=>x"8100", 11=>x"8200", 12=>x"7e00",
---- 13=>x"7e00", 14=>x"8100", 15=>x"8300", 16=>x"7d00",
---- 17=>x"7e00", 18=>x"7f00", 19=>x"7f00", 20=>x"7f00",
---- 21=>x"8000", 22=>x"7e00", 23=>x"7f00", 24=>x"7f00",
---- 25=>x"8100", 26=>x"8000", 27=>x"8200", 28=>x"8000",
---- 29=>x"7f00", 30=>x"7f00", 31=>x"8100", 32=>x"7f00",
---- 33=>x"7b00", 34=>x"8000", 35=>x"8100", 36=>x"8100",
---- 37=>x"7e00", 38=>x"7f00", 39=>x"7e00", 40=>x"8300",
---- 41=>x"7e00", 42=>x"7d00", 43=>x"7f00", 44=>x"7d00",
---- 45=>x"7f00", 46=>x"7d00", 47=>x"8000", 48=>x"7e00",
---- 49=>x"7d00", 50=>x"7c00", 51=>x"7e00", 52=>x"8000",
---- 53=>x"7e00", 54=>x"7e00", 55=>x"7f00", 56=>x"7d00",
---- 57=>x"7f00", 58=>x"7f00", 59=>x"7d00", 60=>x"8100",
---- 61=>x"7e00", 62=>x"7c00", 63=>x"7f00", 64=>x"8000",
---- 65=>x"7e00", 66=>x"7c00", 67=>x"7f00", 68=>x"8100",
---- 69=>x"7d00", 70=>x"7d00", 71=>x"7e00", 72=>x"7e00",
---- 73=>x"7e00", 74=>x"7c00", 75=>x"7d00", 76=>x"7e00",
---- 77=>x"8000", 78=>x"7e00", 79=>x"7d00", 80=>x"7e00",
---- 81=>x"7d00", 82=>x"7e00", 83=>x"7f00", 84=>x"7f00",
---- 85=>x"7c00", 86=>x"8200", 87=>x"8200", 88=>x"8200",
---- 89=>x"7e00", 90=>x"8000", 91=>x"8000", 92=>x"8300",
---- 93=>x"7f00", 94=>x"8000", 95=>x"7d00", 96=>x"8300",
---- 97=>x"8300", 98=>x"8200", 99=>x"7d00", 100=>x"8100",
---- 101=>x"8100", 102=>x"8000", 103=>x"7d00", 104=>x"7d00",
---- 105=>x"7f00", 106=>x"7f00", 107=>x"7e00", 108=>x"7d00",
---- 109=>x"7f00", 110=>x"7f00", 111=>x"8100", 112=>x"7e00",
---- 113=>x"8100", 114=>x"7f00", 115=>x"7e00", 116=>x"7a00",
---- 117=>x"7d00", 118=>x"8000", 119=>x"7b00", 120=>x"7600",
---- 121=>x"7500", 122=>x"7700", 123=>x"7900", 124=>x"7100",
---- 125=>x"7100", 126=>x"7600", 127=>x"7800", 128=>x"6a00",
---- 129=>x"6d00", 130=>x"7200", 131=>x"7200", 132=>x"8500",
---- 133=>x"9700", 134=>x"6700", 135=>x"6b00", 136=>x"c300",
---- 137=>x"9e00", 138=>x"6c00", 139=>x"6300", 140=>x"cc00",
---- 141=>x"ca00", 142=>x"ab00", 143=>x"7200", 144=>x"ca00",
---- 145=>x"ca00", 146=>x"d000", 147=>x"b100", 148=>x"c400",
---- 149=>x"c100", 150=>x"c400", 151=>x"cc00", 152=>x"bc00",
---- 153=>x"c100", 154=>x"cb00", 155=>x"d500", 156=>x"d300",
---- 157=>x"d700", 158=>x"d900", 159=>x"db00", 160=>x"d800",
---- 161=>x"d600", 162=>x"d500", 163=>x"d700", 164=>x"d200",
---- 165=>x"d600", 166=>x"d200", 167=>x"d300", 168=>x"d000",
---- 169=>x"d200", 170=>x"d300", 171=>x"ce00", 172=>x"cf00",
---- 173=>x"cd00", 174=>x"d200", 175=>x"d500", 176=>x"3200",
---- 177=>x"cf00", 178=>x"cf00", 179=>x"d200", 180=>x"ce00",
---- 181=>x"cb00", 182=>x"cf00", 183=>x"3200", 184=>x"cc00",
---- 185=>x"ca00", 186=>x"ca00", 187=>x"cf00", 188=>x"ca00",
---- 189=>x"ce00", 190=>x"d600", 191=>x"d900", 192=>x"d100",
---- 193=>x"cb00", 194=>x"cf00", 195=>x"ce00", 196=>x"c800",
---- 197=>x"c500", 198=>x"c700", 199=>x"c800", 200=>x"c900",
---- 201=>x"cb00", 202=>x"d000", 203=>x"cd00", 204=>x"cf00",
---- 205=>x"ce00", 206=>x"cd00", 207=>x"cf00", 208=>x"d200",
---- 209=>x"cf00", 210=>x"cf00", 211=>x"cf00", 212=>x"ce00",
---- 213=>x"cd00", 214=>x"d000", 215=>x"cc00", 216=>x"c300",
---- 217=>x"cf00", 218=>x"d000", 219=>x"cf00", 220=>x"c800",
---- 221=>x"cc00", 222=>x"cd00", 223=>x"cc00", 224=>x"ce00",
---- 225=>x"ca00", 226=>x"cd00", 227=>x"cf00", 228=>x"ca00",
---- 229=>x"cc00", 230=>x"c700", 231=>x"c600", 232=>x"c400",
---- 233=>x"c100", 234=>x"ca00", 235=>x"cb00", 236=>x"c400",
---- 237=>x"c800", 238=>x"ce00", 239=>x"cf00", 240=>x"cc00",
---- 241=>x"ca00", 242=>x"ca00", 243=>x"cd00", 244=>x"cc00",
---- 245=>x"c800", 246=>x"ca00", 247=>x"cc00", 248=>x"c500",
---- 249=>x"3900", 250=>x"cb00", 251=>x"cb00", 252=>x"c000",
---- 253=>x"bb00", 254=>x"c400", 255=>x"cb00", 256=>x"c800",
---- 257=>x"c100", 258=>x"bc00", 259=>x"c700", 260=>x"c500",
---- 261=>x"c700", 262=>x"c300", 263=>x"c000", 264=>x"c300",
---- 265=>x"c300", 266=>x"c400", 267=>x"c900", 268=>x"c500",
---- 269=>x"c900", 270=>x"c500", 271=>x"c600", 272=>x"c000",
---- 273=>x"ca00", 274=>x"c800", 275=>x"c600", 276=>x"be00",
---- 277=>x"c700", 278=>x"3200", 279=>x"cd00", 280=>x"c300",
---- 281=>x"be00", 282=>x"c400", 283=>x"be00", 284=>x"b200",
---- 285=>x"a200", 286=>x"ab00", 287=>x"ad00", 288=>x"a100",
---- 289=>x"ae00", 290=>x"ba00", 291=>x"b800", 292=>x"b300",
---- 293=>x"b400", 294=>x"b600", 295=>x"b900", 296=>x"b700",
---- 297=>x"b600", 298=>x"b900", 299=>x"b300", 300=>x"b200",
---- 301=>x"b400", 302=>x"b800", 303=>x"ad00", 304=>x"b000",
---- 305=>x"b200", 306=>x"b800", 307=>x"b700", 308=>x"af00",
---- 309=>x"b200", 310=>x"b700", 311=>x"bc00", 312=>x"b000",
---- 313=>x"b200", 314=>x"b000", 315=>x"ba00", 316=>x"ac00",
---- 317=>x"af00", 318=>x"ae00", 319=>x"ae00", 320=>x"b000",
---- 321=>x"ad00", 322=>x"a700", 323=>x"a900", 324=>x"b100",
---- 325=>x"a900", 326=>x"a300", 327=>x"ab00", 328=>x"ac00",
---- 329=>x"ab00", 330=>x"a400", 331=>x"a400", 332=>x"a600",
---- 333=>x"a600", 334=>x"a600", 335=>x"a800", 336=>x"a700",
---- 337=>x"a200", 338=>x"a600", 339=>x"a600", 340=>x"9e00",
---- 341=>x"a300", 342=>x"a100", 343=>x"a500", 344=>x"9600",
---- 345=>x"8f00", 346=>x"8700", 347=>x"6700", 348=>x"a600",
---- 349=>x"7a00", 350=>x"7a00", 351=>x"5000", 352=>x"6700",
---- 353=>x"4f00", 354=>x"6700", 355=>x"7500", 356=>x"2900",
---- 357=>x"3400", 358=>x"2c00", 359=>x"3c00", 360=>x"2b00",
---- 361=>x"2f00", 362=>x"2d00", 363=>x"2200", 364=>x"2d00",
---- 365=>x"3700", 366=>x"2600", 367=>x"4f00", 368=>x"2300",
---- 369=>x"1e00", 370=>x"3300", 371=>x"9600", 372=>x"1d00",
---- 373=>x"4000", 374=>x"9100", 375=>x"ba00", 376=>x"5600",
---- 377=>x"a600", 378=>x"b900", 379=>x"8400", 380=>x"ac00",
---- 381=>x"b000", 382=>x"8100", 383=>x"7400", 384=>x"a400",
---- 385=>x"7b00", 386=>x"8300", 387=>x"ad00", 388=>x"7600",
---- 389=>x"8700", 390=>x"b500", 391=>x"c700", 392=>x"8e00",
---- 393=>x"b100", 394=>x"c400", 395=>x"c700", 396=>x"bd00",
---- 397=>x"be00", 398=>x"c300", 399=>x"c700", 400=>x"c800",
---- 401=>x"c200", 402=>x"c000", 403=>x"c100", 404=>x"c600",
---- 405=>x"c200", 406=>x"bf00", 407=>x"be00", 408=>x"c200",
---- 409=>x"c100", 410=>x"be00", 411=>x"bb00", 412=>x"c100",
---- 413=>x"c100", 414=>x"b900", 415=>x"b800", 416=>x"bf00",
---- 417=>x"bc00", 418=>x"ba00", 419=>x"b700", 420=>x"bb00",
---- 421=>x"b800", 422=>x"b500", 423=>x"af00", 424=>x"b600",
---- 425=>x"b300", 426=>x"ac00", 427=>x"ab00", 428=>x"b300",
---- 429=>x"ad00", 430=>x"ab00", 431=>x"a800", 432=>x"b300",
---- 433=>x"aa00", 434=>x"a300", 435=>x"a500", 436=>x"ac00",
---- 437=>x"a300", 438=>x"5f00", 439=>x"a500", 440=>x"5900",
---- 441=>x"a200", 442=>x"9e00", 443=>x"a300", 444=>x"a400",
---- 445=>x"a200", 446=>x"a000", 447=>x"a100", 448=>x"a800",
---- 449=>x"a500", 450=>x"a400", 451=>x"a700", 452=>x"aa00",
---- 453=>x"ab00", 454=>x"aa00", 455=>x"ae00", 456=>x"ab00",
---- 457=>x"aa00", 458=>x"a900", 459=>x"9e00", 460=>x"a600",
---- 461=>x"a300", 462=>x"9b00", 463=>x"9400", 464=>x"a500",
---- 465=>x"9b00", 466=>x"9700", 467=>x"9e00", 468=>x"9c00",
---- 469=>x"9b00", 470=>x"a100", 471=>x"a100", 472=>x"9a00",
---- 473=>x"9d00", 474=>x"a200", 475=>x"a200", 476=>x"a200",
---- 477=>x"9f00", 478=>x"a300", 479=>x"a500", 480=>x"a400",
---- 481=>x"a300", 482=>x"a500", 483=>x"a700", 484=>x"a600",
---- 485=>x"a600", 486=>x"aa00", 487=>x"aa00", 488=>x"9800",
---- 489=>x"9d00", 490=>x"a700", 491=>x"ac00", 492=>x"7400",
---- 493=>x"8000", 494=>x"9100", 495=>x"a200", 496=>x"4300",
---- 497=>x"4c00", 498=>x"5b00", 499=>x"7100", 500=>x"4e00",
---- 501=>x"4700", 502=>x"4000", 503=>x"4000", 504=>x"6900",
---- 505=>x"5f00", 506=>x"5800", 507=>x"4d00", 508=>x"6100",
---- 509=>x"7500", 510=>x"6d00", 511=>x"6600", 512=>x"5200",
---- 513=>x"7d00", 514=>x"6700", 515=>x"7600", 516=>x"2d00",
---- 517=>x"4500", 518=>x"6a00", 519=>x"8e00", 520=>x"2b00",
---- 521=>x"2700", 522=>x"3f00", 523=>x"7200", 524=>x"2700",
---- 525=>x"2900", 526=>x"2300", 527=>x"4000", 528=>x"4300",
---- 529=>x"2b00", 530=>x"4800", 531=>x"4200", 532=>x"8d00",
---- 533=>x"4600", 534=>x"6400", 535=>x"6c00", 536=>x"b800",
---- 537=>x"6900", 538=>x"4f00", 539=>x"7700", 540=>x"b200",
---- 541=>x"8500", 542=>x"6300", 543=>x"7600", 544=>x"6b00",
---- 545=>x"8e00", 546=>x"8600", 547=>x"6f00", 548=>x"9e00",
---- 549=>x"9100", 550=>x"8500", 551=>x"7a00", 552=>x"b100",
---- 553=>x"ad00", 554=>x"a600", 555=>x"9200", 556=>x"9b00",
---- 557=>x"a700", 558=>x"9e00", 559=>x"8b00", 560=>x"9700",
---- 561=>x"9300", 562=>x"9200", 563=>x"9300", 564=>x"a200",
---- 565=>x"9b00", 566=>x"a400", 567=>x"9800", 568=>x"a300",
---- 569=>x"a500", 570=>x"a500", 571=>x"9000", 572=>x"a700",
---- 573=>x"a800", 574=>x"9e00", 575=>x"8d00", 576=>x"a800",
---- 577=>x"a100", 578=>x"9a00", 579=>x"8e00", 580=>x"a800",
---- 581=>x"9d00", 582=>x"9800", 583=>x"9400", 584=>x"a800",
---- 585=>x"a300", 586=>x"9900", 587=>x"9200", 588=>x"a500",
---- 589=>x"a000", 590=>x"9b00", 591=>x"9600", 592=>x"a400",
---- 593=>x"9f00", 594=>x"9900", 595=>x"9600", 596=>x"a000",
---- 597=>x"9d00", 598=>x"9900", 599=>x"9300", 600=>x"a000",
---- 601=>x"9b00", 602=>x"9100", 603=>x"8e00", 604=>x"9f00",
---- 605=>x"9a00", 606=>x"9200", 607=>x"8f00", 608=>x"9d00",
---- 609=>x"9600", 610=>x"9200", 611=>x"8800", 612=>x"9b00",
---- 613=>x"9800", 614=>x"8e00", 615=>x"8500", 616=>x"9b00",
---- 617=>x"9700", 618=>x"8c00", 619=>x"8600", 620=>x"9b00",
---- 621=>x"9400", 622=>x"8c00", 623=>x"8600", 624=>x"9700",
---- 625=>x"9000", 626=>x"8900", 627=>x"8100", 628=>x"9400",
---- 629=>x"9000", 630=>x"8900", 631=>x"7b00", 632=>x"9200",
---- 633=>x"8f00", 634=>x"8100", 635=>x"7100", 636=>x"6e00",
---- 637=>x"8f00", 638=>x"7f00", 639=>x"6b00", 640=>x"9200",
---- 641=>x"9100", 642=>x"8100", 643=>x"6c00", 644=>x"9200",
---- 645=>x"8e00", 646=>x"8500", 647=>x"7500", 648=>x"9500",
---- 649=>x"9300", 650=>x"8b00", 651=>x"7a00", 652=>x"9500",
---- 653=>x"9400", 654=>x"9200", 655=>x"8400", 656=>x"9800",
---- 657=>x"9500", 658=>x"9400", 659=>x"8e00", 660=>x"9b00",
---- 661=>x"9a00", 662=>x"9700", 663=>x"9400", 664=>x"9b00",
---- 665=>x"9e00", 666=>x"9900", 667=>x"9500", 668=>x"9a00",
---- 669=>x"9600", 670=>x"9900", 671=>x"9600", 672=>x"9900",
---- 673=>x"9500", 674=>x"9600", 675=>x"9700", 676=>x"9a00",
---- 677=>x"9200", 678=>x"9100", 679=>x"9600", 680=>x"9600",
---- 681=>x"9600", 682=>x"9200", 683=>x"9300", 684=>x"9100",
---- 685=>x"9100", 686=>x"9200", 687=>x"9200", 688=>x"9100",
---- 689=>x"8f00", 690=>x"8f00", 691=>x"7000", 692=>x"8e00",
---- 693=>x"8f00", 694=>x"8f00", 695=>x"9000", 696=>x"8600",
---- 697=>x"8400", 698=>x"8300", 699=>x"7f00", 700=>x"9500",
---- 701=>x"6900", 702=>x"7000", 703=>x"6a00", 704=>x"6600",
---- 705=>x"6b00", 706=>x"7300", 707=>x"7000", 708=>x"7900",
---- 709=>x"7d00", 710=>x"8400", 711=>x"8700", 712=>x"7900",
---- 713=>x"7900", 714=>x"7f00", 715=>x"8600", 716=>x"8000",
---- 717=>x"7f00", 718=>x"7f00", 719=>x"7e00", 720=>x"7b00",
---- 721=>x"8100", 722=>x"8300", 723=>x"8000", 724=>x"7e00",
---- 725=>x"7c00", 726=>x"7b00", 727=>x"7c00", 728=>x"8500",
---- 729=>x"8000", 730=>x"7c00", 731=>x"7700", 732=>x"8400",
---- 733=>x"8000", 734=>x"8200", 735=>x"8300", 736=>x"8700",
---- 737=>x"8500", 738=>x"8900", 739=>x"8e00", 740=>x"8e00",
---- 741=>x"8d00", 742=>x"9500", 743=>x"9900", 744=>x"9700",
---- 745=>x"9300", 746=>x"9500", 747=>x"9b00", 748=>x"9f00",
---- 749=>x"9c00", 750=>x"9900", 751=>x"a000", 752=>x"a600",
---- 753=>x"a700", 754=>x"a300", 755=>x"a200", 756=>x"5900",
---- 757=>x"ac00", 758=>x"a800", 759=>x"a600", 760=>x"9e00",
---- 761=>x"a700", 762=>x"a400", 763=>x"a700", 764=>x"9c00",
---- 765=>x"9c00", 766=>x"a200", 767=>x"a800", 768=>x"9900",
---- 769=>x"6b00", 770=>x"9900", 771=>x"a300", 772=>x"9600",
---- 773=>x"9400", 774=>x"9700", 775=>x"9d00", 776=>x"9e00",
---- 777=>x"a100", 778=>x"a000", 779=>x"a000", 780=>x"9b00",
---- 781=>x"9e00", 782=>x"9a00", 783=>x"9900", 784=>x"9400",
---- 785=>x"9900", 786=>x"9700", 787=>x"9600", 788=>x"9500",
---- 789=>x"9300", 790=>x"9200", 791=>x"9100", 792=>x"9100",
---- 793=>x"8d00", 794=>x"8f00", 795=>x"8d00", 796=>x"8c00",
---- 797=>x"8c00", 798=>x"8d00", 799=>x"8c00", 800=>x"8e00",
---- 801=>x"8d00", 802=>x"8900", 803=>x"8d00", 804=>x"8d00",
---- 805=>x"8a00", 806=>x"8a00", 807=>x"9000", 808=>x"8c00",
---- 809=>x"8900", 810=>x"8b00", 811=>x"9100", 812=>x"8700",
---- 813=>x"8700", 814=>x"8b00", 815=>x"9100", 816=>x"8800",
---- 817=>x"8a00", 818=>x"8c00", 819=>x"9000", 820=>x"8a00",
---- 821=>x"8d00", 822=>x"8e00", 823=>x"9300", 824=>x"8a00",
---- 825=>x"8f00", 826=>x"9400", 827=>x"9600", 828=>x"8c00",
---- 829=>x"8f00", 830=>x"6a00", 831=>x"9600", 832=>x"9100",
---- 833=>x"8f00", 834=>x"9200", 835=>x"9500", 836=>x"8f00",
---- 837=>x"9100", 838=>x"9100", 839=>x"9400", 840=>x"8e00",
---- 841=>x"8f00", 842=>x"9200", 843=>x"9700", 844=>x"8d00",
---- 845=>x"9000", 846=>x"9200", 847=>x"9600", 848=>x"9100",
---- 849=>x"9400", 850=>x"9500", 851=>x"9700", 852=>x"9100",
---- 853=>x"9500", 854=>x"9400", 855=>x"9100", 856=>x"8f00",
---- 857=>x"8f00", 858=>x"9400", 859=>x"9000", 860=>x"8d00",
---- 861=>x"9100", 862=>x"9200", 863=>x"8f00", 864=>x"8f00",
---- 865=>x"9100", 866=>x"9100", 867=>x"9300", 868=>x"9000",
---- 869=>x"9000", 870=>x"9200", 871=>x"9000", 872=>x"8d00",
---- 873=>x"8d00", 874=>x"9000", 875=>x"9000", 876=>x"8e00",
---- 877=>x"8f00", 878=>x"9000", 879=>x"9000", 880=>x"8c00",
---- 881=>x"8c00", 882=>x"8d00", 883=>x"8d00", 884=>x"8a00",
---- 885=>x"8c00", 886=>x"8d00", 887=>x"8f00", 888=>x"8b00",
---- 889=>x"8a00", 890=>x"8e00", 891=>x"9000", 892=>x"8a00",
---- 893=>x"8800", 894=>x"8c00", 895=>x"8f00", 896=>x"8a00",
---- 897=>x"8b00", 898=>x"8c00", 899=>x"8c00", 900=>x"8a00",
---- 901=>x"8c00", 902=>x"8a00", 903=>x"8b00", 904=>x"8c00",
---- 905=>x"8b00", 906=>x"8800", 907=>x"8c00", 908=>x"8700",
---- 909=>x"8800", 910=>x"8800", 911=>x"8a00", 912=>x"8700",
---- 913=>x"8900", 914=>x"8500", 915=>x"8b00", 916=>x"8a00",
---- 917=>x"8c00", 918=>x"8900", 919=>x"8c00", 920=>x"8900",
---- 921=>x"8b00", 922=>x"8b00", 923=>x"8c00", 924=>x"8b00",
---- 925=>x"8700", 926=>x"8700", 927=>x"8800", 928=>x"8a00",
---- 929=>x"8700", 930=>x"8800", 931=>x"8900", 932=>x"8a00",
---- 933=>x"8700", 934=>x"8800", 935=>x"8600", 936=>x"8a00",
---- 937=>x"8600", 938=>x"8500", 939=>x"8800", 940=>x"8900",
---- 941=>x"8800", 942=>x"8700", 943=>x"8800", 944=>x"8900",
---- 945=>x"8900", 946=>x"8a00", 947=>x"8700", 948=>x"8900",
---- 949=>x"8800", 950=>x"8a00", 951=>x"8600", 952=>x"8a00",
---- 953=>x"7500", 954=>x"8a00", 955=>x"8b00", 956=>x"8a00",
---- 957=>x"8c00", 958=>x"8b00", 959=>x"8a00", 960=>x"8d00",
---- 961=>x"8b00", 962=>x"8a00", 963=>x"8900", 964=>x"8f00",
---- 965=>x"8e00", 966=>x"7400", 967=>x"8a00", 968=>x"8c00",
---- 969=>x"8d00", 970=>x"8e00", 971=>x"8a00", 972=>x"8f00",
---- 973=>x"8e00", 974=>x"8f00", 975=>x"8d00", 976=>x"9100",
---- 977=>x"8f00", 978=>x"9100", 979=>x"8e00", 980=>x"9100",
---- 981=>x"9100", 982=>x"8e00", 983=>x"8d00", 984=>x"9100",
---- 985=>x"9100", 986=>x"8f00", 987=>x"8d00", 988=>x"9100",
---- 989=>x"9000", 990=>x"9200", 991=>x"8f00", 992=>x"9000",
---- 993=>x"8d00", 994=>x"9300", 995=>x"9000", 996=>x"9100",
---- 997=>x"9100", 998=>x"9200", 999=>x"9300", 1000=>x"9100",
---- 1001=>x"9000", 1002=>x"9400", 1003=>x"9200", 1004=>x"9500",
---- 1005=>x"9300", 1006=>x"9400", 1007=>x"9400", 1008=>x"9000",
---- 1009=>x"9000", 1010=>x"9500", 1011=>x"9300", 1012=>x"9200",
---- 1013=>x"9300", 1014=>x"8f00", 1015=>x"9000", 1016=>x"9200",
---- 1017=>x"9400", 1018=>x"8c00", 1019=>x"9100", 1020=>x"8f00",
---- 1021=>x"9000", 1022=>x"8e00", 1023=>x"9100"),
----
---- 36 => (0=>x"8000", 1=>x"8200", 2=>x"8100", 3=>x"8100", 4=>x"8000",
---- 5=>x"8300", 6=>x"8000", 7=>x"8000", 8=>x"7f00",
---- 9=>x"8100", 10=>x"8200", 11=>x"8000", 12=>x"7f00",
---- 13=>x"8100", 14=>x"8200", 15=>x"7f00", 16=>x"8000",
---- 17=>x"8300", 18=>x"7f00", 19=>x"7f00", 20=>x"7d00",
---- 21=>x"8000", 22=>x"8200", 23=>x"7f00", 24=>x"7f00",
---- 25=>x"7c00", 26=>x"8000", 27=>x"8100", 28=>x"7f00",
---- 29=>x"7e00", 30=>x"8000", 31=>x"8300", 32=>x"8100",
---- 33=>x"8200", 34=>x"8000", 35=>x"8100", 36=>x"8000",
---- 37=>x"8200", 38=>x"8300", 39=>x"8100", 40=>x"7f00",
---- 41=>x"7e00", 42=>x"8300", 43=>x"8200", 44=>x"7f00",
---- 45=>x"7c00", 46=>x"7f00", 47=>x"7f00", 48=>x"7e00",
---- 49=>x"8000", 50=>x"7f00", 51=>x"7d00", 52=>x"7f00",
---- 53=>x"7f00", 54=>x"7f00", 55=>x"7e00", 56=>x"7d00",
---- 57=>x"7e00", 58=>x"7e00", 59=>x"7e00", 60=>x"7c00",
---- 61=>x"7d00", 62=>x"7c00", 63=>x"7f00", 64=>x"7f00",
---- 65=>x"7d00", 66=>x"7e00", 67=>x"7e00", 68=>x"8000",
---- 69=>x"7f00", 70=>x"7b00", 71=>x"7d00", 72=>x"7a00",
---- 73=>x"7f00", 74=>x"7f00", 75=>x"7d00", 76=>x"7d00",
---- 77=>x"7c00", 78=>x"7e00", 79=>x"7d00", 80=>x"8000",
---- 81=>x"7e00", 82=>x"7d00", 83=>x"7f00", 84=>x"7c00",
---- 85=>x"7f00", 86=>x"7d00", 87=>x"7e00", 88=>x"7e00",
---- 89=>x"8000", 90=>x"8200", 91=>x"7f00", 92=>x"7d00",
---- 93=>x"7e00", 94=>x"8100", 95=>x"7e00", 96=>x"8000",
---- 97=>x"7d00", 98=>x"7e00", 99=>x"7f00", 100=>x"8000",
---- 101=>x"7e00", 102=>x"7c00", 103=>x"8100", 104=>x"7e00",
---- 105=>x"8000", 106=>x"7d00", 107=>x"8000", 108=>x"7e00",
---- 109=>x"7e00", 110=>x"7a00", 111=>x"7e00", 112=>x"7e00",
---- 113=>x"7b00", 114=>x"7d00", 115=>x"8000", 116=>x"7800",
---- 117=>x"7900", 118=>x"7e00", 119=>x"7d00", 120=>x"7900",
---- 121=>x"7900", 122=>x"7700", 123=>x"7a00", 124=>x"7700",
---- 125=>x"7600", 126=>x"7a00", 127=>x"7900", 128=>x"7400",
---- 129=>x"7700", 130=>x"7800", 131=>x"7800", 132=>x"6e00",
---- 133=>x"7500", 134=>x"7400", 135=>x"7100", 136=>x"6c00",
---- 137=>x"6c00", 138=>x"6a00", 139=>x"6c00", 140=>x"6200",
---- 141=>x"6500", 142=>x"6800", 143=>x"6900", 144=>x"7500",
---- 145=>x"5900", 146=>x"5d00", 147=>x"6000", 148=>x"bb00",
---- 149=>x"7b00", 150=>x"7200", 151=>x"6400", 152=>x"da00",
---- 153=>x"d500", 154=>x"cf00", 155=>x"b900", 156=>x"dc00",
---- 157=>x"e400", 158=>x"e600", 159=>x"e900", 160=>x"d600",
---- 161=>x"da00", 162=>x"e100", 163=>x"e300", 164=>x"d800",
---- 165=>x"d700", 166=>x"dd00", 167=>x"e200", 168=>x"d000",
---- 169=>x"d600", 170=>x"d800", 171=>x"df00", 172=>x"cd00",
---- 173=>x"d000", 174=>x"d800", 175=>x"da00", 176=>x"d300",
---- 177=>x"ce00", 178=>x"d000", 179=>x"d400", 180=>x"cd00",
---- 181=>x"d200", 182=>x"d200", 183=>x"d600", 184=>x"d100",
---- 185=>x"d400", 186=>x"2600", 187=>x"d900", 188=>x"d700",
---- 189=>x"d200", 190=>x"d500", 191=>x"d200", 192=>x"cb00",
---- 193=>x"ca00", 194=>x"cc00", 195=>x"ce00", 196=>x"c700",
---- 197=>x"ce00", 198=>x"d100", 199=>x"d100", 200=>x"ce00",
---- 201=>x"cf00", 202=>x"d100", 203=>x"d300", 204=>x"d000",
---- 205=>x"d000", 206=>x"ce00", 207=>x"d200", 208=>x"cf00",
---- 209=>x"d000", 210=>x"cd00", 211=>x"cb00", 212=>x"ce00",
---- 213=>x"d100", 214=>x"cf00", 215=>x"ce00", 216=>x"ce00",
---- 217=>x"d200", 218=>x"cf00", 219=>x"cf00", 220=>x"cd00",
---- 221=>x"cb00", 222=>x"cc00", 223=>x"cb00", 224=>x"cb00",
---- 225=>x"c300", 226=>x"c400", 227=>x"c900", 228=>x"c800",
---- 229=>x"cb00", 230=>x"c800", 231=>x"cb00", 232=>x"cb00",
---- 233=>x"d400", 234=>x"cd00", 235=>x"c400", 236=>x"cc00",
---- 237=>x"ca00", 238=>x"d200", 239=>x"cd00", 240=>x"ce00",
---- 241=>x"c900", 242=>x"c900", 243=>x"cd00", 244=>x"cb00",
---- 245=>x"c800", 246=>x"c600", 247=>x"c300", 248=>x"c500",
---- 249=>x"c600", 250=>x"ca00", 251=>x"c700", 252=>x"ca00",
---- 253=>x"c600", 254=>x"c800", 255=>x"3400", 256=>x"cb00",
---- 257=>x"c900", 258=>x"c600", 259=>x"c800", 260=>x"c600",
---- 261=>x"cc00", 262=>x"c900", 263=>x"c300", 264=>x"c000",
---- 265=>x"c900", 266=>x"cc00", 267=>x"c900", 268=>x"c700",
---- 269=>x"c600", 270=>x"cb00", 271=>x"bc00", 272=>x"ca00",
---- 273=>x"ca00", 274=>x"af00", 275=>x"9900", 276=>x"c400",
---- 277=>x"b100", 278=>x"a800", 279=>x"b100", 280=>x"aa00",
---- 281=>x"ab00", 282=>x"c000", 283=>x"c300", 284=>x"b200",
---- 285=>x"bf00", 286=>x"bb00", 287=>x"b600", 288=>x"bc00",
---- 289=>x"bc00", 290=>x"af00", 291=>x"ab00", 292=>x"c100",
---- 293=>x"bd00", 294=>x"bb00", 295=>x"b600", 296=>x"b500",
---- 297=>x"bc00", 298=>x"bd00", 299=>x"c000", 300=>x"b200",
---- 301=>x"b900", 302=>x"4600", 303=>x"c100", 304=>x"af00",
---- 305=>x"b500", 306=>x"b900", 307=>x"bd00", 308=>x"b600",
---- 309=>x"ae00", 310=>x"b700", 311=>x"be00", 312=>x"bc00",
---- 313=>x"b700", 314=>x"b000", 315=>x"b500", 316=>x"ba00",
---- 317=>x"bb00", 318=>x"b400", 319=>x"ae00", 320=>x"af00",
---- 321=>x"ba00", 322=>x"b400", 323=>x"af00", 324=>x"a700",
---- 325=>x"ac00", 326=>x"b200", 327=>x"ac00", 328=>x"a900",
---- 329=>x"a300", 330=>x"a100", 331=>x"a400", 332=>x"9f00",
---- 333=>x"a400", 334=>x"a000", 335=>x"a000", 336=>x"a600",
---- 337=>x"9a00", 338=>x"a300", 339=>x"a900", 340=>x"a500",
---- 341=>x"a200", 342=>x"9e00", 343=>x"a100", 344=>x"9800",
---- 345=>x"a400", 346=>x"9e00", 347=>x"9100", 348=>x"3f00",
---- 349=>x"7f00", 350=>x"a100", 351=>x"9100", 352=>x"2d00",
---- 353=>x"3e00", 354=>x"9a00", 355=>x"9600", 356=>x"2900",
---- 357=>x"2600", 358=>x"7b00", 359=>x"bc00", 360=>x"2400",
---- 361=>x"5200", 362=>x"a800", 363=>x"bf00", 364=>x"7000",
---- 365=>x"b200", 366=>x"b400", 367=>x"8b00", 368=>x"be00",
---- 369=>x"a100", 370=>x"8900", 371=>x"9800", 372=>x"9200",
---- 373=>x"7300", 374=>x"9e00", 375=>x"c400", 376=>x"6b00",
---- 377=>x"9800", 378=>x"c300", 379=>x"c700", 380=>x"a100",
---- 381=>x"bb00", 382=>x"c200", 383=>x"be00", 384=>x"c700",
---- 385=>x"be00", 386=>x"bf00", 387=>x"b700", 388=>x"c300",
---- 389=>x"bc00", 390=>x"ba00", 391=>x"b700", 392=>x"be00",
---- 393=>x"b600", 394=>x"b700", 395=>x"b200", 396=>x"bb00",
---- 397=>x"b400", 398=>x"b000", 399=>x"b300", 400=>x"bc00",
---- 401=>x"b500", 402=>x"b300", 403=>x"b300", 404=>x"bd00",
---- 405=>x"b900", 406=>x"b600", 407=>x"b700", 408=>x"ba00",
---- 409=>x"b500", 410=>x"4a00", 411=>x"b100", 412=>x"b600",
---- 413=>x"b300", 414=>x"b200", 415=>x"b200", 416=>x"b400",
---- 417=>x"b200", 418=>x"b400", 419=>x"b100", 420=>x"ad00",
---- 421=>x"af00", 422=>x"b200", 423=>x"af00", 424=>x"a500",
---- 425=>x"ad00", 426=>x"b000", 427=>x"ab00", 428=>x"a900",
---- 429=>x"b100", 430=>x"ae00", 431=>x"b000", 432=>x"aa00",
---- 433=>x"ac00", 434=>x"b200", 435=>x"b300", 436=>x"a600",
---- 437=>x"a900", 438=>x"b300", 439=>x"b500", 440=>x"a900",
---- 441=>x"b000", 442=>x"b700", 443=>x"b300", 444=>x"ad00",
---- 445=>x"b900", 446=>x"b400", 447=>x"a100", 448=>x"b500",
---- 449=>x"ae00", 450=>x"9500", 451=>x"9e00", 452=>x"a600",
---- 453=>x"9400", 454=>x"9a00", 455=>x"a400", 456=>x"9400",
---- 457=>x"9700", 458=>x"a400", 459=>x"a800", 460=>x"9e00",
---- 461=>x"9f00", 462=>x"a400", 463=>x"ab00", 464=>x"9f00",
---- 465=>x"a600", 466=>x"a800", 467=>x"ac00", 468=>x"a500",
---- 469=>x"ab00", 470=>x"ac00", 471=>x"ad00", 472=>x"a800",
---- 473=>x"ad00", 474=>x"ab00", 475=>x"ae00", 476=>x"aa00",
---- 477=>x"ae00", 478=>x"ac00", 479=>x"ae00", 480=>x"ab00",
---- 481=>x"b000", 482=>x"b000", 483=>x"af00", 484=>x"af00",
---- 485=>x"af00", 486=>x"b200", 487=>x"b200", 488=>x"af00",
---- 489=>x"b100", 490=>x"b300", 491=>x"b500", 492=>x"ab00",
---- 493=>x"b200", 494=>x"b600", 495=>x"b500", 496=>x"8d00",
---- 497=>x"a600", 498=>x"b100", 499=>x"b200", 500=>x"4e00",
---- 501=>x"6a00", 502=>x"8f00", 503=>x"5700", 504=>x"4800",
---- 505=>x"4800", 506=>x"6300", 507=>x"8700", 508=>x"6600",
---- 509=>x"6100", 510=>x"6500", 511=>x"7700", 512=>x"7800",
---- 513=>x"7500", 514=>x"7300", 515=>x"7900", 516=>x"8100",
---- 517=>x"7d00", 518=>x"7e00", 519=>x"7e00", 520=>x"8800",
---- 521=>x"8400", 522=>x"8000", 523=>x"7f00", 524=>x"7700",
---- 525=>x"7700", 526=>x"8000", 527=>x"7e00", 528=>x"6600",
---- 529=>x"8200", 530=>x"7800", 531=>x"7c00", 532=>x"5c00",
---- 533=>x"7b00", 534=>x"7200", 535=>x"7800", 536=>x"6000",
---- 537=>x"6c00", 538=>x"6f00", 539=>x"7300", 540=>x"7300",
---- 541=>x"6a00", 542=>x"7800", 543=>x"7500", 544=>x"8000",
---- 545=>x"7600", 546=>x"7600", 547=>x"7900", 548=>x"8400",
---- 549=>x"8000", 550=>x"7700", 551=>x"8800", 552=>x"8200",
---- 553=>x"7d00", 554=>x"7a00", 555=>x"7a00", 556=>x"7c00",
---- 557=>x"7700", 558=>x"7f00", 559=>x"8400", 560=>x"8000",
---- 561=>x"7800", 562=>x"8400", 563=>x"8500", 564=>x"8300",
---- 565=>x"8100", 566=>x"8600", 567=>x"8800", 568=>x"8200",
---- 569=>x"8400", 570=>x"8a00", 571=>x"8900", 572=>x"8800",
---- 573=>x"8d00", 574=>x"8f00", 575=>x"8800", 576=>x"8900",
---- 577=>x"8f00", 578=>x"8b00", 579=>x"8500", 580=>x"8b00",
---- 581=>x"8f00", 582=>x"9000", 583=>x"8800", 584=>x"9400",
---- 585=>x"9200", 586=>x"8f00", 587=>x"8a00", 588=>x"9200",
---- 589=>x"9200", 590=>x"8f00", 591=>x"8a00", 592=>x"9400",
---- 593=>x"9200", 594=>x"9200", 595=>x"8c00", 596=>x"9300",
---- 597=>x"9300", 598=>x"9000", 599=>x"8b00", 600=>x"8d00",
---- 601=>x"9000", 602=>x"8f00", 603=>x"8900", 604=>x"8900",
---- 605=>x"8b00", 606=>x"8c00", 607=>x"8800", 608=>x"8700",
---- 609=>x"8600", 610=>x"7600", 611=>x"8700", 612=>x"7a00",
---- 613=>x"8500", 614=>x"8600", 615=>x"8300", 616=>x"8400",
---- 617=>x"8400", 618=>x"8500", 619=>x"8100", 620=>x"8400",
---- 621=>x"8200", 622=>x"8400", 623=>x"7f00", 624=>x"7f00",
---- 625=>x"7d00", 626=>x"8000", 627=>x"8500", 628=>x"7500",
---- 629=>x"7c00", 630=>x"8400", 631=>x"8900", 632=>x"7100",
---- 633=>x"8000", 634=>x"8700", 635=>x"8800", 636=>x"7500",
---- 637=>x"8500", 638=>x"8c00", 639=>x"8b00", 640=>x"7900",
---- 641=>x"8600", 642=>x"8900", 643=>x"8800", 644=>x"8000",
---- 645=>x"8500", 646=>x"8400", 647=>x"5b00", 648=>x"7a00",
---- 649=>x"8500", 650=>x"7c00", 651=>x"5400", 652=>x"7700",
---- 653=>x"7c00", 654=>x"7d00", 655=>x"7e00", 656=>x"8600",
---- 657=>x"8200", 658=>x"7c00", 659=>x"7f00", 660=>x"9100",
---- 661=>x"8f00", 662=>x"7a00", 663=>x"8300", 664=>x"9300",
---- 665=>x"9200", 666=>x"8f00", 667=>x"8a00", 668=>x"9400",
---- 669=>x"9400", 670=>x"9000", 671=>x"8f00", 672=>x"9300",
---- 673=>x"9300", 674=>x"9200", 675=>x"9400", 676=>x"9700",
---- 677=>x"9400", 678=>x"9700", 679=>x"9900", 680=>x"9500",
---- 681=>x"9900", 682=>x"9a00", 683=>x"9b00", 684=>x"9400",
---- 685=>x"9500", 686=>x"9900", 687=>x"9c00", 688=>x"9400",
---- 689=>x"9a00", 690=>x"9d00", 691=>x"a000", 692=>x"9400",
---- 693=>x"9200", 694=>x"9300", 695=>x"8d00", 696=>x"7b00",
---- 697=>x"7a00", 698=>x"7d00", 699=>x"7900", 700=>x"6300",
---- 701=>x"6100", 702=>x"5d00", 703=>x"5800", 704=>x"7000",
---- 705=>x"6e00", 706=>x"6a00", 707=>x"6600", 708=>x"8400",
---- 709=>x"8c00", 710=>x"9400", 711=>x"9300", 712=>x"8900",
---- 713=>x"9900", 714=>x"a900", 715=>x"b400", 716=>x"8500",
---- 717=>x"9500", 718=>x"9600", 719=>x"9d00", 720=>x"8000",
---- 721=>x"8900", 722=>x"8e00", 723=>x"9000", 724=>x"7b00",
---- 725=>x"8100", 726=>x"8700", 727=>x"7900", 728=>x"7600",
---- 729=>x"7600", 730=>x"7700", 731=>x"7800", 732=>x"7e00",
---- 733=>x"7b00", 734=>x"7600", 735=>x"7700", 736=>x"8f00",
---- 737=>x"9000", 738=>x"9000", 739=>x"9200", 740=>x"9900",
---- 741=>x"9f00", 742=>x"a400", 743=>x"a300", 744=>x"a400",
---- 745=>x"a600", 746=>x"a900", 747=>x"ac00", 748=>x"a600",
---- 749=>x"a900", 750=>x"ab00", 751=>x"a900", 752=>x"a400",
---- 753=>x"aa00", 754=>x"a600", 755=>x"a200", 756=>x"a700",
---- 757=>x"a800", 758=>x"a600", 759=>x"a500", 760=>x"aa00",
---- 761=>x"ab00", 762=>x"a800", 763=>x"a600", 764=>x"a800",
---- 765=>x"ac00", 766=>x"a800", 767=>x"a200", 768=>x"a400",
---- 769=>x"a400", 770=>x"5d00", 771=>x"9a00", 772=>x"a200",
---- 773=>x"a400", 774=>x"5f00", 775=>x"9800", 776=>x"a200",
---- 777=>x"a700", 778=>x"a600", 779=>x"a800", 780=>x"9a00",
---- 781=>x"9d00", 782=>x"9e00", 783=>x"a000", 784=>x"9700",
---- 785=>x"9500", 786=>x"9400", 787=>x"9600", 788=>x"8f00",
---- 789=>x"9000", 790=>x"9100", 791=>x"9200", 792=>x"8e00",
---- 793=>x"9000", 794=>x"8f00", 795=>x"9500", 796=>x"8e00",
---- 797=>x"8f00", 798=>x"9000", 799=>x"9500", 800=>x"8f00",
---- 801=>x"9000", 802=>x"9400", 803=>x"9800", 804=>x"8e00",
---- 805=>x"9500", 806=>x"9700", 807=>x"9d00", 808=>x"9100",
---- 809=>x"9300", 810=>x"9900", 811=>x"9d00", 812=>x"9200",
---- 813=>x"9700", 814=>x"9c00", 815=>x"a200", 816=>x"9500",
---- 817=>x"9b00", 818=>x"9e00", 819=>x"a100", 820=>x"9800",
---- 821=>x"9b00", 822=>x"9f00", 823=>x"a100", 824=>x"9800",
---- 825=>x"9c00", 826=>x"a200", 827=>x"a200", 828=>x"9900",
---- 829=>x"9d00", 830=>x"a100", 831=>x"a000", 832=>x"6800",
---- 833=>x"9900", 834=>x"a000", 835=>x"a100", 836=>x"9700",
---- 837=>x"9800", 838=>x"9c00", 839=>x"a000", 840=>x"9700",
---- 841=>x"9800", 842=>x"9b00", 843=>x"9e00", 844=>x"9500",
---- 845=>x"9800", 846=>x"9a00", 847=>x"9d00", 848=>x"9400",
---- 849=>x"9600", 850=>x"9900", 851=>x"9b00", 852=>x"9500",
---- 853=>x"9600", 854=>x"9700", 855=>x"9a00", 856=>x"9300",
---- 857=>x"9600", 858=>x"9900", 859=>x"9e00", 860=>x"9000",
---- 861=>x"9500", 862=>x"9900", 863=>x"6600", 864=>x"9200",
---- 865=>x"9300", 866=>x"9700", 867=>x"9900", 868=>x"9200",
---- 869=>x"9200", 870=>x"9500", 871=>x"9700", 872=>x"9300",
---- 873=>x"9400", 874=>x"9500", 875=>x"9600", 876=>x"9100",
---- 877=>x"9300", 878=>x"9500", 879=>x"9400", 880=>x"8f00",
---- 881=>x"9200", 882=>x"9300", 883=>x"9200", 884=>x"8d00",
---- 885=>x"9000", 886=>x"9300", 887=>x"9400", 888=>x"8c00",
---- 889=>x"8e00", 890=>x"9400", 891=>x"9700", 892=>x"8f00",
---- 893=>x"8e00", 894=>x"9300", 895=>x"9300", 896=>x"8e00",
---- 897=>x"8e00", 898=>x"9100", 899=>x"9200", 900=>x"8e00",
---- 901=>x"8e00", 902=>x"9100", 903=>x"9000", 904=>x"8b00",
---- 905=>x"8e00", 906=>x"9200", 907=>x"9200", 908=>x"8e00",
---- 909=>x"8e00", 910=>x"8f00", 911=>x"9200", 912=>x"9000",
---- 913=>x"8d00", 914=>x"8f00", 915=>x"9200", 916=>x"8e00",
---- 917=>x"8d00", 918=>x"8f00", 919=>x"9000", 920=>x"8c00",
---- 921=>x"8f00", 922=>x"8e00", 923=>x"9000", 924=>x"8b00",
---- 925=>x"8d00", 926=>x"9100", 927=>x"9100", 928=>x"8c00",
---- 929=>x"8a00", 930=>x"8e00", 931=>x"9100", 932=>x"7500",
---- 933=>x"8a00", 934=>x"8e00", 935=>x"8e00", 936=>x"8600",
---- 937=>x"8900", 938=>x"8e00", 939=>x"8c00", 940=>x"8800",
---- 941=>x"7400", 942=>x"8c00", 943=>x"8b00", 944=>x"8a00",
---- 945=>x"8a00", 946=>x"8a00", 947=>x"8700", 948=>x"8600",
---- 949=>x"8d00", 950=>x"8900", 951=>x"8900", 952=>x"8900",
---- 953=>x"8c00", 954=>x"8a00", 955=>x"8b00", 956=>x"8800",
---- 957=>x"8800", 958=>x"8900", 959=>x"8c00", 960=>x"8700",
---- 961=>x"8900", 962=>x"8b00", 963=>x"8b00", 964=>x"7800",
---- 965=>x"8b00", 966=>x"8b00", 967=>x"7200", 968=>x"8a00",
---- 969=>x"8d00", 970=>x"8a00", 971=>x"8e00", 972=>x"8b00",
---- 973=>x"8e00", 974=>x"8b00", 975=>x"8e00", 976=>x"8e00",
---- 977=>x"8d00", 978=>x"8b00", 979=>x"8c00", 980=>x"8f00",
---- 981=>x"9000", 982=>x"8b00", 983=>x"8900", 984=>x"8e00",
---- 985=>x"8e00", 986=>x"8c00", 987=>x"8900", 988=>x"9000",
---- 989=>x"8d00", 990=>x"9000", 991=>x"8e00", 992=>x"9000",
---- 993=>x"8f00", 994=>x"9200", 995=>x"8e00", 996=>x"9100",
---- 997=>x"8f00", 998=>x"9500", 999=>x"9300", 1000=>x"9100",
---- 1001=>x"6f00", 1002=>x"9400", 1003=>x"9200", 1004=>x"9100",
---- 1005=>x"9200", 1006=>x"9700", 1007=>x"9100", 1008=>x"9300",
---- 1009=>x"9200", 1010=>x"9200", 1011=>x"9300", 1012=>x"9400",
---- 1013=>x"9100", 1014=>x"9100", 1015=>x"9100", 1016=>x"9200",
---- 1017=>x"9200", 1018=>x"9300", 1019=>x"9200", 1020=>x"9300",
---- 1021=>x"9000", 1022=>x"9200", 1023=>x"9000"),
----
---- 37 => (0=>x"7f00", 1=>x"7f00", 2=>x"7f00", 3=>x"8000", 4=>x"7f00",
---- 5=>x"7f00", 6=>x"7f00", 7=>x"8000", 8=>x"8000",
---- 9=>x"7f00", 10=>x"8000", 11=>x"8000", 12=>x"8000",
---- 13=>x"8100", 14=>x"7e00", 15=>x"7c00", 16=>x"8100",
---- 17=>x"7e00", 18=>x"7d00", 19=>x"7e00", 20=>x"8000",
---- 21=>x"7e00", 22=>x"7f00", 23=>x"7f00", 24=>x"7e00",
---- 25=>x"7f00", 26=>x"8100", 27=>x"7f00", 28=>x"7f00",
---- 29=>x"8100", 30=>x"8200", 31=>x"7f00", 32=>x"8000",
---- 33=>x"8000", 34=>x"8100", 35=>x"8200", 36=>x"8200",
---- 37=>x"7d00", 38=>x"7e00", 39=>x"8200", 40=>x"7e00",
---- 41=>x"7e00", 42=>x"8000", 43=>x"7f00", 44=>x"7e00",
---- 45=>x"7d00", 46=>x"8300", 47=>x"7f00", 48=>x"7d00",
---- 49=>x"7b00", 50=>x"8000", 51=>x"8100", 52=>x"7e00",
---- 53=>x"8000", 54=>x"8000", 55=>x"7e00", 56=>x"7c00",
---- 57=>x"8000", 58=>x"8100", 59=>x"7d00", 60=>x"7e00",
---- 61=>x"7f00", 62=>x"8000", 63=>x"8200", 64=>x"7f00",
---- 65=>x"8000", 66=>x"7f00", 67=>x"8000", 68=>x"8000",
---- 69=>x"7f00", 70=>x"8000", 71=>x"7f00", 72=>x"7c00",
---- 73=>x"7d00", 74=>x"7e00", 75=>x"7e00", 76=>x"8000",
---- 77=>x"7d00", 78=>x"7d00", 79=>x"7f00", 80=>x"7d00",
---- 81=>x"7c00", 82=>x"8000", 83=>x"7e00", 84=>x"7e00",
---- 85=>x"7e00", 86=>x"8000", 87=>x"7e00", 88=>x"7f00",
---- 89=>x"7d00", 90=>x"7e00", 91=>x"8000", 92=>x"7f00",
---- 93=>x"8000", 94=>x"8100", 95=>x"7f00", 96=>x"7e00",
---- 97=>x"8000", 98=>x"7d00", 99=>x"7d00", 100=>x"7f00",
---- 101=>x"7d00", 102=>x"8000", 103=>x"7c00", 104=>x"7c00",
---- 105=>x"7c00", 106=>x"7d00", 107=>x"7e00", 108=>x"7e00",
---- 109=>x"7b00", 110=>x"7b00", 111=>x"7a00", 112=>x"7c00",
---- 113=>x"7a00", 114=>x"7b00", 115=>x"7900", 116=>x"7900",
---- 117=>x"7d00", 118=>x"7b00", 119=>x"7a00", 120=>x"7600",
---- 121=>x"7900", 122=>x"7a00", 123=>x"7800", 124=>x"7800",
---- 125=>x"7600", 126=>x"7700", 127=>x"7800", 128=>x"7700",
---- 129=>x"7800", 130=>x"7700", 131=>x"7700", 132=>x"7300",
---- 133=>x"7300", 134=>x"7300", 135=>x"7700", 136=>x"6e00",
---- 137=>x"7100", 138=>x"7100", 139=>x"7300", 140=>x"6a00",
---- 141=>x"6c00", 142=>x"6e00", 143=>x"7200", 144=>x"6400",
---- 145=>x"6700", 146=>x"6b00", 147=>x"6c00", 148=>x"a700",
---- 149=>x"6100", 150=>x"6300", 151=>x"6900", 152=>x"7600",
---- 153=>x"5500", 154=>x"5e00", 155=>x"6500", 156=>x"c400",
---- 157=>x"6500", 158=>x"5500", 159=>x"5a00", 160=>x"e600",
---- 161=>x"9d00", 162=>x"4e00", 163=>x"5200", 164=>x"e300",
---- 165=>x"d000", 166=>x"7700", 167=>x"4b00", 168=>x"e000",
---- 169=>x"e300", 170=>x"c400", 171=>x"6000", 172=>x"e000",
---- 173=>x"de00", 174=>x"e200", 175=>x"a500", 176=>x"d500",
---- 177=>x"df00", 178=>x"df00", 179=>x"da00", 180=>x"d500",
---- 181=>x"de00", 182=>x"e100", 183=>x"de00", 184=>x"da00",
---- 185=>x"df00", 186=>x"e500", 187=>x"e000", 188=>x"d400",
---- 189=>x"d800", 190=>x"dc00", 191=>x"e100", 192=>x"ce00",
---- 193=>x"d100", 194=>x"d400", 195=>x"d600", 196=>x"d400",
---- 197=>x"d300", 198=>x"d400", 199=>x"d400", 200=>x"d000",
---- 201=>x"d300", 202=>x"d200", 203=>x"d400", 204=>x"d100",
---- 205=>x"d100", 206=>x"d400", 207=>x"ce00", 208=>x"cf00",
---- 209=>x"d000", 210=>x"d100", 211=>x"cc00", 212=>x"d200",
---- 213=>x"d100", 214=>x"d300", 215=>x"d100", 216=>x"cf00",
---- 217=>x"cc00", 218=>x"ca00", 219=>x"cd00", 220=>x"ca00",
---- 221=>x"cd00", 222=>x"cb00", 223=>x"cd00", 224=>x"ca00",
---- 225=>x"d100", 226=>x"d400", 227=>x"d100", 228=>x"ce00",
---- 229=>x"cf00", 230=>x"d000", 231=>x"d400", 232=>x"ca00",
---- 233=>x"ce00", 234=>x"cf00", 235=>x"d000", 236=>x"c800",
---- 237=>x"cb00", 238=>x"ce00", 239=>x"cf00", 240=>x"cf00",
---- 241=>x"c700", 242=>x"ca00", 243=>x"d000", 244=>x"c900",
---- 245=>x"c700", 246=>x"c400", 247=>x"3300", 248=>x"c200",
---- 249=>x"c900", 250=>x"c700", 251=>x"c900", 252=>x"cb00",
---- 253=>x"c800", 254=>x"cb00", 255=>x"cb00", 256=>x"ca00",
---- 257=>x"d000", 258=>x"cf00", 259=>x"cb00", 260=>x"c200",
---- 261=>x"ca00", 262=>x"bf00", 263=>x"ba00", 264=>x"b100",
---- 265=>x"a200", 266=>x"b200", 267=>x"c600", 268=>x"9e00",
---- 269=>x"a800", 270=>x"c200", 271=>x"c600", 272=>x"b300",
---- 273=>x"c200", 274=>x"bd00", 275=>x"c000", 276=>x"bd00",
---- 277=>x"be00", 278=>x"c100", 279=>x"c600", 280=>x"be00",
---- 281=>x"bd00", 282=>x"ba00", 283=>x"bd00", 284=>x"b200",
---- 285=>x"b500", 286=>x"b500", 287=>x"b900", 288=>x"bb00",
---- 289=>x"bc00", 290=>x"c200", 291=>x"be00", 292=>x"bc00",
---- 293=>x"bf00", 294=>x"c200", 295=>x"c000", 296=>x"ba00",
---- 297=>x"bb00", 298=>x"c000", 299=>x"bd00", 300=>x"bf00",
---- 301=>x"b800", 302=>x"bb00", 303=>x"bf00", 304=>x"c000",
---- 305=>x"bd00", 306=>x"b600", 307=>x"b500", 308=>x"bd00",
---- 309=>x"bc00", 310=>x"b400", 311=>x"af00", 312=>x"b700",
---- 313=>x"b200", 314=>x"b200", 315=>x"b100", 316=>x"af00",
---- 317=>x"b200", 318=>x"af00", 319=>x"ae00", 320=>x"5600",
---- 321=>x"aa00", 322=>x"ae00", 323=>x"5000", 324=>x"ab00",
---- 325=>x"a600", 326=>x"aa00", 327=>x"af00", 328=>x"ad00",
---- 329=>x"5500", 330=>x"a300", 331=>x"a700", 332=>x"a300",
---- 333=>x"ab00", 334=>x"9f00", 335=>x"9f00", 336=>x"9800",
---- 337=>x"9d00", 338=>x"9f00", 339=>x"9600", 340=>x"9c00",
---- 341=>x"9000", 342=>x"9b00", 343=>x"9400", 344=>x"9b00",
---- 345=>x"8a00", 346=>x"9700", 347=>x"b300", 348=>x"8800",
---- 349=>x"a100", 350=>x"bb00", 351=>x"c100", 352=>x"a100",
---- 353=>x"c300", 354=>x"b400", 355=>x"9e00", 356=>x"c100",
---- 357=>x"a400", 358=>x"9700", 359=>x"a100", 360=>x"9900",
---- 361=>x"9200", 362=>x"ae00", 363=>x"c000", 364=>x"9600",
---- 365=>x"b900", 366=>x"cb00", 367=>x"cc00", 368=>x"b300",
---- 369=>x"c600", 370=>x"c900", 371=>x"cb00", 372=>x"be00",
---- 373=>x"bc00", 374=>x"be00", 375=>x"3f00", 376=>x"bf00",
---- 377=>x"b800", 378=>x"b800", 379=>x"b800", 380=>x"b500",
---- 381=>x"b200", 382=>x"b400", 383=>x"b900", 384=>x"b300",
---- 385=>x"b500", 386=>x"ba00", 387=>x"bc00", 388=>x"b400",
---- 389=>x"b400", 390=>x"b800", 391=>x"bb00", 392=>x"b300",
---- 393=>x"b700", 394=>x"ba00", 395=>x"b700", 396=>x"b700",
---- 397=>x"b600", 398=>x"b800", 399=>x"b600", 400=>x"b700",
---- 401=>x"b400", 402=>x"b300", 403=>x"b600", 404=>x"b500",
---- 405=>x"b300", 406=>x"b700", 407=>x"b300", 408=>x"b400",
---- 409=>x"b800", 410=>x"b800", 411=>x"b300", 412=>x"b400",
---- 413=>x"b500", 414=>x"b400", 415=>x"ad00", 416=>x"b400",
---- 417=>x"b200", 418=>x"ad00", 419=>x"ac00", 420=>x"ae00",
---- 421=>x"ae00", 422=>x"af00", 423=>x"b000", 424=>x"ae00",
---- 425=>x"af00", 426=>x"b200", 427=>x"ad00", 428=>x"b100",
---- 429=>x"b000", 430=>x"ab00", 431=>x"af00", 432=>x"b000",
---- 433=>x"a600", 434=>x"9f00", 435=>x"ac00", 436=>x"ab00",
---- 437=>x"9d00", 438=>x"9f00", 439=>x"a800", 440=>x"a400",
---- 441=>x"a000", 442=>x"a900", 443=>x"ae00", 444=>x"9c00",
---- 445=>x"a600", 446=>x"ab00", 447=>x"b100", 448=>x"5a00",
---- 449=>x"ac00", 450=>x"b100", 451=>x"b700", 452=>x"a900",
---- 453=>x"ad00", 454=>x"b000", 455=>x"bb00", 456=>x"a900",
---- 457=>x"5100", 458=>x"b500", 459=>x"be00", 460=>x"a900",
---- 461=>x"ae00", 462=>x"b800", 463=>x"bb00", 464=>x"a900",
---- 465=>x"b100", 466=>x"b700", 467=>x"4400", 468=>x"af00",
---- 469=>x"af00", 470=>x"b500", 471=>x"b900", 472=>x"b100",
---- 473=>x"b200", 474=>x"b400", 475=>x"b800", 476=>x"af00",
---- 477=>x"b400", 478=>x"b400", 479=>x"b600", 480=>x"b000",
---- 481=>x"b200", 482=>x"b000", 483=>x"b200", 484=>x"b200",
---- 485=>x"b100", 486=>x"b200", 487=>x"b700", 488=>x"b100",
---- 489=>x"af00", 490=>x"b000", 491=>x"b100", 492=>x"b100",
---- 493=>x"b100", 494=>x"b200", 495=>x"af00", 496=>x"af00",
---- 497=>x"b400", 498=>x"b200", 499=>x"ad00", 500=>x"ac00",
---- 501=>x"ad00", 502=>x"ab00", 503=>x"ab00", 504=>x"a300",
---- 505=>x"a700", 506=>x"a700", 507=>x"a900", 508=>x"9400",
---- 509=>x"9d00", 510=>x"9e00", 511=>x"a400", 512=>x"8600",
---- 513=>x"9400", 514=>x"9b00", 515=>x"a100", 516=>x"8900",
---- 517=>x"8c00", 518=>x"9400", 519=>x"9d00", 520=>x"8800",
---- 521=>x"8d00", 522=>x"6e00", 523=>x"9600", 524=>x"8500",
---- 525=>x"8900", 526=>x"9100", 527=>x"9500", 528=>x"8600",
---- 529=>x"8800", 530=>x"8f00", 531=>x"9200", 532=>x"8300",
---- 533=>x"8600", 534=>x"8b00", 535=>x"8e00", 536=>x"7a00",
---- 537=>x"8200", 538=>x"8700", 539=>x"8d00", 540=>x"7800",
---- 541=>x"8100", 542=>x"8800", 543=>x"8e00", 544=>x"7d00",
---- 545=>x"8100", 546=>x"8500", 547=>x"8900", 548=>x"7f00",
---- 549=>x"8000", 550=>x"8000", 551=>x"8c00", 552=>x"7d00",
---- 553=>x"8000", 554=>x"8000", 555=>x"8b00", 556=>x"8000",
---- 557=>x"8100", 558=>x"7f00", 559=>x"8900", 560=>x"8200",
---- 561=>x"8100", 562=>x"7d00", 563=>x"8400", 564=>x"8400",
---- 565=>x"8000", 566=>x"7f00", 567=>x"8000", 568=>x"8100",
---- 569=>x"7f00", 570=>x"8100", 571=>x"8000", 572=>x"8400",
---- 573=>x"8100", 574=>x"8300", 575=>x"7f00", 576=>x"8300",
---- 577=>x"8200", 578=>x"8100", 579=>x"8000", 580=>x"8100",
---- 581=>x"8200", 582=>x"7f00", 583=>x"7c00", 584=>x"8300",
---- 585=>x"8600", 586=>x"8100", 587=>x"8100", 588=>x"8300",
---- 589=>x"8500", 590=>x"8300", 591=>x"8000", 592=>x"8700",
---- 593=>x"8400", 594=>x"8000", 595=>x"8100", 596=>x"8700",
---- 597=>x"8100", 598=>x"7e00", 599=>x"8500", 600=>x"8500",
---- 601=>x"7d00", 602=>x"7e00", 603=>x"8200", 604=>x"8100",
---- 605=>x"7d00", 606=>x"7d00", 607=>x"8000", 608=>x"7d00",
---- 609=>x"7f00", 610=>x"7c00", 611=>x"7e00", 612=>x"8000",
---- 613=>x"7c00", 614=>x"7900", 615=>x"7c00", 616=>x"8000",
---- 617=>x"7b00", 618=>x"7800", 619=>x"7c00", 620=>x"7c00",
---- 621=>x"7b00", 622=>x"7800", 623=>x"7a00", 624=>x"7e00",
---- 625=>x"7b00", 626=>x"7b00", 627=>x"7600", 628=>x"8200",
---- 629=>x"7d00", 630=>x"7c00", 631=>x"7900", 632=>x"8900",
---- 633=>x"8900", 634=>x"8300", 635=>x"7c00", 636=>x"8c00",
---- 637=>x"8e00", 638=>x"8d00", 639=>x"8200", 640=>x"8500",
---- 641=>x"8b00", 642=>x"8900", 643=>x"8700", 644=>x"3e00",
---- 645=>x"4f00", 646=>x"6900", 647=>x"7200", 648=>x"3c00",
---- 649=>x"5000", 650=>x"6000", 651=>x"a700", 652=>x"7c00",
---- 653=>x"8000", 654=>x"8100", 655=>x"7600", 656=>x"8300",
---- 657=>x"8400", 658=>x"8600", 659=>x"7d00", 660=>x"8100",
---- 661=>x"8600", 662=>x"9100", 663=>x"8e00", 664=>x"8b00",
---- 665=>x"9300", 666=>x"a700", 667=>x"b300", 668=>x"9500",
---- 669=>x"a000", 670=>x"b900", 671=>x"c500", 672=>x"9900",
---- 673=>x"a700", 674=>x"c400", 675=>x"cc00", 676=>x"9f00",
---- 677=>x"ae00", 678=>x"cc00", 679=>x"ce00", 680=>x"a200",
---- 681=>x"b200", 682=>x"d100", 683=>x"cf00", 684=>x"a200",
---- 685=>x"b500", 686=>x"cd00", 687=>x"d400", 688=>x"a400",
---- 689=>x"a900", 690=>x"b400", 691=>x"bb00", 692=>x"8b00",
---- 693=>x"8600", 694=>x"8e00", 695=>x"9000", 696=>x"7800",
---- 697=>x"7400", 698=>x"7c00", 699=>x"8500", 700=>x"5e00",
---- 701=>x"6400", 702=>x"8f00", 703=>x"7600", 704=>x"6a00",
---- 705=>x"6c00", 706=>x"7500", 707=>x"7d00", 708=>x"9700",
---- 709=>x"9900", 710=>x"9f00", 711=>x"ae00", 712=>x"b800",
---- 713=>x"b900", 714=>x"b800", 715=>x"c800", 716=>x"a500",
---- 717=>x"a300", 718=>x"9a00", 719=>x"9e00", 720=>x"9200",
---- 721=>x"9600", 722=>x"9100", 723=>x"8b00", 724=>x"8e00",
---- 725=>x"8d00", 726=>x"8900", 727=>x"8700", 728=>x"7d00",
---- 729=>x"7800", 730=>x"7600", 731=>x"7700", 732=>x"7900",
---- 733=>x"7d00", 734=>x"8100", 735=>x"7300", 736=>x"9000",
---- 737=>x"6a00", 738=>x"9a00", 739=>x"9b00", 740=>x"9e00",
---- 741=>x"9b00", 742=>x"9c00", 743=>x"9e00", 744=>x"a400",
---- 745=>x"9e00", 746=>x"9c00", 747=>x"9d00", 748=>x"a900",
---- 749=>x"a300", 750=>x"a300", 751=>x"a200", 752=>x"a900",
---- 753=>x"a800", 754=>x"a700", 755=>x"a400", 756=>x"a900",
---- 757=>x"ad00", 758=>x"af00", 759=>x"a400", 760=>x"a900",
---- 761=>x"aa00", 762=>x"a800", 763=>x"9f00", 764=>x"a300",
---- 765=>x"a300", 766=>x"9e00", 767=>x"9b00", 768=>x"9a00",
---- 769=>x"9a00", 770=>x"9b00", 771=>x"9400", 772=>x"9800",
---- 773=>x"9900", 774=>x"9200", 775=>x"8500", 776=>x"ad00",
---- 777=>x"aa00", 778=>x"a200", 779=>x"9d00", 780=>x"a100",
---- 781=>x"a000", 782=>x"a900", 783=>x"b200", 784=>x"9900",
---- 785=>x"9c00", 786=>x"a600", 787=>x"ad00", 788=>x"6700",
---- 789=>x"a100", 790=>x"aa00", 791=>x"ae00", 792=>x"9800",
---- 793=>x"a400", 794=>x"ac00", 795=>x"b000", 796=>x"9a00",
---- 797=>x"a600", 798=>x"ab00", 799=>x"b300", 800=>x"9f00",
---- 801=>x"a700", 802=>x"ae00", 803=>x"b700", 804=>x"a200",
---- 805=>x"a900", 806=>x"ae00", 807=>x"b500", 808=>x"a600",
---- 809=>x"ad00", 810=>x"b100", 811=>x"b500", 812=>x"a400",
---- 813=>x"a900", 814=>x"ac00", 815=>x"b300", 816=>x"a400",
---- 817=>x"a700", 818=>x"a800", 819=>x"b000", 820=>x"a300",
---- 821=>x"a600", 822=>x"a900", 823=>x"4f00", 824=>x"a400",
---- 825=>x"a800", 826=>x"a700", 827=>x"aa00", 828=>x"a200",
---- 829=>x"a500", 830=>x"a500", 831=>x"a900", 832=>x"a100",
---- 833=>x"a200", 834=>x"a500", 835=>x"a800", 836=>x"a100",
---- 837=>x"a100", 838=>x"a400", 839=>x"a500", 840=>x"9f00",
---- 841=>x"a200", 842=>x"a200", 843=>x"a500", 844=>x"a100",
---- 845=>x"a000", 846=>x"a300", 847=>x"a500", 848=>x"9e00",
---- 849=>x"9f00", 850=>x"a200", 851=>x"a400", 852=>x"9b00",
---- 853=>x"9e00", 854=>x"9f00", 855=>x"a200", 856=>x"9c00",
---- 857=>x"9d00", 858=>x"a000", 859=>x"9f00", 860=>x"9a00",
---- 861=>x"9c00", 862=>x"9b00", 863=>x"a000", 864=>x"9a00",
---- 865=>x"9b00", 866=>x"9e00", 867=>x"a000", 868=>x"9900",
---- 869=>x"9a00", 870=>x"9d00", 871=>x"a100", 872=>x"9c00",
---- 873=>x"9c00", 874=>x"9f00", 875=>x"9f00", 876=>x"9b00",
---- 877=>x"9b00", 878=>x"9d00", 879=>x"9e00", 880=>x"9700",
---- 881=>x"9a00", 882=>x"9b00", 883=>x"9d00", 884=>x"9500",
---- 885=>x"9900", 886=>x"9b00", 887=>x"9e00", 888=>x"9600",
---- 889=>x"9a00", 890=>x"9c00", 891=>x"9b00", 892=>x"9600",
---- 893=>x"9800", 894=>x"9700", 895=>x"9a00", 896=>x"9400",
---- 897=>x"9400", 898=>x"9600", 899=>x"9d00", 900=>x"9300",
---- 901=>x"9500", 902=>x"9800", 903=>x"9b00", 904=>x"9400",
---- 905=>x"6b00", 906=>x"9600", 907=>x"9a00", 908=>x"9400",
---- 909=>x"9600", 910=>x"9700", 911=>x"9800", 912=>x"9200",
---- 913=>x"9400", 914=>x"9300", 915=>x"9800", 916=>x"9400",
---- 917=>x"9400", 918=>x"9400", 919=>x"9700", 920=>x"9400",
---- 921=>x"9500", 922=>x"9400", 923=>x"9700", 924=>x"9400",
---- 925=>x"9500", 926=>x"9600", 927=>x"9700", 928=>x"9000",
---- 929=>x"9100", 930=>x"9500", 931=>x"6900", 932=>x"8f00",
---- 933=>x"9200", 934=>x"9100", 935=>x"9500", 936=>x"8f00",
---- 937=>x"8e00", 938=>x"9000", 939=>x"9300", 940=>x"8f00",
---- 941=>x"9200", 942=>x"8f00", 943=>x"9200", 944=>x"8c00",
---- 945=>x"8f00", 946=>x"8f00", 947=>x"9100", 948=>x"8b00",
---- 949=>x"8d00", 950=>x"7200", 951=>x"8f00", 952=>x"8c00",
---- 953=>x"8b00", 954=>x"8b00", 955=>x"8e00", 956=>x"8c00",
---- 957=>x"8800", 958=>x"8b00", 959=>x"8e00", 960=>x"8c00",
---- 961=>x"8a00", 962=>x"8b00", 963=>x"8c00", 964=>x"8c00",
---- 965=>x"8e00", 966=>x"7300", 967=>x"8c00", 968=>x"8900",
---- 969=>x"8a00", 970=>x"8900", 971=>x"8a00", 972=>x"8b00",
---- 973=>x"8a00", 974=>x"8b00", 975=>x"8a00", 976=>x"8b00",
---- 977=>x"8b00", 978=>x"8c00", 979=>x"8b00", 980=>x"8c00",
---- 981=>x"8f00", 982=>x"8d00", 983=>x"8d00", 984=>x"8900",
---- 985=>x"8c00", 986=>x"8f00", 987=>x"8e00", 988=>x"8b00",
---- 989=>x"8e00", 990=>x"8f00", 991=>x"8e00", 992=>x"8d00",
---- 993=>x"8f00", 994=>x"8b00", 995=>x"8d00", 996=>x"8e00",
---- 997=>x"8f00", 998=>x"8f00", 999=>x"9200", 1000=>x"9100",
---- 1001=>x"9000", 1002=>x"8f00", 1003=>x"9100", 1004=>x"6a00",
---- 1005=>x"9400", 1006=>x"9000", 1007=>x"9400", 1008=>x"9500",
---- 1009=>x"9100", 1010=>x"9100", 1011=>x"9700", 1012=>x"9700",
---- 1013=>x"9500", 1014=>x"6a00", 1015=>x"9600", 1016=>x"9500",
---- 1017=>x"9500", 1018=>x"9400", 1019=>x"9100", 1020=>x"9400",
---- 1021=>x"9400", 1022=>x"9700", 1023=>x"9600"),
----
---- 38 => (0=>x"7d00", 1=>x"7c00", 2=>x"7800", 3=>x"7a00", 4=>x"8300",
---- 5=>x"7b00", 6=>x"7800", 7=>x"7900", 8=>x"7a00",
---- 9=>x"7a00", 10=>x"7a00", 11=>x"7800", 12=>x"7c00",
---- 13=>x"7900", 14=>x"7b00", 15=>x"7800", 16=>x"7c00",
---- 17=>x"7c00", 18=>x"7800", 19=>x"7700", 20=>x"7c00",
---- 21=>x"7b00", 22=>x"7600", 23=>x"7700", 24=>x"7c00",
---- 25=>x"7b00", 26=>x"7a00", 27=>x"7a00", 28=>x"7b00",
---- 29=>x"8300", 30=>x"7c00", 31=>x"7900", 32=>x"8000",
---- 33=>x"7c00", 34=>x"7900", 35=>x"7900", 36=>x"7e00",
---- 37=>x"7d00", 38=>x"7d00", 39=>x"7a00", 40=>x"7e00",
---- 41=>x"7c00", 42=>x"7b00", 43=>x"7b00", 44=>x"7e00",
---- 45=>x"7b00", 46=>x"7b00", 47=>x"7a00", 48=>x"7d00",
---- 49=>x"7c00", 50=>x"7e00", 51=>x"7900", 52=>x"7e00",
---- 53=>x"7c00", 54=>x"7a00", 55=>x"7a00", 56=>x"7d00",
---- 57=>x"7b00", 58=>x"7b00", 59=>x"7900", 60=>x"8000",
---- 61=>x"8100", 62=>x"7d00", 63=>x"7700", 64=>x"7c00",
---- 65=>x"8000", 66=>x"7c00", 67=>x"7900", 68=>x"7d00",
---- 69=>x"7e00", 70=>x"7d00", 71=>x"7a00", 72=>x"8000",
---- 73=>x"7c00", 74=>x"7b00", 75=>x"7900", 76=>x"8100",
---- 77=>x"7d00", 78=>x"7c00", 79=>x"7a00", 80=>x"7d00",
---- 81=>x"7c00", 82=>x"7c00", 83=>x"7800", 84=>x"7d00",
---- 85=>x"7900", 86=>x"7a00", 87=>x"7a00", 88=>x"7d00",
---- 89=>x"7a00", 90=>x"7c00", 91=>x"7a00", 92=>x"7b00",
---- 93=>x"7e00", 94=>x"7d00", 95=>x"7800", 96=>x"8100",
---- 97=>x"7d00", 98=>x"7a00", 99=>x"7700", 100=>x"7d00",
---- 101=>x"7c00", 102=>x"7900", 103=>x"7700", 104=>x"7c00",
---- 105=>x"7600", 106=>x"7700", 107=>x"7900", 108=>x"7b00",
---- 109=>x"7800", 110=>x"7900", 111=>x"7800", 112=>x"7b00",
---- 113=>x"7700", 114=>x"7600", 115=>x"7500", 116=>x"7700",
---- 117=>x"7400", 118=>x"7100", 119=>x"7300", 120=>x"7800",
---- 121=>x"7500", 122=>x"7300", 123=>x"7400", 124=>x"7700",
---- 125=>x"7600", 126=>x"7500", 127=>x"7300", 128=>x"7500",
---- 129=>x"7400", 130=>x"7500", 131=>x"7200", 132=>x"7400",
---- 133=>x"7500", 134=>x"7400", 135=>x"7100", 136=>x"7300",
---- 137=>x"7200", 138=>x"7200", 139=>x"7100", 140=>x"7200",
---- 141=>x"7100", 142=>x"8d00", 143=>x"6f00", 144=>x"7200",
---- 145=>x"6e00", 146=>x"7000", 147=>x"6f00", 148=>x"6e00",
---- 149=>x"6c00", 150=>x"6e00", 151=>x"6d00", 152=>x"6c00",
---- 153=>x"6c00", 154=>x"6c00", 155=>x"6b00", 156=>x"6600",
---- 157=>x"9700", 158=>x"9600", 159=>x"6a00", 160=>x"5d00",
---- 161=>x"6200", 162=>x"6700", 163=>x"6500", 164=>x"5900",
---- 165=>x"5b00", 166=>x"6400", 167=>x"6500", 168=>x"b000",
---- 169=>x"5700", 170=>x"5c00", 171=>x"6000", 172=>x"5400",
---- 173=>x"4e00", 174=>x"5400", 175=>x"5c00", 176=>x"9a00",
---- 177=>x"4f00", 178=>x"4e00", 179=>x"5400", 180=>x"d500",
---- 181=>x"7900", 182=>x"4800", 183=>x"5100", 184=>x"de00",
---- 185=>x"bf00", 186=>x"6100", 187=>x"4800", 188=>x"df00",
---- 189=>x"e400", 190=>x"a200", 191=>x"4d00", 192=>x"d900",
---- 193=>x"de00", 194=>x"d300", 195=>x"9b00", 196=>x"d600",
---- 197=>x"da00", 198=>x"e000", 199=>x"e200", 200=>x"d600",
---- 201=>x"d900", 202=>x"da00", 203=>x"de00", 204=>x"d300",
---- 205=>x"d600", 206=>x"d500", 207=>x"d500", 208=>x"d200",
---- 209=>x"d600", 210=>x"d300", 211=>x"d300", 212=>x"cd00",
---- 213=>x"d600", 214=>x"d900", 215=>x"d700", 216=>x"c900",
---- 217=>x"cf00", 218=>x"d300", 219=>x"d700", 220=>x"cc00",
---- 221=>x"d000", 222=>x"d400", 223=>x"d700", 224=>x"cd00",
---- 225=>x"ce00", 226=>x"d200", 227=>x"d400", 228=>x"d000",
---- 229=>x"ca00", 230=>x"cf00", 231=>x"d300", 232=>x"d300",
---- 233=>x"cb00", 234=>x"cd00", 235=>x"d400", 236=>x"cf00",
---- 237=>x"d100", 238=>x"d100", 239=>x"d000", 240=>x"ce00",
---- 241=>x"ce00", 242=>x"cf00", 243=>x"cd00", 244=>x"cf00",
---- 245=>x"cc00", 246=>x"ca00", 247=>x"cc00", 248=>x"ce00",
---- 249=>x"d000", 250=>x"cb00", 251=>x"d000", 252=>x"d100",
---- 253=>x"d100", 254=>x"cd00", 255=>x"ce00", 256=>x"ca00",
---- 257=>x"c600", 258=>x"c300", 259=>x"c700", 260=>x"c400",
---- 261=>x"3f00", 262=>x"c500", 263=>x"cc00", 264=>x"cb00",
---- 265=>x"c700", 266=>x"c600", 267=>x"cc00", 268=>x"c700",
---- 269=>x"c800", 270=>x"c800", 271=>x"cd00", 272=>x"c400",
---- 273=>x"c900", 274=>x"c900", 275=>x"c900", 276=>x"c600",
---- 277=>x"c700", 278=>x"c500", 279=>x"c600", 280=>x"c000",
---- 281=>x"c100", 282=>x"c000", 283=>x"c400", 284=>x"c000",
---- 285=>x"bf00", 286=>x"c000", 287=>x"c700", 288=>x"c400",
---- 289=>x"c500", 290=>x"bf00", 291=>x"c400", 292=>x"bc00",
---- 293=>x"c300", 294=>x"bf00", 295=>x"b700", 296=>x"bd00",
---- 297=>x"b900", 298=>x"bc00", 299=>x"b500", 300=>x"b900",
---- 301=>x"b500", 302=>x"b100", 303=>x"b100", 304=>x"b300",
---- 305=>x"b700", 306=>x"b900", 307=>x"ae00", 308=>x"b200",
---- 309=>x"b400", 310=>x"b400", 311=>x"b900", 312=>x"aa00",
---- 313=>x"b400", 314=>x"b700", 315=>x"b600", 316=>x"a700",
---- 317=>x"a700", 318=>x"b200", 319=>x"b700", 320=>x"a700",
---- 321=>x"a900", 322=>x"a700", 323=>x"b600", 324=>x"a300",
---- 325=>x"a600", 326=>x"a700", 327=>x"a500", 328=>x"a900",
---- 329=>x"9b00", 330=>x"9e00", 331=>x"6a00", 332=>x"a500",
---- 333=>x"9600", 334=>x"9500", 335=>x"5300", 336=>x"9600",
---- 337=>x"a300", 338=>x"b500", 339=>x"c500", 340=>x"a600",
---- 341=>x"c700", 342=>x"bf00", 343=>x"af00", 344=>x"c600",
---- 345=>x"b900", 346=>x"a800", 347=>x"aa00", 348=>x"ab00",
---- 349=>x"a500", 350=>x"ab00", 351=>x"c000", 352=>x"a000",
---- 353=>x"ac00", 354=>x"bd00", 355=>x"bd00", 356=>x"b200",
---- 357=>x"c500", 358=>x"c900", 359=>x"c200", 360=>x"c500",
---- 361=>x"c900", 362=>x"c800", 363=>x"c300", 364=>x"ca00",
---- 365=>x"c500", 366=>x"c400", 367=>x"c100", 368=>x"c600",
---- 369=>x"c500", 370=>x"c500", 371=>x"c200", 372=>x"3e00",
---- 373=>x"c400", 374=>x"c400", 375=>x"c000", 376=>x"bf00",
---- 377=>x"c200", 378=>x"c100", 379=>x"be00", 380=>x"bf00",
---- 381=>x"bf00", 382=>x"bc00", 383=>x"be00", 384=>x"bc00",
---- 385=>x"bc00", 386=>x"bc00", 387=>x"bd00", 388=>x"b800",
---- 389=>x"4600", 390=>x"b800", 391=>x"b900", 392=>x"b500",
---- 393=>x"b400", 394=>x"b300", 395=>x"b500", 396=>x"b500",
---- 397=>x"b300", 398=>x"b300", 399=>x"b300", 400=>x"b500",
---- 401=>x"af00", 402=>x"b000", 403=>x"b300", 404=>x"b000",
---- 405=>x"ad00", 406=>x"ac00", 407=>x"b400", 408=>x"aa00",
---- 409=>x"a700", 410=>x"ae00", 411=>x"b700", 412=>x"aa00",
---- 413=>x"ab00", 414=>x"b300", 415=>x"b800", 416=>x"b000",
---- 417=>x"5200", 418=>x"b500", 419=>x"b900", 420=>x"b000",
---- 421=>x"ac00", 422=>x"b300", 423=>x"b300", 424=>x"ae00",
---- 425=>x"b100", 426=>x"ab00", 427=>x"ac00", 428=>x"b000",
---- 429=>x"a700", 430=>x"a600", 431=>x"b800", 432=>x"a700",
---- 433=>x"ab00", 434=>x"bb00", 435=>x"c400", 436=>x"b200",
---- 437=>x"bb00", 438=>x"bd00", 439=>x"c300", 440=>x"b800",
---- 441=>x"b900", 442=>x"bc00", 443=>x"c500", 444=>x"b800",
---- 445=>x"bd00", 446=>x"c000", 447=>x"c400", 448=>x"b800",
---- 449=>x"c100", 450=>x"c300", 451=>x"c800", 452=>x"ba00",
---- 453=>x"bf00", 454=>x"c000", 455=>x"c500", 456=>x"bc00",
---- 457=>x"be00", 458=>x"c300", 459=>x"c600", 460=>x"c000",
---- 461=>x"c300", 462=>x"c300", 463=>x"c400", 464=>x"c100",
---- 465=>x"c300", 466=>x"c400", 467=>x"c500", 468=>x"c000",
---- 469=>x"c100", 470=>x"3d00", 471=>x"c600", 472=>x"bf00",
---- 473=>x"c300", 474=>x"c400", 475=>x"c400", 476=>x"be00",
---- 477=>x"bf00", 478=>x"c400", 479=>x"c600", 480=>x"bb00",
---- 481=>x"bd00", 482=>x"c100", 483=>x"c500", 484=>x"b700",
---- 485=>x"ba00", 486=>x"be00", 487=>x"c200", 488=>x"b500",
---- 489=>x"b800", 490=>x"bc00", 491=>x"c300", 492=>x"af00",
---- 493=>x"b700", 494=>x"b900", 495=>x"be00", 496=>x"ad00",
---- 497=>x"b000", 498=>x"b900", 499=>x"bf00", 500=>x"af00",
---- 501=>x"b100", 502=>x"b800", 503=>x"bd00", 504=>x"aa00",
---- 505=>x"b000", 506=>x"b500", 507=>x"bb00", 508=>x"a300",
---- 509=>x"aa00", 510=>x"b500", 511=>x"bb00", 512=>x"9f00",
---- 513=>x"5800", 514=>x"b200", 515=>x"c000", 516=>x"9d00",
---- 517=>x"a500", 518=>x"b200", 519=>x"be00", 520=>x"9d00",
---- 521=>x"a500", 522=>x"b300", 523=>x"be00", 524=>x"9a00",
---- 525=>x"a400", 526=>x"b300", 527=>x"bf00", 528=>x"9a00",
---- 529=>x"a300", 530=>x"ae00", 531=>x"c400", 532=>x"6700",
---- 533=>x"a500", 534=>x"b400", 535=>x"c800", 536=>x"9b00",
---- 537=>x"a700", 538=>x"b800", 539=>x"ca00", 540=>x"9d00",
---- 541=>x"a900", 542=>x"bc00", 543=>x"d400", 544=>x"9800",
---- 545=>x"ab00", 546=>x"c500", 547=>x"da00", 548=>x"9b00",
---- 549=>x"ad00", 550=>x"c400", 551=>x"db00", 552=>x"9600",
---- 553=>x"a800", 554=>x"c100", 555=>x"da00", 556=>x"9400",
---- 557=>x"a300", 558=>x"bb00", 559=>x"d900", 560=>x"9200",
---- 561=>x"a400", 562=>x"ba00", 563=>x"d600", 564=>x"8e00",
---- 565=>x"a500", 566=>x"bb00", 567=>x"d200", 568=>x"8e00",
---- 569=>x"a200", 570=>x"b600", 571=>x"cf00", 572=>x"8a00",
---- 573=>x"a200", 574=>x"b500", 575=>x"3100", 576=>x"8700",
---- 577=>x"9a00", 578=>x"b500", 579=>x"cc00", 580=>x"8300",
---- 581=>x"9800", 582=>x"b000", 583=>x"c900", 584=>x"8500",
---- 585=>x"9200", 586=>x"a900", 587=>x"c900", 588=>x"8100",
---- 589=>x"6e00", 590=>x"ab00", 591=>x"c800", 592=>x"8400",
---- 593=>x"9300", 594=>x"a400", 595=>x"c400", 596=>x"8600",
---- 597=>x"8f00", 598=>x"a300", 599=>x"c000", 600=>x"8600",
---- 601=>x"9100", 602=>x"a100", 603=>x"bc00", 604=>x"8400",
---- 605=>x"9000", 606=>x"9d00", 607=>x"b000", 608=>x"8600",
---- 609=>x"8c00", 610=>x"9800", 611=>x"ac00", 612=>x"8200",
---- 613=>x"8600", 614=>x"9900", 615=>x"af00", 616=>x"7e00",
---- 617=>x"8800", 618=>x"9800", 619=>x"ac00", 620=>x"7e00",
---- 621=>x"8800", 622=>x"9400", 623=>x"a400", 624=>x"7f00",
---- 625=>x"8600", 626=>x"9300", 627=>x"a200", 628=>x"7f00",
---- 629=>x"8700", 630=>x"9000", 631=>x"a100", 632=>x"7f00",
---- 633=>x"8700", 634=>x"8d00", 635=>x"a100", 636=>x"7900",
---- 637=>x"7c00", 638=>x"8a00", 639=>x"9e00", 640=>x"7900",
---- 641=>x"7600", 642=>x"8400", 643=>x"9600", 644=>x"7a00",
---- 645=>x"7b00", 646=>x"7d00", 647=>x"8500", 648=>x"5c00",
---- 649=>x"6d00", 650=>x"7900", 651=>x"7e00", 652=>x"6a00",
---- 653=>x"6500", 654=>x"7300", 655=>x"7700", 656=>x"7600",
---- 657=>x"7d00", 658=>x"8b00", 659=>x"9c00", 660=>x"8400",
---- 661=>x"9a00", 662=>x"bb00", 663=>x"c800", 664=>x"9a00",
---- 665=>x"a000", 666=>x"be00", 667=>x"c600", 668=>x"a900",
---- 669=>x"a600", 670=>x"bf00", 671=>x"c700", 672=>x"b500",
---- 673=>x"aa00", 674=>x"c200", 675=>x"c800", 676=>x"bd00",
---- 677=>x"ac00", 678=>x"c200", 679=>x"ce00", 680=>x"c000",
---- 681=>x"a900", 682=>x"b900", 683=>x"cd00", 684=>x"c300",
---- 685=>x"b200", 686=>x"c800", 687=>x"d200", 688=>x"c500",
---- 689=>x"cc00", 690=>x"c000", 691=>x"b400", 692=>x"9a00",
---- 693=>x"a600", 694=>x"9b00", 695=>x"9600", 696=>x"8900",
---- 697=>x"8d00", 698=>x"7800", 699=>x"6600", 700=>x"7c00",
---- 701=>x"7400", 702=>x"5b00", 703=>x"5200", 704=>x"8000",
---- 705=>x"8100", 706=>x"8300", 707=>x"7b00", 708=>x"b100",
---- 709=>x"b400", 710=>x"a200", 711=>x"8900", 712=>x"c800",
---- 713=>x"c400", 714=>x"a000", 715=>x"8700", 716=>x"a400",
---- 717=>x"a600", 718=>x"8f00", 719=>x"8700", 720=>x"8f00",
---- 721=>x"8e00", 722=>x"8400", 723=>x"8e00", 724=>x"8100",
---- 725=>x"8200", 726=>x"8d00", 727=>x"9700", 728=>x"8000",
---- 729=>x"9400", 730=>x"9a00", 731=>x"9300", 732=>x"9600",
---- 733=>x"9b00", 734=>x"9600", 735=>x"8c00", 736=>x"9800",
---- 737=>x"9900", 738=>x"8d00", 739=>x"8b00", 740=>x"9b00",
---- 741=>x"9600", 742=>x"9000", 743=>x"9000", 744=>x"9b00",
---- 745=>x"9600", 746=>x"9200", 747=>x"9500", 748=>x"9c00",
---- 749=>x"9600", 750=>x"9500", 751=>x"9800", 752=>x"9900",
---- 753=>x"9100", 754=>x"9800", 755=>x"6c00", 756=>x"9700",
---- 757=>x"9100", 758=>x"9900", 759=>x"8000", 760=>x"9400",
---- 761=>x"9400", 762=>x"9100", 763=>x"6f00", 764=>x"9400",
---- 765=>x"9100", 766=>x"8a00", 767=>x"6e00", 768=>x"8e00",
---- 769=>x"8900", 770=>x"8600", 771=>x"6100", 772=>x"8200",
---- 773=>x"8400", 774=>x"7d00", 775=>x"5500", 776=>x"9e00",
---- 777=>x"a300", 778=>x"9700", 779=>x"7100", 780=>x"4600",
---- 781=>x"bf00", 782=>x"c400", 783=>x"bd00", 784=>x"b300",
---- 785=>x"bf00", 786=>x"c300", 787=>x"c700", 788=>x"b700",
---- 789=>x"bf00", 790=>x"c400", 791=>x"c500", 792=>x"b700",
---- 793=>x"bf00", 794=>x"c300", 795=>x"c500", 796=>x"bb00",
---- 797=>x"bd00", 798=>x"c200", 799=>x"c400", 800=>x"bc00",
---- 801=>x"bf00", 802=>x"c100", 803=>x"c200", 804=>x"ba00",
---- 805=>x"bd00", 806=>x"be00", 807=>x"be00", 808=>x"b900",
---- 809=>x"bd00", 810=>x"be00", 811=>x"bd00", 812=>x"b900",
---- 813=>x"bd00", 814=>x"ba00", 815=>x"bc00", 816=>x"b400",
---- 817=>x"b700", 818=>x"b900", 819=>x"b900", 820=>x"b300",
---- 821=>x"b400", 822=>x"b500", 823=>x"b800", 824=>x"af00",
---- 825=>x"b000", 826=>x"b400", 827=>x"b300", 828=>x"af00",
---- 829=>x"ac00", 830=>x"af00", 831=>x"b100", 832=>x"ad00",
---- 833=>x"b000", 834=>x"ad00", 835=>x"b000", 836=>x"a800",
---- 837=>x"ae00", 838=>x"ad00", 839=>x"ae00", 840=>x"a900",
---- 841=>x"ac00", 842=>x"ad00", 843=>x"ad00", 844=>x"a500",
---- 845=>x"a800", 846=>x"aa00", 847=>x"ad00", 848=>x"a500",
---- 849=>x"a900", 850=>x"ab00", 851=>x"ad00", 852=>x"a400",
---- 853=>x"a700", 854=>x"ac00", 855=>x"ac00", 856=>x"a300",
---- 857=>x"a700", 858=>x"aa00", 859=>x"aa00", 860=>x"a600",
---- 861=>x"a600", 862=>x"a700", 863=>x"aa00", 864=>x"a300",
---- 865=>x"a600", 866=>x"a600", 867=>x"a800", 868=>x"a200",
---- 869=>x"a400", 870=>x"a400", 871=>x"a600", 872=>x"a100",
---- 873=>x"a300", 874=>x"a300", 875=>x"5900", 876=>x"9f00",
---- 877=>x"a100", 878=>x"a300", 879=>x"a500", 880=>x"9e00",
---- 881=>x"a100", 882=>x"a300", 883=>x"a400", 884=>x"9f00",
---- 885=>x"a000", 886=>x"a000", 887=>x"a300", 888=>x"9b00",
---- 889=>x"9f00", 890=>x"5f00", 891=>x"a200", 892=>x"9e00",
---- 893=>x"9c00", 894=>x"9d00", 895=>x"a100", 896=>x"9f00",
---- 897=>x"9e00", 898=>x"9d00", 899=>x"a100", 900=>x"6400",
---- 901=>x"9c00", 902=>x"a000", 903=>x"a300", 904=>x"9b00",
---- 905=>x"9c00", 906=>x"9f00", 907=>x"a100", 908=>x"9a00",
---- 909=>x"9b00", 910=>x"9d00", 911=>x"9e00", 912=>x"9800",
---- 913=>x"9a00", 914=>x"9b00", 915=>x"9f00", 916=>x"9800",
---- 917=>x"9800", 918=>x"9a00", 919=>x"9c00", 920=>x"9600",
---- 921=>x"9900", 922=>x"9900", 923=>x"9b00", 924=>x"9a00",
---- 925=>x"9a00", 926=>x"9900", 927=>x"9800", 928=>x"9500",
---- 929=>x"9700", 930=>x"9900", 931=>x"9d00", 932=>x"9300",
---- 933=>x"9800", 934=>x"9900", 935=>x"9b00", 936=>x"9400",
---- 937=>x"9600", 938=>x"9700", 939=>x"9700", 940=>x"9400",
---- 941=>x"9500", 942=>x"9600", 943=>x"9600", 944=>x"9500",
---- 945=>x"9700", 946=>x"9600", 947=>x"9900", 948=>x"9200",
---- 949=>x"9300", 950=>x"9400", 951=>x"9900", 952=>x"9100",
---- 953=>x"9200", 954=>x"9200", 955=>x"9400", 956=>x"9000",
---- 957=>x"9300", 958=>x"9100", 959=>x"9300", 960=>x"8f00",
---- 961=>x"9200", 962=>x"9100", 963=>x"9500", 964=>x"9100",
---- 965=>x"9000", 966=>x"9100", 967=>x"9300", 968=>x"9000",
---- 969=>x"9100", 970=>x"9000", 971=>x"9200", 972=>x"8d00",
---- 973=>x"8e00", 974=>x"8f00", 975=>x"9500", 976=>x"8a00",
---- 977=>x"8e00", 978=>x"9000", 979=>x"9000", 980=>x"8c00",
---- 981=>x"8d00", 982=>x"9100", 983=>x"8e00", 984=>x"8d00",
---- 985=>x"8d00", 986=>x"8e00", 987=>x"9000", 988=>x"8e00",
---- 989=>x"8c00", 990=>x"8f00", 991=>x"8d00", 992=>x"8d00",
---- 993=>x"8f00", 994=>x"9000", 995=>x"8e00", 996=>x"8e00",
---- 997=>x"9100", 998=>x"9100", 999=>x"9200", 1000=>x"8f00",
---- 1001=>x"9200", 1002=>x"9200", 1003=>x"9200", 1004=>x"9200",
---- 1005=>x"9300", 1006=>x"9200", 1007=>x"9000", 1008=>x"9300",
---- 1009=>x"9300", 1010=>x"9200", 1011=>x"9200", 1012=>x"9400",
---- 1013=>x"9400", 1014=>x"9100", 1015=>x"9200", 1016=>x"9300",
---- 1017=>x"9500", 1018=>x"9600", 1019=>x"9100", 1020=>x"9500",
---- 1021=>x"9600", 1022=>x"9700", 1023=>x"9300"),
----
---- 39 => (0=>x"7500", 1=>x"7100", 2=>x"7000", 3=>x"6600", 4=>x"7600",
---- 5=>x"7100", 6=>x"7000", 7=>x"6600", 8=>x"7300",
---- 9=>x"7200", 10=>x"6f00", 11=>x"6600", 12=>x"7300",
---- 13=>x"7100", 14=>x"6c00", 15=>x"6700", 16=>x"7400",
---- 17=>x"7000", 18=>x"6f00", 19=>x"6d00", 20=>x"7500",
---- 21=>x"7200", 22=>x"6f00", 23=>x"6b00", 24=>x"7500",
---- 25=>x"7100", 26=>x"6f00", 27=>x"6e00", 28=>x"7600",
---- 29=>x"7200", 30=>x"6e00", 31=>x"7300", 32=>x"7600",
---- 33=>x"7500", 34=>x"7200", 35=>x"7700", 36=>x"7400",
---- 37=>x"7200", 38=>x"7100", 39=>x"7200", 40=>x"8000",
---- 41=>x"7900", 42=>x"7100", 43=>x"7100", 44=>x"7900",
---- 45=>x"7800", 46=>x"7200", 47=>x"7100", 48=>x"7900",
---- 49=>x"7800", 50=>x"7300", 51=>x"6e00", 52=>x"7e00",
---- 53=>x"7d00", 54=>x"7400", 55=>x"6e00", 56=>x"7900",
---- 57=>x"7900", 58=>x"7700", 59=>x"7100", 60=>x"7400",
---- 61=>x"7700", 62=>x"7600", 63=>x"7400", 64=>x"7700",
---- 65=>x"7800", 66=>x"7300", 67=>x"7000", 68=>x"7a00",
---- 69=>x"7700", 70=>x"7400", 71=>x"6f00", 72=>x"7800",
---- 73=>x"7500", 74=>x"7700", 75=>x"7400", 76=>x"7800",
---- 77=>x"7500", 78=>x"7800", 79=>x"7900", 80=>x"7500",
---- 81=>x"8c00", 82=>x"7400", 83=>x"7300", 84=>x"7500",
---- 85=>x"7600", 86=>x"7300", 87=>x"7300", 88=>x"7600",
---- 89=>x"7700", 90=>x"6f00", 91=>x"7300", 92=>x"7500",
---- 93=>x"7300", 94=>x"7300", 95=>x"7100", 96=>x"7900",
---- 97=>x"7700", 98=>x"7200", 99=>x"7100", 100=>x"7800",
---- 101=>x"7800", 102=>x"7500", 103=>x"6f00", 104=>x"7500",
---- 105=>x"7500", 106=>x"7600", 107=>x"7100", 108=>x"8a00",
---- 109=>x"7000", 110=>x"7400", 111=>x"7000", 112=>x"7400",
---- 113=>x"7100", 114=>x"7300", 115=>x"6f00", 116=>x"7100",
---- 117=>x"7000", 118=>x"7000", 119=>x"6f00", 120=>x"7300",
---- 121=>x"7200", 122=>x"7000", 123=>x"6d00", 124=>x"7100",
---- 125=>x"7100", 126=>x"6d00", 127=>x"6b00", 128=>x"8f00",
---- 129=>x"7100", 130=>x"7000", 131=>x"6f00", 132=>x"7100",
---- 133=>x"6f00", 134=>x"6e00", 135=>x"6f00", 136=>x"6d00",
---- 137=>x"6d00", 138=>x"6e00", 139=>x"6a00", 140=>x"6f00",
---- 141=>x"6f00", 142=>x"6e00", 143=>x"6a00", 144=>x"6c00",
---- 145=>x"6a00", 146=>x"6a00", 147=>x"6c00", 148=>x"6b00",
---- 149=>x"6a00", 150=>x"6b00", 151=>x"6900", 152=>x"6a00",
---- 153=>x"6800", 154=>x"6700", 155=>x"6800", 156=>x"6500",
---- 157=>x"6400", 158=>x"6500", 159=>x"6800", 160=>x"6400",
---- 161=>x"6600", 162=>x"6400", 163=>x"6600", 164=>x"6700",
---- 165=>x"6500", 166=>x"6500", 167=>x"6400", 168=>x"6000",
---- 169=>x"6400", 170=>x"6200", 171=>x"6100", 172=>x"5d00",
---- 173=>x"6300", 174=>x"6100", 175=>x"6100", 176=>x"5900",
---- 177=>x"5e00", 178=>x"6200", 179=>x"6000", 180=>x"5500",
---- 181=>x"5800", 182=>x"5900", 183=>x"5c00", 184=>x"5000",
---- 185=>x"5100", 186=>x"5400", 187=>x"5700", 188=>x"4b00",
---- 189=>x"4a00", 190=>x"5000", 191=>x"5300", 192=>x"6700",
---- 193=>x"5000", 194=>x"4d00", 195=>x"4c00", 196=>x"cb00",
---- 197=>x"9000", 198=>x"4b00", 199=>x"4600", 200=>x"e600",
---- 201=>x"db00", 202=>x"9400", 203=>x"5f00", 204=>x"da00",
---- 205=>x"e200", 206=>x"df00", 207=>x"9600", 208=>x"d400",
---- 209=>x"da00", 210=>x"e100", 211=>x"d600", 212=>x"d800",
---- 213=>x"da00", 214=>x"d600", 215=>x"e000", 216=>x"d700",
---- 217=>x"dd00", 218=>x"dc00", 219=>x"dd00", 220=>x"d800",
---- 221=>x"d800", 222=>x"df00", 223=>x"e100", 224=>x"d500",
---- 225=>x"d300", 226=>x"d900", 227=>x"df00", 228=>x"d100",
---- 229=>x"d500", 230=>x"d700", 231=>x"df00", 232=>x"d100",
---- 233=>x"d200", 234=>x"d600", 235=>x"d800", 236=>x"d000",
---- 237=>x"d200", 238=>x"d200", 239=>x"d400", 240=>x"ca00",
---- 241=>x"cc00", 242=>x"cd00", 243=>x"d200", 244=>x"cd00",
---- 245=>x"cb00", 246=>x"d000", 247=>x"cf00", 248=>x"d100",
---- 249=>x"d200", 250=>x"d100", 251=>x"d100", 252=>x"cd00",
---- 253=>x"cc00", 254=>x"cb00", 255=>x"cc00", 256=>x"c900",
---- 257=>x"cb00", 258=>x"cc00", 259=>x"ce00", 260=>x"cd00",
---- 261=>x"ce00", 262=>x"c900", 263=>x"cc00", 264=>x"ca00",
---- 265=>x"c900", 266=>x"c900", 267=>x"c800", 268=>x"c900",
---- 269=>x"c800", 270=>x"cb00", 271=>x"c900", 272=>x"c800",
---- 273=>x"ca00", 274=>x"c900", 275=>x"c900", 276=>x"c300",
---- 277=>x"c800", 278=>x"c600", 279=>x"c700", 280=>x"c300",
---- 281=>x"c100", 282=>x"c500", 283=>x"c100", 284=>x"c700",
---- 285=>x"c000", 286=>x"ba00", 287=>x"c100", 288=>x"c300",
---- 289=>x"bc00", 290=>x"b600", 291=>x"bb00", 292=>x"bb00",
---- 293=>x"b800", 294=>x"b600", 295=>x"b900", 296=>x"af00",
---- 297=>x"b100", 298=>x"b800", 299=>x"ba00", 300=>x"b000",
---- 301=>x"ab00", 302=>x"b300", 303=>x"ba00", 304=>x"aa00",
---- 305=>x"b000", 306=>x"ac00", 307=>x"b500", 308=>x"b500",
---- 309=>x"ac00", 310=>x"b100", 311=>x"a800", 312=>x"b800",
---- 313=>x"ac00", 314=>x"aa00", 315=>x"a400", 316=>x"b100",
---- 317=>x"ac00", 318=>x"6100", 319=>x"a000", 320=>x"af00",
---- 321=>x"a500", 322=>x"9700", 323=>x"9800", 324=>x"a600",
---- 325=>x"9d00", 326=>x"a500", 327=>x"bc00", 328=>x"9900",
---- 329=>x"b400", 330=>x"c600", 331=>x"be00", 332=>x"bc00",
---- 333=>x"c400", 334=>x"b300", 335=>x"aa00", 336=>x"b800",
---- 337=>x"aa00", 338=>x"b600", 339=>x"b500", 340=>x"a800",
---- 341=>x"b100", 342=>x"c200", 343=>x"c300", 344=>x"bb00",
---- 345=>x"c100", 346=>x"c400", 347=>x"c900", 348=>x"ca00",
---- 349=>x"cd00", 350=>x"ca00", 351=>x"c600", 352=>x"c400",
---- 353=>x"c900", 354=>x"c700", 355=>x"c100", 356=>x"c400",
---- 357=>x"c600", 358=>x"c300", 359=>x"be00", 360=>x"c600",
---- 361=>x"c400", 362=>x"c100", 363=>x"c100", 364=>x"c100",
---- 365=>x"c000", 366=>x"c000", 367=>x"c100", 368=>x"c000",
---- 369=>x"c200", 370=>x"c000", 371=>x"c000", 372=>x"c100",
---- 373=>x"c200", 374=>x"be00", 375=>x"c000", 376=>x"be00",
---- 377=>x"3c00", 378=>x"bb00", 379=>x"b900", 380=>x"bf00",
---- 381=>x"bc00", 382=>x"ba00", 383=>x"bc00", 384=>x"bd00",
---- 385=>x"b900", 386=>x"bb00", 387=>x"bb00", 388=>x"bb00",
---- 389=>x"b600", 390=>x"b800", 391=>x"bc00", 392=>x"b500",
---- 393=>x"b700", 394=>x"b800", 395=>x"b900", 396=>x"af00",
---- 397=>x"b200", 398=>x"b900", 399=>x"bc00", 400=>x"ae00",
---- 401=>x"af00", 402=>x"b700", 403=>x"bf00", 404=>x"b700",
---- 405=>x"af00", 406=>x"b600", 407=>x"bd00", 408=>x"b400",
---- 409=>x"b400", 410=>x"b600", 411=>x"bd00", 412=>x"b600",
---- 413=>x"b600", 414=>x"ba00", 415=>x"ba00", 416=>x"4700",
---- 417=>x"b600", 418=>x"b800", 419=>x"b600", 420=>x"b300",
---- 421=>x"b400", 422=>x"bb00", 423=>x"bf00", 424=>x"b600",
---- 425=>x"c000", 426=>x"c600", 427=>x"c100", 428=>x"c200",
---- 429=>x"c400", 430=>x"c800", 431=>x"c300", 432=>x"c400",
---- 433=>x"c500", 434=>x"cb00", 435=>x"c500", 436=>x"c500",
---- 437=>x"c400", 438=>x"cc00", 439=>x"c800", 440=>x"c200",
---- 441=>x"3a00", 442=>x"c900", 443=>x"c800", 444=>x"c300",
---- 445=>x"c500", 446=>x"ca00", 447=>x"ca00", 448=>x"c600",
---- 449=>x"c700", 450=>x"cb00", 451=>x"ca00", 452=>x"c500",
---- 453=>x"c700", 454=>x"c900", 455=>x"c900", 456=>x"c800",
---- 457=>x"c600", 458=>x"c900", 459=>x"cb00", 460=>x"c800",
---- 461=>x"c900", 462=>x"c900", 463=>x"cd00", 464=>x"c400",
---- 465=>x"c900", 466=>x"cb00", 467=>x"cc00", 468=>x"c600",
---- 469=>x"c600", 470=>x"cc00", 471=>x"cc00", 472=>x"c800",
---- 473=>x"c700", 474=>x"c800", 475=>x"ca00", 476=>x"c500",
---- 477=>x"c600", 478=>x"c500", 479=>x"c500", 480=>x"c600",
---- 481=>x"c400", 482=>x"c200", 483=>x"c500", 484=>x"c500",
---- 485=>x"c300", 486=>x"c300", 487=>x"c400", 488=>x"c400",
---- 489=>x"c400", 490=>x"c200", 491=>x"bf00", 492=>x"c200",
---- 493=>x"c200", 494=>x"bd00", 495=>x"be00", 496=>x"c200",
---- 497=>x"c200", 498=>x"be00", 499=>x"4400", 500=>x"bf00",
---- 501=>x"c000", 502=>x"be00", 503=>x"ba00", 504=>x"c000",
---- 505=>x"bf00", 506=>x"bf00", 507=>x"bc00", 508=>x"c100",
---- 509=>x"c400", 510=>x"c100", 511=>x"bc00", 512=>x"c200",
---- 513=>x"c400", 514=>x"c300", 515=>x"be00", 516=>x"c200",
---- 517=>x"c300", 518=>x"c700", 519=>x"c600", 520=>x"c700",
---- 521=>x"ca00", 522=>x"cb00", 523=>x"c900", 524=>x"cc00",
---- 525=>x"cf00", 526=>x"cf00", 527=>x"cd00", 528=>x"d100",
---- 529=>x"d600", 530=>x"d700", 531=>x"af00", 532=>x"d700",
---- 533=>x"dc00", 534=>x"c700", 535=>x"7300", 536=>x"d700",
---- 537=>x"d900", 538=>x"a700", 539=>x"5a00", 540=>x"da00",
---- 541=>x"d500", 542=>x"8b00", 543=>x"6400", 544=>x"dd00",
---- 545=>x"cb00", 546=>x"7f00", 547=>x"5e00", 548=>x"df00",
---- 549=>x"c500", 550=>x"8800", 551=>x"6500", 552=>x"e000",
---- 553=>x"c700", 554=>x"aa00", 555=>x"a100", 556=>x"e000",
---- 557=>x"cc00", 558=>x"ab00", 559=>x"a200", 560=>x"e200",
---- 561=>x"d000", 562=>x"b200", 563=>x"9f00", 564=>x"df00",
---- 565=>x"d400", 566=>x"bb00", 567=>x"b000", 568=>x"de00",
---- 569=>x"d600", 570=>x"bf00", 571=>x"ba00", 572=>x"de00",
---- 573=>x"d700", 574=>x"c100", 575=>x"b800", 576=>x"db00",
---- 577=>x"db00", 578=>x"c300", 579=>x"b600", 580=>x"dc00",
---- 581=>x"de00", 582=>x"c900", 583=>x"b600", 584=>x"dd00",
---- 585=>x"dc00", 586=>x"cd00", 587=>x"b700", 588=>x"d900",
---- 589=>x"dc00", 590=>x"d000", 591=>x"ba00", 592=>x"dc00",
---- 593=>x"e000", 594=>x"d400", 595=>x"b800", 596=>x"d900",
---- 597=>x"df00", 598=>x"d500", 599=>x"b900", 600=>x"d600",
---- 601=>x"df00", 602=>x"d900", 603=>x"bc00", 604=>x"cd00",
---- 605=>x"df00", 606=>x"dc00", 607=>x"be00", 608=>x"ca00",
---- 609=>x"dd00", 610=>x"dc00", 611=>x"c400", 612=>x"c900",
---- 613=>x"db00", 614=>x"df00", 615=>x"cb00", 616=>x"c200",
---- 617=>x"d500", 618=>x"e300", 619=>x"d600", 620=>x"b800",
---- 621=>x"d400", 622=>x"e500", 623=>x"dd00", 624=>x"b200",
---- 625=>x"d200", 626=>x"e400", 627=>x"df00", 628=>x"ae00",
---- 629=>x"cc00", 630=>x"e600", 631=>x"1d00", 632=>x"b300",
---- 633=>x"cb00", 634=>x"e700", 635=>x"e300", 636=>x"b500",
---- 637=>x"c800", 638=>x"dd00", 639=>x"e000", 640=>x"ac00",
---- 641=>x"c500", 642=>x"cf00", 643=>x"d400", 644=>x"a100",
---- 645=>x"bc00", 646=>x"cc00", 647=>x"bc00", 648=>x"9300",
---- 649=>x"b100", 650=>x"c300", 651=>x"ac00", 652=>x"8900",
---- 653=>x"b200", 654=>x"b800", 655=>x"aa00", 656=>x"b100",
---- 657=>x"be00", 658=>x"b300", 659=>x"a600", 660=>x"c400",
---- 661=>x"be00", 662=>x"b000", 663=>x"a700", 664=>x"c000",
---- 665=>x"bf00", 666=>x"b300", 667=>x"a600", 668=>x"c000",
---- 669=>x"c100", 670=>x"b200", 671=>x"a200", 672=>x"c500",
---- 673=>x"c500", 674=>x"b100", 675=>x"a000", 676=>x"c500",
---- 677=>x"c000", 678=>x"af00", 679=>x"a000", 680=>x"c700",
---- 681=>x"be00", 682=>x"b000", 683=>x"9b00", 684=>x"cb00",
---- 685=>x"c300", 686=>x"b400", 687=>x"9800", 688=>x"ac00",
---- 689=>x"b500", 690=>x"b400", 691=>x"9300", 692=>x"9200",
---- 693=>x"9b00", 694=>x"9900", 695=>x"7b00", 696=>x"7200",
---- 697=>x"7900", 698=>x"6a00", 699=>x"6000", 700=>x"5f00",
---- 701=>x"6f00", 702=>x"7000", 703=>x"7300", 704=>x"7900",
---- 705=>x"8700", 706=>x"8500", 707=>x"8500", 708=>x"8600",
---- 709=>x"8d00", 710=>x"9000", 711=>x"9000", 712=>x"8800",
---- 713=>x"8f00", 714=>x"9500", 715=>x"8f00", 716=>x"9000",
---- 717=>x"9300", 718=>x"9700", 719=>x"8e00", 720=>x"9300",
---- 721=>x"9700", 722=>x"8f00", 723=>x"8b00", 724=>x"9300",
---- 725=>x"9300", 726=>x"8d00", 727=>x"7900", 728=>x"8f00",
---- 729=>x"9000", 730=>x"8000", 731=>x"4e00", 732=>x"8d00",
---- 733=>x"9100", 734=>x"5c00", 735=>x"3c00", 736=>x"9000",
---- 737=>x"8200", 738=>x"3500", 739=>x"3f00", 740=>x"9200",
---- 741=>x"5c00", 742=>x"d700", 743=>x"4800", 744=>x"8600",
---- 745=>x"3300", 746=>x"2800", 747=>x"4000", 748=>x"6c00",
---- 749=>x"2500", 750=>x"3100", 751=>x"4400", 752=>x"4c00",
---- 753=>x"2500", 754=>x"3a00", 755=>x"4500", 756=>x"3700",
---- 757=>x"2700", 758=>x"3e00", 759=>x"3c00", 760=>x"3200",
---- 761=>x"2900", 762=>x"3f00", 763=>x"3500", 764=>x"3500",
---- 765=>x"2b00", 766=>x"3d00", 767=>x"3700", 768=>x"3300",
---- 769=>x"2e00", 770=>x"3700", 771=>x"3700", 772=>x"3200",
---- 773=>x"3200", 774=>x"3400", 775=>x"3600", 776=>x"4400",
---- 777=>x"3900", 778=>x"3300", 779=>x"3800", 780=>x"a900",
---- 781=>x"8900", 782=>x"a100", 783=>x"4100", 784=>x"cc00",
---- 785=>x"cb00", 786=>x"c000", 787=>x"a000", 788=>x"c600",
---- 789=>x"c800", 790=>x"cd00", 791=>x"d000", 792=>x"c800",
---- 793=>x"c800", 794=>x"c900", 795=>x"c900", 796=>x"c800",
---- 797=>x"c700", 798=>x"c900", 799=>x"c800", 800=>x"c300",
---- 801=>x"c400", 802=>x"c900", 803=>x"c800", 804=>x"be00",
---- 805=>x"c100", 806=>x"c500", 807=>x"c500", 808=>x"bd00",
---- 809=>x"c200", 810=>x"c300", 811=>x"c200", 812=>x"4100",
---- 813=>x"c000", 814=>x"c000", 815=>x"c100", 816=>x"be00",
---- 817=>x"be00", 818=>x"be00", 819=>x"bd00", 820=>x"ba00",
---- 821=>x"bb00", 822=>x"bd00", 823=>x"bf00", 824=>x"b400",
---- 825=>x"bb00", 826=>x"bd00", 827=>x"bd00", 828=>x"b300",
---- 829=>x"b500", 830=>x"b900", 831=>x"b800", 832=>x"b300",
---- 833=>x"b500", 834=>x"b700", 835=>x"b600", 836=>x"b300",
---- 837=>x"b400", 838=>x"b500", 839=>x"ba00", 840=>x"b200",
---- 841=>x"b100", 842=>x"b500", 843=>x"b900", 844=>x"b100",
---- 845=>x"b200", 846=>x"b700", 847=>x"b700", 848=>x"af00",
---- 849=>x"b200", 850=>x"b600", 851=>x"b300", 852=>x"af00",
---- 853=>x"b200", 854=>x"b100", 855=>x"b500", 856=>x"af00",
---- 857=>x"af00", 858=>x"b000", 859=>x"b900", 860=>x"ab00",
---- 861=>x"af00", 862=>x"b200", 863=>x"b300", 864=>x"ac00",
---- 865=>x"ad00", 866=>x"4f00", 867=>x"b400", 868=>x"ab00",
---- 869=>x"b000", 870=>x"af00", 871=>x"b100", 872=>x"ab00",
---- 873=>x"b000", 874=>x"ac00", 875=>x"b100", 876=>x"a700",
---- 877=>x"ac00", 878=>x"af00", 879=>x"b200", 880=>x"a800",
---- 881=>x"ab00", 882=>x"b100", 883=>x"b200", 884=>x"a500",
---- 885=>x"a900", 886=>x"aa00", 887=>x"ac00", 888=>x"a600",
---- 889=>x"aa00", 890=>x"a800", 891=>x"a900", 892=>x"a700",
---- 893=>x"a700", 894=>x"a900", 895=>x"aa00", 896=>x"a400",
---- 897=>x"a700", 898=>x"a700", 899=>x"ad00", 900=>x"a400",
---- 901=>x"a700", 902=>x"a500", 903=>x"a900", 904=>x"a400",
---- 905=>x"a600", 906=>x"a700", 907=>x"a500", 908=>x"a100",
---- 909=>x"a500", 910=>x"a400", 911=>x"a600", 912=>x"9c00",
---- 913=>x"a200", 914=>x"a300", 915=>x"a500", 916=>x"9d00",
---- 917=>x"9f00", 918=>x"a000", 919=>x"a500", 920=>x"9d00",
---- 921=>x"a100", 922=>x"a300", 923=>x"a500", 924=>x"a000",
---- 925=>x"a200", 926=>x"a100", 927=>x"a400", 928=>x"9d00",
---- 929=>x"9f00", 930=>x"a000", 931=>x"a300", 932=>x"6300",
---- 933=>x"9f00", 934=>x"6000", 935=>x"a200", 936=>x"9a00",
---- 937=>x"9f00", 938=>x"a000", 939=>x"a100", 940=>x"9900",
---- 941=>x"9b00", 942=>x"9e00", 943=>x"9d00", 944=>x"9c00",
---- 945=>x"9b00", 946=>x"9c00", 947=>x"9f00", 948=>x"9a00",
---- 949=>x"6400", 950=>x"9d00", 951=>x"9d00", 952=>x"9a00",
---- 953=>x"9b00", 954=>x"9d00", 955=>x"9b00", 956=>x"9800",
---- 957=>x"6600", 958=>x"9b00", 959=>x"9b00", 960=>x"9800",
---- 961=>x"9700", 962=>x"9800", 963=>x"9c00", 964=>x"9400",
---- 965=>x"9500", 966=>x"9700", 967=>x"9a00", 968=>x"9400",
---- 969=>x"9300", 970=>x"9800", 971=>x"9a00", 972=>x"9400",
---- 973=>x"9200", 974=>x"9500", 975=>x"9a00", 976=>x"9400",
---- 977=>x"9300", 978=>x"9600", 979=>x"9700", 980=>x"9100",
---- 981=>x"9600", 982=>x"9500", 983=>x"9700", 984=>x"9100",
---- 985=>x"9300", 986=>x"9500", 987=>x"9600", 988=>x"9100",
---- 989=>x"9500", 990=>x"9700", 991=>x"9700", 992=>x"9100",
---- 993=>x"9300", 994=>x"9400", 995=>x"9400", 996=>x"9300",
---- 997=>x"9400", 998=>x"9200", 999=>x"9700", 1000=>x"9300",
---- 1001=>x"9400", 1002=>x"9400", 1003=>x"6900", 1004=>x"9500",
---- 1005=>x"9500", 1006=>x"9400", 1007=>x"9600", 1008=>x"9300",
---- 1009=>x"9700", 1010=>x"9600", 1011=>x"9b00", 1012=>x"9300",
---- 1013=>x"9600", 1014=>x"9600", 1015=>x"9b00", 1016=>x"9400",
---- 1017=>x"9600", 1018=>x"9500", 1019=>x"9500", 1020=>x"9700",
---- 1021=>x"9600", 1022=>x"9700", 1023=>x"9600"),
----
---- 40 => (0=>x"6900", 1=>x"7400", 2=>x"7b00", 3=>x"8800", 4=>x"6900",
---- 5=>x"7400", 6=>x"7b00", 7=>x"8800", 8=>x"6900",
---- 9=>x"7300", 10=>x"7c00", 11=>x"8600", 12=>x"6500",
---- 13=>x"6f00", 14=>x"7b00", 15=>x"8000", 16=>x"6500",
---- 17=>x"6a00", 18=>x"7200", 19=>x"7b00", 20=>x"6b00",
---- 21=>x"6700", 22=>x"6c00", 23=>x"7400", 24=>x"6d00",
---- 25=>x"6a00", 26=>x"6600", 27=>x"9000", 28=>x"6e00",
---- 29=>x"6b00", 30=>x"6600", 31=>x"6c00", 32=>x"6e00",
---- 33=>x"6b00", 34=>x"6a00", 35=>x"6900", 36=>x"6f00",
---- 37=>x"6f00", 38=>x"6800", 39=>x"6500", 40=>x"6e00",
---- 41=>x"6b00", 42=>x"6c00", 43=>x"6700", 44=>x"6e00",
---- 45=>x"6f00", 46=>x"6a00", 47=>x"6800", 48=>x"6e00",
---- 49=>x"6d00", 50=>x"6a00", 51=>x"6a00", 52=>x"6e00",
---- 53=>x"6d00", 54=>x"6a00", 55=>x"6900", 56=>x"7000",
---- 57=>x"6f00", 58=>x"6b00", 59=>x"6a00", 60=>x"7000",
---- 61=>x"7000", 62=>x"6e00", 63=>x"6c00", 64=>x"9200",
---- 65=>x"6e00", 66=>x"6c00", 67=>x"6b00", 68=>x"6f00",
---- 69=>x"7200", 70=>x"6c00", 71=>x"6b00", 72=>x"7200",
---- 73=>x"7200", 74=>x"6e00", 75=>x"6b00", 76=>x"7400",
---- 77=>x"6f00", 78=>x"6c00", 79=>x"6900", 80=>x"7100",
---- 81=>x"7300", 82=>x"7000", 83=>x"6e00", 84=>x"8d00",
---- 85=>x"7300", 86=>x"6f00", 87=>x"6d00", 88=>x"7400",
---- 89=>x"7000", 90=>x"6d00", 91=>x"6a00", 92=>x"7500",
---- 93=>x"6f00", 94=>x"6e00", 95=>x"6900", 96=>x"7200",
---- 97=>x"7200", 98=>x"6e00", 99=>x"6c00", 100=>x"7000",
---- 101=>x"9100", 102=>x"6d00", 103=>x"6b00", 104=>x"7100",
---- 105=>x"6f00", 106=>x"6c00", 107=>x"6900", 108=>x"7000",
---- 109=>x"7400", 110=>x"6e00", 111=>x"6700", 112=>x"7200",
---- 113=>x"6d00", 114=>x"6f00", 115=>x"6a00", 116=>x"6d00",
---- 117=>x"6b00", 118=>x"6900", 119=>x"6b00", 120=>x"6c00",
---- 121=>x"6b00", 122=>x"6700", 123=>x"6600", 124=>x"6c00",
---- 125=>x"6900", 126=>x"6900", 127=>x"6300", 128=>x"6a00",
---- 129=>x"6a00", 130=>x"6900", 131=>x"6500", 132=>x"9400",
---- 133=>x"6a00", 134=>x"6500", 135=>x"6500", 136=>x"6b00",
---- 137=>x"6a00", 138=>x"6900", 139=>x"6500", 140=>x"6a00",
---- 141=>x"6c00", 142=>x"6900", 143=>x"6400", 144=>x"6f00",
---- 145=>x"6d00", 146=>x"9600", 147=>x"9800", 148=>x"6b00",
---- 149=>x"6a00", 150=>x"6600", 151=>x"6400", 152=>x"6a00",
---- 153=>x"6900", 154=>x"6700", 155=>x"6300", 156=>x"6800",
---- 157=>x"9900", 158=>x"6700", 159=>x"6200", 160=>x"6500",
---- 161=>x"6600", 162=>x"6400", 163=>x"6100", 164=>x"6500",
---- 165=>x"6400", 166=>x"6500", 167=>x"5e00", 168=>x"6200",
---- 169=>x"6100", 170=>x"6200", 171=>x"6000", 172=>x"6700",
---- 173=>x"6000", 174=>x"6000", 175=>x"5e00", 176=>x"6000",
---- 177=>x"5e00", 178=>x"6000", 179=>x"5e00", 180=>x"6000",
---- 181=>x"a000", 182=>x"5f00", 183=>x"5e00", 184=>x"5800",
---- 185=>x"5800", 186=>x"5b00", 187=>x"5a00", 188=>x"5400",
---- 189=>x"5800", 190=>x"5a00", 191=>x"5800", 192=>x"4f00",
---- 193=>x"5400", 194=>x"5700", 195=>x"5700", 196=>x"4900",
---- 197=>x"4d00", 198=>x"5500", 199=>x"5400", 200=>x"4500",
---- 201=>x"4900", 202=>x"4f00", 203=>x"5100", 204=>x"4300",
---- 205=>x"4200", 206=>x"4700", 207=>x"4d00", 208=>x"7500",
---- 209=>x"3200", 210=>x"4000", 211=>x"4800", 212=>x"c200",
---- 213=>x"4d00", 214=>x"3900", 215=>x"4500", 216=>x"dc00",
---- 217=>x"8000", 218=>x"4d00", 219=>x"4600", 220=>x"e300",
---- 221=>x"cb00", 222=>x"8900", 223=>x"3900", 224=>x"e200",
---- 225=>x"e600", 226=>x"c100", 227=>x"4a00", 228=>x"1e00",
---- 229=>x"1d00", 230=>x"e200", 231=>x"7500", 232=>x"e100",
---- 233=>x"de00", 234=>x"e300", 235=>x"a400", 236=>x"da00",
---- 237=>x"e100", 238=>x"e100", 239=>x"cc00", 240=>x"d600",
---- 241=>x"dd00", 242=>x"e100", 243=>x"df00", 244=>x"d000",
---- 245=>x"d900", 246=>x"e000", 247=>x"e000", 248=>x"cd00",
---- 249=>x"d300", 250=>x"da00", 251=>x"de00", 252=>x"cd00",
---- 253=>x"d000", 254=>x"d100", 255=>x"d600", 256=>x"ce00",
---- 257=>x"cf00", 258=>x"cf00", 259=>x"d300", 260=>x"ce00",
---- 261=>x"ce00", 262=>x"cf00", 263=>x"cf00", 264=>x"ca00",
---- 265=>x"cd00", 266=>x"cb00", 267=>x"cb00", 268=>x"c800",
---- 269=>x"c600", 270=>x"c400", 271=>x"c700", 272=>x"c800",
---- 273=>x"c600", 274=>x"c500", 275=>x"c200", 276=>x"c800",
---- 277=>x"c900", 278=>x"c600", 279=>x"c400", 280=>x"c000",
---- 281=>x"c400", 282=>x"c400", 283=>x"c500", 284=>x"bd00",
---- 285=>x"bc00", 286=>x"c100", 287=>x"c200", 288=>x"be00",
---- 289=>x"bf00", 290=>x"bb00", 291=>x"be00", 292=>x"bb00",
---- 293=>x"bc00", 294=>x"b700", 295=>x"4600", 296=>x"ba00",
---- 297=>x"b300", 298=>x"b900", 299=>x"4900", 300=>x"b900",
---- 301=>x"b600", 302=>x"b000", 303=>x"b300", 304=>x"b900",
---- 305=>x"b800", 306=>x"aa00", 307=>x"ae00", 308=>x"b500",
---- 309=>x"b300", 310=>x"a700", 311=>x"a000", 312=>x"ab00",
---- 313=>x"a800", 314=>x"9c00", 315=>x"a400", 316=>x"9800",
---- 317=>x"a600", 318=>x"b700", 319=>x"c700", 320=>x"aa00",
---- 321=>x"c600", 322=>x"c500", 323=>x"b500", 324=>x"c800",
---- 325=>x"b700", 326=>x"a900", 327=>x"b200", 328=>x"af00",
---- 329=>x"af00", 330=>x"b500", 331=>x"bf00", 332=>x"b200",
---- 333=>x"bc00", 334=>x"c200", 335=>x"c600", 336=>x"ba00",
---- 337=>x"ca00", 338=>x"cd00", 339=>x"c800", 340=>x"c100",
---- 341=>x"cc00", 342=>x"c800", 343=>x"bf00", 344=>x"c500",
---- 345=>x"c600", 346=>x"c200", 347=>x"bc00", 348=>x"c100",
---- 349=>x"c500", 350=>x"c200", 351=>x"c100", 352=>x"3f00",
---- 353=>x"c300", 354=>x"c300", 355=>x"c300", 356=>x"c200",
---- 357=>x"c500", 358=>x"c500", 359=>x"c100", 360=>x"c300",
---- 361=>x"c500", 362=>x"c300", 363=>x"c100", 364=>x"c200",
---- 365=>x"c100", 366=>x"c300", 367=>x"c300", 368=>x"c300",
---- 369=>x"c500", 370=>x"c200", 371=>x"c200", 372=>x"4000",
---- 373=>x"c100", 374=>x"c300", 375=>x"c300", 376=>x"be00",
---- 377=>x"3e00", 378=>x"be00", 379=>x"be00", 380=>x"be00",
---- 381=>x"bd00", 382=>x"bf00", 383=>x"be00", 384=>x"bb00",
---- 385=>x"be00", 386=>x"c000", 387=>x"be00", 388=>x"4400",
---- 389=>x"be00", 390=>x"bf00", 391=>x"be00", 392=>x"bd00",
---- 393=>x"bf00", 394=>x"c100", 395=>x"bf00", 396=>x"bd00",
---- 397=>x"bd00", 398=>x"be00", 399=>x"bd00", 400=>x"bd00",
---- 401=>x"c100", 402=>x"c000", 403=>x"bd00", 404=>x"c000",
---- 405=>x"c000", 406=>x"c100", 407=>x"bf00", 408=>x"bc00",
---- 409=>x"bc00", 410=>x"b900", 411=>x"b600", 412=>x"b700",
---- 413=>x"b600", 414=>x"b300", 415=>x"b900", 416=>x"ba00",
---- 417=>x"ba00", 418=>x"bc00", 419=>x"c100", 420=>x"c000",
---- 421=>x"c100", 422=>x"c200", 423=>x"c300", 424=>x"c100",
---- 425=>x"3f00", 426=>x"c300", 427=>x"c500", 428=>x"c300",
---- 429=>x"3b00", 430=>x"c500", 431=>x"c600", 432=>x"c500",
---- 433=>x"c400", 434=>x"c600", 435=>x"c400", 436=>x"c700",
---- 437=>x"c400", 438=>x"c400", 439=>x"c700", 440=>x"c800",
---- 441=>x"c700", 442=>x"c900", 443=>x"c900", 444=>x"c800",
---- 445=>x"3600", 446=>x"cc00", 447=>x"cc00", 448=>x"c700",
---- 449=>x"c800", 450=>x"cb00", 451=>x"ce00", 452=>x"c900",
---- 453=>x"c900", 454=>x"ce00", 455=>x"d000", 456=>x"ca00",
---- 457=>x"cb00", 458=>x"d000", 459=>x"d200", 460=>x"cb00",
---- 461=>x"cb00", 462=>x"ce00", 463=>x"d100", 464=>x"cc00",
---- 465=>x"cc00", 466=>x"d000", 467=>x"cf00", 468=>x"cb00",
---- 469=>x"cd00", 470=>x"ce00", 471=>x"d000", 472=>x"cb00",
---- 473=>x"cc00", 474=>x"cc00", 475=>x"cf00", 476=>x"c900",
---- 477=>x"ca00", 478=>x"cd00", 479=>x"cc00", 480=>x"c800",
---- 481=>x"c900", 482=>x"ca00", 483=>x"cb00", 484=>x"c600",
---- 485=>x"c600", 486=>x"c900", 487=>x"cc00", 488=>x"c300",
---- 489=>x"c500", 490=>x"c800", 491=>x"c900", 492=>x"c000",
---- 493=>x"c100", 494=>x"c400", 495=>x"c800", 496=>x"bd00",
---- 497=>x"c000", 498=>x"c300", 499=>x"c700", 500=>x"c300",
---- 501=>x"c100", 502=>x"be00", 503=>x"c200", 504=>x"c100",
---- 505=>x"bf00", 506=>x"b900", 507=>x"bb00", 508=>x"be00",
---- 509=>x"ba00", 510=>x"b000", 511=>x"a700", 512=>x"bf00",
---- 513=>x"bd00", 514=>x"aa00", 515=>x"9300", 516=>x"bf00",
---- 517=>x"b800", 518=>x"9b00", 519=>x"7500", 520=>x"be00",
---- 521=>x"9900", 522=>x"6000", 523=>x"4000", 524=>x"9a00",
---- 525=>x"4500", 526=>x"3200", 527=>x"3000", 528=>x"5000",
---- 529=>x"2c00", 530=>x"3100", 531=>x"2c00", 532=>x"4000",
---- 533=>x"3600", 534=>x"4400", 535=>x"3400", 536=>x"6200",
---- 537=>x"4500", 538=>x"5300", 539=>x"5800", 540=>x"8400",
---- 541=>x"7500", 542=>x"4900", 543=>x"5d00", 544=>x"7800",
---- 545=>x"9100", 546=>x"7400", 547=>x"5900", 548=>x"6100",
---- 549=>x"7700", 550=>x"8c00", 551=>x"8c00", 552=>x"9500",
---- 553=>x"8600", 554=>x"9100", 555=>x"8f00", 556=>x"9800",
---- 557=>x"9000", 558=>x"8f00", 559=>x"7d00", 560=>x"9500",
---- 561=>x"8d00", 562=>x"8500", 563=>x"8000", 564=>x"a300",
---- 565=>x"9d00", 566=>x"9100", 567=>x"8c00", 568=>x"aa00",
---- 569=>x"a000", 570=>x"9c00", 571=>x"9700", 572=>x"b000",
---- 573=>x"a100", 574=>x"9e00", 575=>x"9a00", 576=>x"b500",
---- 577=>x"5500", 578=>x"9f00", 579=>x"9900", 580=>x"af00",
---- 581=>x"ad00", 582=>x"a400", 583=>x"9700", 584=>x"aa00",
---- 585=>x"a800", 586=>x"a500", 587=>x"9e00", 588=>x"aa00",
---- 589=>x"a400", 590=>x"a200", 591=>x"a000", 592=>x"a900",
---- 593=>x"a300", 594=>x"a100", 595=>x"9f00", 596=>x"a900",
---- 597=>x"a400", 598=>x"a400", 599=>x"9e00", 600=>x"a700",
---- 601=>x"a800", 602=>x"a300", 603=>x"9e00", 604=>x"a500",
---- 605=>x"a400", 606=>x"9f00", 607=>x"9a00", 608=>x"a100",
---- 609=>x"a000", 610=>x"a000", 611=>x"9b00", 612=>x"a400",
---- 613=>x"a400", 614=>x"9e00", 615=>x"9b00", 616=>x"a500",
---- 617=>x"9f00", 618=>x"9c00", 619=>x"9800", 620=>x"ab00",
---- 621=>x"9b00", 622=>x"9b00", 623=>x"9800", 624=>x"b300",
---- 625=>x"9900", 626=>x"9d00", 627=>x"9600", 628=>x"ba00",
---- 629=>x"9300", 630=>x"6800", 631=>x"9700", 632=>x"bb00",
---- 633=>x"8e00", 634=>x"9300", 635=>x"9500", 636=>x"b700",
---- 637=>x"8d00", 638=>x"9700", 639=>x"6c00", 640=>x"a800",
---- 641=>x"8f00", 642=>x"9400", 643=>x"9400", 644=>x"9900",
---- 645=>x"9400", 646=>x"9300", 647=>x"9600", 648=>x"a100",
---- 649=>x"9700", 650=>x"9200", 651=>x"9200", 652=>x"a200",
---- 653=>x"9900", 654=>x"9400", 655=>x"8e00", 656=>x"9e00",
---- 657=>x"9900", 658=>x"9500", 659=>x"8f00", 660=>x"9b00",
---- 661=>x"9600", 662=>x"9500", 663=>x"8f00", 664=>x"9a00",
---- 665=>x"9700", 666=>x"9100", 667=>x"8d00", 668=>x"9900",
---- 669=>x"9100", 670=>x"9200", 671=>x"8e00", 672=>x"9700",
---- 673=>x"9000", 674=>x"9200", 675=>x"8c00", 676=>x"9400",
---- 677=>x"9000", 678=>x"9000", 679=>x"8a00", 680=>x"8d00",
---- 681=>x"9200", 682=>x"8d00", 683=>x"8800", 684=>x"8d00",
---- 685=>x"8e00", 686=>x"8b00", 687=>x"8a00", 688=>x"8300",
---- 689=>x"8600", 690=>x"8a00", 691=>x"8d00", 692=>x"7700",
---- 693=>x"7900", 694=>x"8c00", 695=>x"8c00", 696=>x"7800",
---- 697=>x"8e00", 698=>x"9000", 699=>x"7e00", 700=>x"8700",
---- 701=>x"9000", 702=>x"9300", 703=>x"5d00", 704=>x"9100",
---- 705=>x"9200", 706=>x"8100", 707=>x"3700", 708=>x"9000",
---- 709=>x"8c00", 710=>x"ad00", 711=>x"2800", 712=>x"8c00",
---- 713=>x"7000", 714=>x"3100", 715=>x"2c00", 716=>x"8800",
---- 717=>x"4400", 718=>x"2800", 719=>x"2d00", 720=>x"6900",
---- 721=>x"2e00", 722=>x"2e00", 723=>x"2f00", 724=>x"4d00",
---- 725=>x"2900", 726=>x"2f00", 727=>x"3000", 728=>x"4100",
---- 729=>x"2a00", 730=>x"2c00", 731=>x"2900", 732=>x"4100",
---- 733=>x"2900", 734=>x"2e00", 735=>x"2b00", 736=>x"3e00",
---- 737=>x"2e00", 738=>x"2c00", 739=>x"2d00", 740=>x"3800",
---- 741=>x"2a00", 742=>x"2b00", 743=>x"2e00", 744=>x"3000",
---- 745=>x"2b00", 746=>x"2e00", 747=>x"3100", 748=>x"2d00",
---- 749=>x"2c00", 750=>x"3000", 751=>x"3000", 752=>x"2b00",
---- 753=>x"3100", 754=>x"3400", 755=>x"2f00", 756=>x"3000",
---- 757=>x"3500", 758=>x"3500", 759=>x"3200", 760=>x"3500",
---- 761=>x"3900", 762=>x"3800", 763=>x"3600", 764=>x"3800",
---- 765=>x"3b00", 766=>x"3a00", 767=>x"3900", 768=>x"3800",
---- 769=>x"3500", 770=>x"3700", 771=>x"3900", 772=>x"3900",
---- 773=>x"3800", 774=>x"3700", 775=>x"3a00", 776=>x"3f00",
---- 777=>x"3c00", 778=>x"3900", 779=>x"3700", 780=>x"3300",
---- 781=>x"3200", 782=>x"3600", 783=>x"3800", 784=>x"6a00",
---- 785=>x"4400", 786=>x"3500", 787=>x"3700", 788=>x"c900",
---- 789=>x"a700", 790=>x"7700", 791=>x"4b00", 792=>x"cb00",
---- 793=>x"cf00", 794=>x"c900", 795=>x"ae00", 796=>x"ca00",
---- 797=>x"c800", 798=>x"cb00", 799=>x"d300", 800=>x"ca00",
---- 801=>x"cb00", 802=>x"3500", 803=>x"cb00", 804=>x"c800",
---- 805=>x"cb00", 806=>x"cb00", 807=>x"cc00", 808=>x"c600",
---- 809=>x"c700", 810=>x"ca00", 811=>x"cc00", 812=>x"c300",
---- 813=>x"c700", 814=>x"c900", 815=>x"cc00", 816=>x"c200",
---- 817=>x"c500", 818=>x"c600", 819=>x"c900", 820=>x"c200",
---- 821=>x"c400", 822=>x"3a00", 823=>x"c700", 824=>x"c000",
---- 825=>x"c100", 826=>x"c100", 827=>x"c700", 828=>x"bc00",
---- 829=>x"c000", 830=>x"c400", 831=>x"c700", 832=>x"b900",
---- 833=>x"c000", 834=>x"c200", 835=>x"c400", 836=>x"ba00",
---- 837=>x"bf00", 838=>x"bf00", 839=>x"c400", 840=>x"b900",
---- 841=>x"be00", 842=>x"bf00", 843=>x"c400", 844=>x"b700",
---- 845=>x"c000", 846=>x"c000", 847=>x"c000", 848=>x"b800",
---- 849=>x"ba00", 850=>x"bd00", 851=>x"c000", 852=>x"b900",
---- 853=>x"bb00", 854=>x"bd00", 855=>x"be00", 856=>x"ba00",
---- 857=>x"ba00", 858=>x"bb00", 859=>x"bb00", 860=>x"b700",
---- 861=>x"bb00", 862=>x"bc00", 863=>x"bd00", 864=>x"b400",
---- 865=>x"bb00", 866=>x"bc00", 867=>x"bd00", 868=>x"b300",
---- 869=>x"ba00", 870=>x"bb00", 871=>x"bc00", 872=>x"b500",
---- 873=>x"ba00", 874=>x"bc00", 875=>x"bc00", 876=>x"b500",
---- 877=>x"b600", 878=>x"ba00", 879=>x"be00", 880=>x"b000",
---- 881=>x"4a00", 882=>x"ba00", 883=>x"bf00", 884=>x"b000",
---- 885=>x"b700", 886=>x"ba00", 887=>x"bd00", 888=>x"b200",
---- 889=>x"b600", 890=>x"b900", 891=>x"bc00", 892=>x"b000",
---- 893=>x"b200", 894=>x"b600", 895=>x"b800", 896=>x"5000",
---- 897=>x"af00", 898=>x"b400", 899=>x"b800", 900=>x"ab00",
---- 901=>x"ae00", 902=>x"b500", 903=>x"b800", 904=>x"a900",
---- 905=>x"af00", 906=>x"b400", 907=>x"b700", 908=>x"aa00",
---- 909=>x"aa00", 910=>x"af00", 911=>x"b300", 912=>x"aa00",
---- 913=>x"ae00", 914=>x"ad00", 915=>x"b300", 916=>x"a700",
---- 917=>x"ae00", 918=>x"af00", 919=>x"b300", 920=>x"a800",
---- 921=>x"ab00", 922=>x"ab00", 923=>x"b000", 924=>x"a600",
---- 925=>x"a900", 926=>x"a900", 927=>x"ab00", 928=>x"a600",
---- 929=>x"aa00", 930=>x"a800", 931=>x"ac00", 932=>x"a700",
---- 933=>x"a900", 934=>x"aa00", 935=>x"ab00", 936=>x"a500",
---- 937=>x"a800", 938=>x"a900", 939=>x"a900", 940=>x"a200",
---- 941=>x"a400", 942=>x"a700", 943=>x"a800", 944=>x"a000",
---- 945=>x"a300", 946=>x"a600", 947=>x"a700", 948=>x"9e00",
---- 949=>x"a100", 950=>x"a500", 951=>x"a600", 952=>x"9c00",
---- 953=>x"9f00", 954=>x"a400", 955=>x"a600", 956=>x"9b00",
---- 957=>x"a100", 958=>x"9f00", 959=>x"a700", 960=>x"6200",
---- 961=>x"a100", 962=>x"a000", 963=>x"a400", 964=>x"9c00",
---- 965=>x"9f00", 966=>x"a200", 967=>x"a600", 968=>x"9900",
---- 969=>x"9e00", 970=>x"a200", 971=>x"a200", 972=>x"9a00",
---- 973=>x"9e00", 974=>x"a100", 975=>x"a100", 976=>x"9a00",
---- 977=>x"9b00", 978=>x"6100", 979=>x"9f00", 980=>x"9800",
---- 981=>x"9b00", 982=>x"9d00", 983=>x"9f00", 984=>x"9900",
---- 985=>x"9d00", 986=>x"9f00", 987=>x"9f00", 988=>x"9700",
---- 989=>x"9a00", 990=>x"9f00", 991=>x"9e00", 992=>x"9400",
---- 993=>x"9a00", 994=>x"9b00", 995=>x"9b00", 996=>x"9600",
---- 997=>x"9900", 998=>x"9b00", 999=>x"9a00", 1000=>x"9600",
---- 1001=>x"9500", 1002=>x"9900", 1003=>x"9b00", 1004=>x"9700",
---- 1005=>x"9700", 1006=>x"9700", 1007=>x"9c00", 1008=>x"9900",
---- 1009=>x"9800", 1010=>x"9700", 1011=>x"9d00", 1012=>x"9900",
---- 1013=>x"9b00", 1014=>x"9900", 1015=>x"9c00", 1016=>x"9a00",
---- 1017=>x"9a00", 1018=>x"9a00", 1019=>x"9d00", 1020=>x"9d00",
---- 1021=>x"6100", 1022=>x"9d00", 1023=>x"9e00"),
----
---- 41 => (0=>x"8e00", 1=>x"9200", 2=>x"9800", 3=>x"9a00", 4=>x"8d00",
---- 5=>x"9200", 6=>x"9800", 7=>x"9a00", 8=>x"8c00",
---- 9=>x"9300", 10=>x"9700", 11=>x"9900", 12=>x"8900",
---- 13=>x"9100", 14=>x"9400", 15=>x"9900", 16=>x"8500",
---- 17=>x"8c00", 18=>x"9300", 19=>x"9800", 20=>x"7f00",
---- 21=>x"8800", 22=>x"8e00", 23=>x"9600", 24=>x"7c00",
---- 25=>x"8700", 26=>x"8d00", 27=>x"9300", 28=>x"7400",
---- 29=>x"8100", 30=>x"8d00", 31=>x"9200", 32=>x"6f00",
---- 33=>x"7b00", 34=>x"8a00", 35=>x"9200", 36=>x"6d00",
---- 37=>x"7900", 38=>x"8400", 39=>x"8c00", 40=>x"6c00",
---- 41=>x"7300", 42=>x"7f00", 43=>x"8a00", 44=>x"6a00",
---- 45=>x"6d00", 46=>x"8400", 47=>x"8800", 48=>x"6f00",
---- 49=>x"7200", 50=>x"7c00", 51=>x"8500", 52=>x"6e00",
---- 53=>x"7500", 54=>x"7900", 55=>x"8500", 56=>x"6e00",
---- 57=>x"7500", 58=>x"7d00", 59=>x"8400", 60=>x"6d00",
---- 61=>x"7600", 62=>x"7e00", 63=>x"8600", 64=>x"6c00",
---- 65=>x"7400", 66=>x"8000", 67=>x"8400", 68=>x"7100",
---- 69=>x"7500", 70=>x"7900", 71=>x"8100", 72=>x"6e00",
---- 73=>x"7500", 74=>x"7900", 75=>x"8100", 76=>x"6b00",
---- 77=>x"7000", 78=>x"7a00", 79=>x"8200", 80=>x"6f00",
---- 81=>x"7500", 82=>x"7c00", 83=>x"8100", 84=>x"6d00",
---- 85=>x"7300", 86=>x"7900", 87=>x"7c00", 88=>x"6e00",
---- 89=>x"7000", 90=>x"7300", 91=>x"7d00", 92=>x"6d00",
---- 93=>x"7300", 94=>x"7500", 95=>x"7e00", 96=>x"6c00",
---- 97=>x"6f00", 98=>x"7700", 99=>x"7c00", 100=>x"6c00",
---- 101=>x"6f00", 102=>x"7600", 103=>x"7c00", 104=>x"6a00",
---- 105=>x"6e00", 106=>x"7300", 107=>x"7e00", 108=>x"6c00",
---- 109=>x"7000", 110=>x"7700", 111=>x"8000", 112=>x"6f00",
---- 113=>x"7200", 114=>x"7700", 115=>x"7f00", 116=>x"6c00",
---- 117=>x"7000", 118=>x"7500", 119=>x"7d00", 120=>x"6c00",
---- 121=>x"6f00", 122=>x"7400", 123=>x"7c00", 124=>x"6b00",
---- 125=>x"6f00", 126=>x"7400", 127=>x"8000", 128=>x"6800",
---- 129=>x"6d00", 130=>x"7200", 131=>x"7e00", 132=>x"6500",
---- 133=>x"6e00", 134=>x"7400", 135=>x"8000", 136=>x"6800",
---- 137=>x"6d00", 138=>x"7400", 139=>x"7e00", 140=>x"6600",
---- 141=>x"6d00", 142=>x"7200", 143=>x"7d00", 144=>x"6500",
---- 145=>x"6a00", 146=>x"7300", 147=>x"7e00", 148=>x"6400",
---- 149=>x"9500", 150=>x"7100", 151=>x"7c00", 152=>x"6400",
---- 153=>x"6f00", 154=>x"7200", 155=>x"7f00", 156=>x"6600",
---- 157=>x"6a00", 158=>x"7000", 159=>x"7f00", 160=>x"6500",
---- 161=>x"6c00", 162=>x"7000", 163=>x"7e00", 164=>x"6000",
---- 165=>x"6b00", 166=>x"6f00", 167=>x"7d00", 168=>x"5f00",
---- 169=>x"6b00", 170=>x"7000", 171=>x"7c00", 172=>x"6000",
---- 173=>x"6800", 174=>x"6f00", 175=>x"7b00", 176=>x"6000",
---- 177=>x"9800", 178=>x"7200", 179=>x"7a00", 180=>x"5f00",
---- 181=>x"6500", 182=>x"6e00", 183=>x"7b00", 184=>x"5d00",
---- 185=>x"6600", 186=>x"6f00", 187=>x"7c00", 188=>x"5e00",
---- 189=>x"6500", 190=>x"7000", 191=>x"7d00", 192=>x"5900",
---- 193=>x"6300", 194=>x"7000", 195=>x"7c00", 196=>x"5900",
---- 197=>x"6100", 198=>x"6e00", 199=>x"7d00", 200=>x"5600",
---- 201=>x"6200", 202=>x"6c00", 203=>x"7900", 204=>x"5300",
---- 205=>x"5c00", 206=>x"6c00", 207=>x"7d00", 208=>x"5200",
---- 209=>x"5d00", 210=>x"6b00", 211=>x"7b00", 212=>x"4e00",
---- 213=>x"5900", 214=>x"6800", 215=>x"7900", 216=>x"4700",
---- 217=>x"5600", 218=>x"6400", 219=>x"7500", 220=>x"4700",
---- 221=>x"4f00", 222=>x"6300", 223=>x"7700", 224=>x"3a00",
---- 225=>x"4c00", 226=>x"6000", 227=>x"7600", 228=>x"3100",
---- 229=>x"4d00", 230=>x"5f00", 231=>x"7200", 232=>x"3900",
---- 233=>x"4700", 234=>x"5a00", 235=>x"7200", 236=>x"a500",
---- 237=>x"3d00", 238=>x"5700", 239=>x"6b00", 240=>x"9b00",
---- 241=>x"4000", 242=>x"5100", 243=>x"6a00", 244=>x"d100",
---- 245=>x"7100", 246=>x"4600", 247=>x"6600", 248=>x"e000",
---- 249=>x"b400", 250=>x"5400", 251=>x"5d00", 252=>x"da00",
---- 253=>x"db00", 254=>x"8800", 255=>x"5400", 256=>x"d500",
---- 257=>x"db00", 258=>x"c000", 259=>x"7800", 260=>x"d200",
---- 261=>x"d700", 262=>x"d900", 263=>x"c400", 264=>x"ce00",
---- 265=>x"d400", 266=>x"d500", 267=>x"d800", 268=>x"cb00",
---- 269=>x"cd00", 270=>x"d200", 271=>x"d400", 272=>x"c600",
---- 273=>x"c800", 274=>x"cb00", 275=>x"cf00", 276=>x"c100",
---- 277=>x"c400", 278=>x"c600", 279=>x"c500", 280=>x"c000",
---- 281=>x"bc00", 282=>x"c300", 283=>x"bf00", 284=>x"c000",
---- 285=>x"b800", 286=>x"bc00", 287=>x"bc00", 288=>x"bb00",
---- 289=>x"b800", 290=>x"b800", 291=>x"bf00", 292=>x"bb00",
---- 293=>x"b600", 294=>x"b200", 295=>x"ba00", 296=>x"b900",
---- 297=>x"b300", 298=>x"ac00", 299=>x"aa00", 300=>x"b000",
---- 301=>x"ae00", 302=>x"a200", 303=>x"a200", 304=>x"a200",
---- 305=>x"9f00", 306=>x"a000", 307=>x"ba00", 308=>x"9b00",
---- 309=>x"b000", 310=>x"c900", 311=>x"cc00", 312=>x"c200",
---- 313=>x"d000", 314=>x"c100", 315=>x"b400", 316=>x"c200",
---- 317=>x"b700", 318=>x"b600", 319=>x"ba00", 320=>x"b100",
---- 321=>x"b300", 322=>x"bc00", 323=>x"c500", 324=>x"bc00",
---- 325=>x"c100", 326=>x"c400", 327=>x"cd00", 328=>x"c400",
---- 329=>x"cc00", 330=>x"cb00", 331=>x"cb00", 332=>x"c700",
---- 333=>x"c700", 334=>x"c400", 335=>x"c200", 336=>x"c000",
---- 337=>x"bd00", 338=>x"b900", 339=>x"b700", 340=>x"bb00",
---- 341=>x"bb00", 342=>x"bb00", 343=>x"bc00", 344=>x"bd00",
---- 345=>x"c000", 346=>x"c100", 347=>x"c000", 348=>x"bf00",
---- 349=>x"c000", 350=>x"c000", 351=>x"c000", 352=>x"c300",
---- 353=>x"c300", 354=>x"be00", 355=>x"bf00", 356=>x"c000",
---- 357=>x"c200", 358=>x"bf00", 359=>x"c000", 360=>x"be00",
---- 361=>x"be00", 362=>x"c100", 363=>x"c300", 364=>x"be00",
---- 365=>x"c000", 366=>x"c100", 367=>x"c400", 368=>x"c200",
---- 369=>x"c000", 370=>x"c200", 371=>x"c200", 372=>x"c000",
---- 373=>x"bf00", 374=>x"c000", 375=>x"c000", 376=>x"bd00",
---- 377=>x"c100", 378=>x"c100", 379=>x"c200", 380=>x"bf00",
---- 381=>x"c100", 382=>x"c000", 383=>x"c100", 384=>x"bf00",
---- 385=>x"be00", 386=>x"c200", 387=>x"c200", 388=>x"bf00",
---- 389=>x"c000", 390=>x"c200", 391=>x"c300", 392=>x"bd00",
---- 393=>x"c200", 394=>x"c300", 395=>x"c300", 396=>x"c200",
---- 397=>x"c200", 398=>x"c400", 399=>x"c800", 400=>x"c100",
---- 401=>x"c300", 402=>x"4100", 403=>x"a100", 404=>x"bc00",
---- 405=>x"b900", 406=>x"ac00", 407=>x"7600", 408=>x"b900",
---- 409=>x"c000", 410=>x"b800", 411=>x"a200", 412=>x"c000",
---- 413=>x"c200", 414=>x"bf00", 415=>x"ae00", 416=>x"c600",
---- 417=>x"c400", 418=>x"bf00", 419=>x"b400", 420=>x"c400",
---- 421=>x"ca00", 422=>x"c500", 423=>x"c000", 424=>x"c300",
---- 425=>x"c600", 426=>x"c600", 427=>x"c400", 428=>x"c500",
---- 429=>x"c500", 430=>x"c800", 431=>x"c500", 432=>x"c600",
---- 433=>x"c600", 434=>x"c500", 435=>x"c500", 436=>x"ca00",
---- 437=>x"c800", 438=>x"c900", 439=>x"c400", 440=>x"cb00",
---- 441=>x"cc00", 442=>x"cc00", 443=>x"ca00", 444=>x"d100",
---- 445=>x"d200", 446=>x"cf00", 447=>x"d100", 448=>x"d100",
---- 449=>x"d300", 450=>x"d100", 451=>x"d200", 452=>x"cf00",
---- 453=>x"d200", 454=>x"d100", 455=>x"d300", 456=>x"2c00",
---- 457=>x"d200", 458=>x"d400", 459=>x"d400", 460=>x"d200",
---- 461=>x"d200", 462=>x"d300", 463=>x"d400", 464=>x"d100",
---- 465=>x"d300", 466=>x"d500", 467=>x"d500", 468=>x"d100",
---- 469=>x"d200", 470=>x"d500", 471=>x"d600", 472=>x"d200",
---- 473=>x"d100", 474=>x"d400", 475=>x"d500", 476=>x"cf00",
---- 477=>x"d100", 478=>x"d200", 479=>x"d300", 480=>x"cd00",
---- 481=>x"d100", 482=>x"d200", 483=>x"d300", 484=>x"ca00",
---- 485=>x"ce00", 486=>x"d100", 487=>x"d400", 488=>x"c900",
---- 489=>x"cb00", 490=>x"ce00", 491=>x"d200", 492=>x"c800",
---- 493=>x"ca00", 494=>x"ce00", 495=>x"ce00", 496=>x"c900",
---- 497=>x"c800", 498=>x"cd00", 499=>x"ca00", 500=>x"c200",
---- 501=>x"b900", 502=>x"a900", 503=>x"8d00", 504=>x"aa00",
---- 505=>x"8700", 506=>x"6200", 507=>x"5200", 508=>x"8400",
---- 509=>x"9200", 510=>x"6800", 511=>x"7000", 512=>x"8400",
---- 513=>x"8000", 514=>x"6f00", 515=>x"5500", 516=>x"5900",
---- 517=>x"4600", 518=>x"3600", 519=>x"3100", 520=>x"3300",
---- 521=>x"3200", 522=>x"3200", 523=>x"3900", 524=>x"3500",
---- 525=>x"3a00", 526=>x"3e00", 527=>x"5600", 528=>x"2e00",
---- 529=>x"3e00", 530=>x"7d00", 531=>x"6e00", 532=>x"2b00",
---- 533=>x"4100", 534=>x"6100", 535=>x"6100", 536=>x"4600",
---- 537=>x"5f00", 538=>x"3f00", 539=>x"6000", 540=>x"5f00",
---- 541=>x"4d00", 542=>x"4f00", 543=>x"9a00", 544=>x"5900",
---- 545=>x"6500", 546=>x"9a00", 547=>x"ba00", 548=>x"7100",
---- 549=>x"a100", 550=>x"b000", 551=>x"5300", 552=>x"8600",
---- 553=>x"9000", 554=>x"9400", 555=>x"8100", 556=>x"6d00",
---- 557=>x"8f00", 558=>x"6f00", 559=>x"5b00", 560=>x"7e00",
---- 561=>x"7d00", 562=>x"7d00", 563=>x"7500", 564=>x"8a00",
---- 565=>x"8400", 566=>x"7e00", 567=>x"7c00", 568=>x"9200",
---- 569=>x"8500", 570=>x"8000", 571=>x"8000", 572=>x"9800",
---- 573=>x"8c00", 574=>x"7900", 575=>x"8300", 576=>x"9500",
---- 577=>x"8e00", 578=>x"8900", 579=>x"8600", 580=>x"9200",
---- 581=>x"8d00", 582=>x"8800", 583=>x"8800", 584=>x"9700",
---- 585=>x"8d00", 586=>x"8900", 587=>x"8500", 588=>x"9700",
---- 589=>x"8f00", 590=>x"8800", 591=>x"8600", 592=>x"9b00",
---- 593=>x"9100", 594=>x"8d00", 595=>x"8700", 596=>x"9800",
---- 597=>x"9400", 598=>x"8f00", 599=>x"8900", 600=>x"9900",
---- 601=>x"9200", 602=>x"9000", 603=>x"8a00", 604=>x"9500",
---- 605=>x"9500", 606=>x"9200", 607=>x"8a00", 608=>x"9400",
---- 609=>x"9600", 610=>x"8f00", 611=>x"8b00", 612=>x"9400",
---- 613=>x"9300", 614=>x"8c00", 615=>x"8800", 616=>x"9500",
---- 617=>x"9100", 618=>x"8e00", 619=>x"8a00", 620=>x"9400",
---- 621=>x"9000", 622=>x"8e00", 623=>x"8900", 624=>x"9600",
---- 625=>x"9400", 626=>x"7400", 627=>x"8900", 628=>x"9800",
---- 629=>x"9300", 630=>x"8a00", 631=>x"8700", 632=>x"9600",
---- 633=>x"9000", 634=>x"8b00", 635=>x"8400", 636=>x"9100",
---- 637=>x"8b00", 638=>x"8800", 639=>x"8200", 640=>x"9100",
---- 641=>x"8e00", 642=>x"8a00", 643=>x"8300", 644=>x"9000",
---- 645=>x"8d00", 646=>x"8600", 647=>x"7f00", 648=>x"8d00",
---- 649=>x"8c00", 650=>x"8700", 651=>x"8100", 652=>x"8c00",
---- 653=>x"8a00", 654=>x"8300", 655=>x"8400", 656=>x"8a00",
---- 657=>x"8500", 658=>x"8400", 659=>x"8100", 660=>x"8b00",
---- 661=>x"8500", 662=>x"8200", 663=>x"7800", 664=>x"7800",
---- 665=>x"8300", 666=>x"8300", 667=>x"6b00", 668=>x"8600",
---- 669=>x"8600", 670=>x"7f00", 671=>x"4b00", 672=>x"8700",
---- 673=>x"8a00", 674=>x"6c00", 675=>x"3100", 676=>x"8800",
---- 677=>x"8400", 678=>x"4d00", 679=>x"2a00", 680=>x"8a00",
---- 681=>x"7300", 682=>x"3600", 683=>x"2e00", 684=>x"8800",
---- 685=>x"5500", 686=>x"2900", 687=>x"2e00", 688=>x"7a00",
---- 689=>x"3a00", 690=>x"2a00", 691=>x"2d00", 692=>x"5700",
---- 693=>x"2b00", 694=>x"2f00", 695=>x"2f00", 696=>x"3900",
---- 697=>x"2e00", 698=>x"2e00", 699=>x"2f00", 700=>x"2a00",
---- 701=>x"2f00", 702=>x"2b00", 703=>x"cf00", 704=>x"2a00",
---- 705=>x"2d00", 706=>x"2e00", 707=>x"3300", 708=>x"2f00",
---- 709=>x"2f00", 710=>x"2f00", 711=>x"3700", 712=>x"2a00",
---- 713=>x"2e00", 714=>x"3300", 715=>x"3500", 716=>x"2b00",
---- 717=>x"2d00", 718=>x"3500", 719=>x"3200", 720=>x"2d00",
---- 721=>x"2f00", 722=>x"3800", 723=>x"3000", 724=>x"2f00",
---- 725=>x"3300", 726=>x"3700", 727=>x"3000", 728=>x"2a00",
---- 729=>x"2f00", 730=>x"2d00", 731=>x"3000", 732=>x"2b00",
---- 733=>x"2f00", 734=>x"3500", 735=>x"3500", 736=>x"2d00",
---- 737=>x"3400", 738=>x"3a00", 739=>x"3400", 740=>x"3100",
---- 741=>x"3200", 742=>x"3300", 743=>x"3c00", 744=>x"2f00",
---- 745=>x"3300", 746=>x"3a00", 747=>x"3f00", 748=>x"3200",
---- 749=>x"3900", 750=>x"3f00", 751=>x"3900", 752=>x"3200",
---- 753=>x"3800", 754=>x"4000", 755=>x"3800", 756=>x"3500",
---- 757=>x"3600", 758=>x"c200", 759=>x"4200", 760=>x"3500",
---- 761=>x"3700", 762=>x"3c00", 763=>x"4600", 764=>x"3800",
---- 765=>x"3700", 766=>x"3c00", 767=>x"4a00", 768=>x"3900",
---- 769=>x"3600", 770=>x"4000", 771=>x"4300", 772=>x"3900",
---- 773=>x"3400", 774=>x"4000", 775=>x"4300", 776=>x"3a00",
---- 777=>x"3400", 778=>x"3d00", 779=>x"4200", 780=>x"3500",
---- 781=>x"3300", 782=>x"3600", 783=>x"3a00", 784=>x"3500",
---- 785=>x"3300", 786=>x"3500", 787=>x"3700", 788=>x"3700",
---- 789=>x"3400", 790=>x"3600", 791=>x"3a00", 792=>x"7d00",
---- 793=>x"4600", 794=>x"2f00", 795=>x"2c00", 796=>x"cf00",
---- 797=>x"b000", 798=>x"7800", 799=>x"3e00", 800=>x"cf00",
---- 801=>x"d500", 802=>x"d000", 803=>x"a600", 804=>x"cc00",
---- 805=>x"ce00", 806=>x"d300", 807=>x"d800", 808=>x"cc00",
---- 809=>x"ce00", 810=>x"cf00", 811=>x"d100", 812=>x"cc00",
---- 813=>x"cd00", 814=>x"d000", 815=>x"d000", 816=>x"cb00",
---- 817=>x"cd00", 818=>x"cf00", 819=>x"d100", 820=>x"ca00",
---- 821=>x"3200", 822=>x"cf00", 823=>x"cf00", 824=>x"c900",
---- 825=>x"ca00", 826=>x"ce00", 827=>x"d000", 828=>x"c900",
---- 829=>x"ca00", 830=>x"cb00", 831=>x"cf00", 832=>x"c800",
---- 833=>x"c900", 834=>x"cd00", 835=>x"cf00", 836=>x"c400",
---- 837=>x"c400", 838=>x"cc00", 839=>x"3200", 840=>x"c500",
---- 841=>x"c700", 842=>x"ca00", 843=>x"cb00", 844=>x"c400",
---- 845=>x"c600", 846=>x"ca00", 847=>x"cc00", 848=>x"c500",
---- 849=>x"c500", 850=>x"c900", 851=>x"cc00", 852=>x"c400",
---- 853=>x"c600", 854=>x"c800", 855=>x"cc00", 856=>x"c200",
---- 857=>x"c600", 858=>x"ca00", 859=>x"cc00", 860=>x"c100",
---- 861=>x"c400", 862=>x"c800", 863=>x"cc00", 864=>x"c300",
---- 865=>x"c400", 866=>x"c700", 867=>x"ca00", 868=>x"c200",
---- 869=>x"c300", 870=>x"c600", 871=>x"cc00", 872=>x"bf00",
---- 873=>x"c200", 874=>x"c400", 875=>x"ca00", 876=>x"c100",
---- 877=>x"c300", 878=>x"c500", 879=>x"c800", 880=>x"c000",
---- 881=>x"c100", 882=>x"c600", 883=>x"c700", 884=>x"c000",
---- 885=>x"c000", 886=>x"c500", 887=>x"c800", 888=>x"bd00",
---- 889=>x"3f00", 890=>x"c400", 891=>x"c700", 892=>x"bd00",
---- 893=>x"c000", 894=>x"c300", 895=>x"c500", 896=>x"bf00",
---- 897=>x"c000", 898=>x"c000", 899=>x"c500", 900=>x"ba00",
---- 901=>x"bf00", 902=>x"c100", 903=>x"c500", 904=>x"b900",
---- 905=>x"be00", 906=>x"c300", 907=>x"c200", 908=>x"ba00",
---- 909=>x"ba00", 910=>x"c000", 911=>x"c100", 912=>x"b700",
---- 913=>x"b900", 914=>x"bf00", 915=>x"c000", 916=>x"b500",
---- 917=>x"b700", 918=>x"bb00", 919=>x"c000", 920=>x"b300",
---- 921=>x"b800", 922=>x"bc00", 923=>x"be00", 924=>x"b100",
---- 925=>x"b700", 926=>x"bb00", 927=>x"bd00", 928=>x"ac00",
---- 929=>x"b200", 930=>x"b900", 931=>x"bd00", 932=>x"ad00",
---- 933=>x"b100", 934=>x"ba00", 935=>x"b900", 936=>x"a900",
---- 937=>x"b100", 938=>x"b600", 939=>x"b800", 940=>x"ad00",
---- 941=>x"b100", 942=>x"b300", 943=>x"b900", 944=>x"ac00",
---- 945=>x"b200", 946=>x"b000", 947=>x"b600", 948=>x"ac00",
---- 949=>x"b300", 950=>x"af00", 951=>x"b500", 952=>x"ab00",
---- 953=>x"ae00", 954=>x"ae00", 955=>x"b400", 956=>x"ab00",
---- 957=>x"a800", 958=>x"ab00", 959=>x"b200", 960=>x"a400",
---- 961=>x"a700", 962=>x"ab00", 963=>x"ad00", 964=>x"a200",
---- 965=>x"a400", 966=>x"ac00", 967=>x"b100", 968=>x"a300",
---- 969=>x"a600", 970=>x"a900", 971=>x"aa00", 972=>x"a200",
---- 973=>x"a800", 974=>x"a800", 975=>x"a700", 976=>x"a100",
---- 977=>x"a800", 978=>x"a800", 979=>x"aa00", 980=>x"a100",
---- 981=>x"a400", 982=>x"a800", 983=>x"aa00", 984=>x"a000",
---- 985=>x"a300", 986=>x"a600", 987=>x"a900", 988=>x"9d00",
---- 989=>x"a400", 990=>x"a500", 991=>x"a600", 992=>x"9d00",
---- 993=>x"a200", 994=>x"a400", 995=>x"aa00", 996=>x"9d00",
---- 997=>x"a000", 998=>x"a400", 999=>x"a600", 1000=>x"9d00",
---- 1001=>x"a200", 1002=>x"a300", 1003=>x"a600", 1004=>x"9e00",
---- 1005=>x"a000", 1006=>x"a500", 1007=>x"a500", 1008=>x"a000",
---- 1009=>x"a200", 1010=>x"a600", 1011=>x"a700", 1012=>x"a000",
---- 1013=>x"a000", 1014=>x"a400", 1015=>x"a300", 1016=>x"9c00",
---- 1017=>x"5e00", 1018=>x"a500", 1019=>x"a400", 1020=>x"9e00",
---- 1021=>x"a100", 1022=>x"a300", 1023=>x"a800"),
----
---- 42 => (0=>x"9f00", 1=>x"a100", 2=>x"a000", 3=>x"9e00", 4=>x"9f00",
---- 5=>x"a000", 6=>x"a100", 7=>x"9d00", 8=>x"9f00",
---- 9=>x"a100", 10=>x"a200", 11=>x"9e00", 12=>x"9d00",
---- 13=>x"a000", 14=>x"a100", 15=>x"9d00", 16=>x"9a00",
---- 17=>x"9d00", 18=>x"a100", 19=>x"a000", 20=>x"9800",
---- 21=>x"9c00", 22=>x"a100", 23=>x"a000", 24=>x"9800",
---- 25=>x"9a00", 26=>x"a100", 27=>x"a000", 28=>x"9700",
---- 29=>x"9900", 30=>x"9d00", 31=>x"a100", 32=>x"9300",
---- 33=>x"9700", 34=>x"9b00", 35=>x"9d00", 36=>x"8f00",
---- 37=>x"9800", 38=>x"6500", 39=>x"9e00", 40=>x"9200",
---- 41=>x"9500", 42=>x"6500", 43=>x"6300", 44=>x"9100",
---- 45=>x"9700", 46=>x"9900", 47=>x"9b00", 48=>x"8d00",
---- 49=>x"9500", 50=>x"9900", 51=>x"9e00", 52=>x"8d00",
---- 53=>x"9100", 54=>x"9900", 55=>x"9e00", 56=>x"8b00",
---- 57=>x"9300", 58=>x"9900", 59=>x"9c00", 60=>x"8a00",
---- 61=>x"9200", 62=>x"9600", 63=>x"9a00", 64=>x"8800",
---- 65=>x"8d00", 66=>x"9300", 67=>x"9900", 68=>x"8900",
---- 69=>x"8d00", 70=>x"9300", 71=>x"9800", 72=>x"8900",
---- 73=>x"8c00", 74=>x"8f00", 75=>x"9500", 76=>x"8700",
---- 77=>x"8b00", 78=>x"8f00", 79=>x"9400", 80=>x"8500",
---- 81=>x"8c00", 82=>x"9000", 83=>x"9300", 84=>x"8600",
---- 85=>x"8a00", 86=>x"8f00", 87=>x"9000", 88=>x"8200",
---- 89=>x"8b00", 90=>x"8c00", 91=>x"9000", 92=>x"8500",
---- 93=>x"8a00", 94=>x"8d00", 95=>x"9100", 96=>x"8200",
---- 97=>x"8a00", 98=>x"8f00", 99=>x"9000", 100=>x"8500",
---- 101=>x"8a00", 102=>x"8c00", 103=>x"9100", 104=>x"8600",
---- 105=>x"8b00", 106=>x"8d00", 107=>x"9500", 108=>x"8500",
---- 109=>x"8a00", 110=>x"8f00", 111=>x"9100", 112=>x"8800",
---- 113=>x"8e00", 114=>x"8f00", 115=>x"9000", 116=>x"8400",
---- 117=>x"8b00", 118=>x"8e00", 119=>x"9200", 120=>x"8500",
---- 121=>x"8c00", 122=>x"8f00", 123=>x"9200", 124=>x"8900",
---- 125=>x"7300", 126=>x"8f00", 127=>x"9200", 128=>x"8600",
---- 129=>x"8c00", 130=>x"9000", 131=>x"9400", 132=>x"8700",
---- 133=>x"8c00", 134=>x"9100", 135=>x"9300", 136=>x"8900",
---- 137=>x"8f00", 138=>x"9300", 139=>x"9600", 140=>x"8700",
---- 141=>x"8e00", 142=>x"9300", 143=>x"9700", 144=>x"8700",
---- 145=>x"8f00", 146=>x"9200", 147=>x"9800", 148=>x"8a00",
---- 149=>x"9600", 150=>x"9500", 151=>x"9900", 152=>x"8b00",
---- 153=>x"9300", 154=>x"9700", 155=>x"9a00", 156=>x"8900",
---- 157=>x"9100", 158=>x"9500", 159=>x"9800", 160=>x"8700",
---- 161=>x"9000", 162=>x"9500", 163=>x"9900", 164=>x"8900",
---- 165=>x"8f00", 166=>x"9400", 167=>x"9600", 168=>x"8500",
---- 169=>x"8e00", 170=>x"9300", 171=>x"9900", 172=>x"8500",
---- 173=>x"8d00", 174=>x"9500", 175=>x"9b00", 176=>x"8500",
---- 177=>x"8d00", 178=>x"9600", 179=>x"9900", 180=>x"8500",
---- 181=>x"8c00", 182=>x"9500", 183=>x"9a00", 184=>x"8600",
---- 185=>x"8d00", 186=>x"9500", 187=>x"9b00", 188=>x"8700",
---- 189=>x"8f00", 190=>x"9500", 191=>x"9900", 192=>x"8600",
---- 193=>x"8d00", 194=>x"9400", 195=>x"9b00", 196=>x"8600",
---- 197=>x"8e00", 198=>x"9300", 199=>x"9a00", 200=>x"8600",
---- 201=>x"8f00", 202=>x"9600", 203=>x"9800", 204=>x"8600",
---- 205=>x"8d00", 206=>x"9500", 207=>x"9b00", 208=>x"8200",
---- 209=>x"8a00", 210=>x"9500", 211=>x"9800", 212=>x"8400",
---- 213=>x"8b00", 214=>x"9400", 215=>x"9700", 216=>x"8000",
---- 217=>x"8c00", 218=>x"9300", 219=>x"9700", 220=>x"8200",
---- 221=>x"8c00", 222=>x"9100", 223=>x"9700", 224=>x"8200",
---- 225=>x"8900", 226=>x"9400", 227=>x"9800", 228=>x"8300",
---- 229=>x"8b00", 230=>x"9300", 231=>x"9700", 232=>x"8100",
---- 233=>x"8b00", 234=>x"9300", 235=>x"9600", 236=>x"7e00",
---- 237=>x"8900", 238=>x"9200", 239=>x"9500", 240=>x"7d00",
---- 241=>x"8800", 242=>x"9700", 243=>x"9600", 244=>x"7b00",
---- 245=>x"8900", 246=>x"8f00", 247=>x"9b00", 248=>x"7b00",
---- 249=>x"8600", 250=>x"8d00", 251=>x"9c00", 252=>x"7900",
---- 253=>x"8600", 254=>x"9000", 255=>x"9800", 256=>x"7100",
---- 257=>x"8200", 258=>x"8f00", 259=>x"9600", 260=>x"9300",
---- 261=>x"7f00", 262=>x"8c00", 263=>x"9600", 264=>x"d500",
---- 265=>x"a200", 266=>x"8500", 267=>x"9400", 268=>x"da00",
---- 269=>x"cf00", 270=>x"9a00", 271=>x"8f00", 272=>x"cf00",
---- 273=>x"d500", 274=>x"ba00", 275=>x"8f00", 276=>x"cd00",
---- 277=>x"d100", 278=>x"cd00", 279=>x"9c00", 280=>x"c200",
---- 281=>x"ca00", 282=>x"d000", 283=>x"a600", 284=>x"b900",
---- 285=>x"c100", 286=>x"ca00", 287=>x"bb00", 288=>x"ba00",
---- 289=>x"bb00", 290=>x"be00", 291=>x"cb00", 292=>x"b900",
---- 293=>x"b800", 294=>x"ba00", 295=>x"c100", 296=>x"b400",
---- 297=>x"b200", 298=>x"ba00", 299=>x"c300", 300=>x"af00",
---- 301=>x"c300", 302=>x"cc00", 303=>x"c300", 304=>x"cb00",
---- 305=>x"c800", 306=>x"b700", 307=>x"aa00", 308=>x"bd00",
---- 309=>x"b200", 310=>x"b700", 311=>x"bb00", 312=>x"b900",
---- 313=>x"c000", 314=>x"c200", 315=>x"c600", 316=>x"c200",
---- 317=>x"c300", 318=>x"c800", 319=>x"ce00", 320=>x"c800",
---- 321=>x"cc00", 322=>x"ce00", 323=>x"cb00", 324=>x"d100",
---- 325=>x"cc00", 326=>x"c900", 327=>x"c500", 328=>x"c800",
---- 329=>x"c500", 330=>x"c300", 331=>x"c100", 332=>x"bb00",
---- 333=>x"b800", 334=>x"be00", 335=>x"c000", 336=>x"b600",
---- 337=>x"b900", 338=>x"bd00", 339=>x"c100", 340=>x"bd00",
---- 341=>x"c000", 342=>x"c300", 343=>x"c400", 344=>x"c000",
---- 345=>x"c100", 346=>x"c300", 347=>x"c600", 348=>x"c300",
---- 349=>x"c000", 350=>x"c500", 351=>x"c800", 352=>x"c300",
---- 353=>x"c400", 354=>x"c600", 355=>x"c900", 356=>x"c400",
---- 357=>x"c400", 358=>x"c700", 359=>x"ca00", 360=>x"c400",
---- 361=>x"c600", 362=>x"c700", 363=>x"c800", 364=>x"c300",
---- 365=>x"c600", 366=>x"c600", 367=>x"c700", 368=>x"c200",
---- 369=>x"c600", 370=>x"c400", 371=>x"c300", 372=>x"c200",
---- 373=>x"c400", 374=>x"c400", 375=>x"c600", 376=>x"c400",
---- 377=>x"c400", 378=>x"c400", 379=>x"c600", 380=>x"c300",
---- 381=>x"c500", 382=>x"c400", 383=>x"c500", 384=>x"c200",
---- 385=>x"c500", 386=>x"c600", 387=>x"c600", 388=>x"c500",
---- 389=>x"c700", 390=>x"cf00", 391=>x"bd00", 392=>x"c800",
---- 393=>x"ca00", 394=>x"6e00", 395=>x"5e00", 396=>x"b700",
---- 397=>x"6200", 398=>x"2c00", 399=>x"5600", 400=>x"5f00",
---- 401=>x"2b00", 402=>x"2c00", 403=>x"5900", 404=>x"4d00",
---- 405=>x"5000", 406=>x"5100", 407=>x"4400", 408=>x"6900",
---- 409=>x"4a00", 410=>x"a500", 411=>x"6400", 412=>x"8400",
---- 413=>x"5d00", 414=>x"4c00", 415=>x"5200", 416=>x"9600",
---- 417=>x"6e00", 418=>x"5d00", 419=>x"5000", 420=>x"ab00",
---- 421=>x"8600", 422=>x"6000", 423=>x"5800", 424=>x"b700",
---- 425=>x"6800", 426=>x"7000", 427=>x"5800", 428=>x"b900",
---- 429=>x"9f00", 430=>x"7700", 431=>x"6100", 432=>x"b700",
---- 433=>x"a500", 434=>x"8500", 435=>x"6300", 436=>x"be00",
---- 437=>x"aa00", 438=>x"8800", 439=>x"6700", 440=>x"c300",
---- 441=>x"b100", 442=>x"9200", 443=>x"6b00", 444=>x"c800",
---- 445=>x"b900", 446=>x"a000", 447=>x"7500", 448=>x"cd00",
---- 449=>x"c100", 450=>x"a800", 451=>x"8000", 452=>x"d000",
---- 453=>x"c300", 454=>x"b200", 455=>x"8e00", 456=>x"cf00",
---- 457=>x"c700", 458=>x"b900", 459=>x"9700", 460=>x"d100",
---- 461=>x"cc00", 462=>x"be00", 463=>x"9f00", 464=>x"d400",
---- 465=>x"d000", 466=>x"c200", 467=>x"a600", 468=>x"d600",
---- 469=>x"d100", 470=>x"c800", 471=>x"ac00", 472=>x"d500",
---- 473=>x"d500", 474=>x"cd00", 475=>x"b300", 476=>x"d500",
---- 477=>x"d100", 478=>x"cc00", 479=>x"be00", 480=>x"d300",
---- 481=>x"d200", 482=>x"cf00", 483=>x"c400", 484=>x"d300",
---- 485=>x"d000", 486=>x"3000", 487=>x"c600", 488=>x"d100",
---- 489=>x"cd00", 490=>x"c900", 491=>x"bd00", 492=>x"ce00",
---- 493=>x"c900", 494=>x"b900", 495=>x"a100", 496=>x"bb00",
---- 497=>x"a300", 498=>x"8900", 499=>x"7600", 500=>x"7300",
---- 501=>x"5e00", 502=>x"4f00", 503=>x"4f00", 504=>x"5c00",
---- 505=>x"5e00", 506=>x"6900", 507=>x"6c00", 508=>x"7b00",
---- 509=>x"9900", 510=>x"6700", 511=>x"6f00", 512=>x"4d00",
---- 513=>x"3800", 514=>x"3900", 515=>x"4100", 516=>x"3000",
---- 517=>x"2f00", 518=>x"3000", 519=>x"3300", 520=>x"3c00",
---- 521=>x"3100", 522=>x"3100", 523=>x"3400", 524=>x"7d00",
---- 525=>x"5800", 526=>x"3400", 527=>x"2a00", 528=>x"a500",
---- 529=>x"8500", 530=>x"4f00", 531=>x"2c00", 532=>x"aa00",
---- 533=>x"9d00", 534=>x"6600", 535=>x"3c00", 536=>x"b000",
---- 537=>x"9d00", 538=>x"7000", 539=>x"4200", 540=>x"b000",
---- 541=>x"9a00", 542=>x"6d00", 543=>x"4300", 544=>x"ae00",
---- 545=>x"9500", 546=>x"6700", 547=>x"4200", 548=>x"9d00",
---- 549=>x"8000", 550=>x"5a00", 551=>x"3600", 552=>x"6700",
---- 553=>x"5700", 554=>x"4000", 555=>x"3000", 556=>x"3d00",
---- 557=>x"4200", 558=>x"4c00", 559=>x"5000", 560=>x"5d00",
---- 561=>x"5b00", 562=>x"5400", 563=>x"6100", 564=>x"6800",
---- 565=>x"6700", 566=>x"6300", 567=>x"6800", 568=>x"7a00",
---- 569=>x"7300", 570=>x"7200", 571=>x"7200", 572=>x"7e00",
---- 573=>x"7700", 574=>x"7400", 575=>x"7200", 576=>x"8000",
---- 577=>x"7d00", 578=>x"7a00", 579=>x"7700", 580=>x"8500",
---- 581=>x"7f00", 582=>x"7c00", 583=>x"7900", 584=>x"8300",
---- 585=>x"8000", 586=>x"8100", 587=>x"7c00", 588=>x"8200",
---- 589=>x"8100", 590=>x"8000", 591=>x"7c00", 592=>x"8500",
---- 593=>x"8100", 594=>x"8000", 595=>x"7e00", 596=>x"8600",
---- 597=>x"8200", 598=>x"8000", 599=>x"7e00", 600=>x"8500",
---- 601=>x"8200", 602=>x"7f00", 603=>x"7d00", 604=>x"8700",
---- 605=>x"8200", 606=>x"8000", 607=>x"7a00", 608=>x"8700",
---- 609=>x"8200", 610=>x"8000", 611=>x"7b00", 612=>x"8500",
---- 613=>x"8200", 614=>x"7f00", 615=>x"7b00", 616=>x"8200",
---- 617=>x"8400", 618=>x"8000", 619=>x"7300", 620=>x"8300",
---- 621=>x"8200", 622=>x"7d00", 623=>x"6e00", 624=>x"8400",
---- 625=>x"8100", 626=>x"7b00", 627=>x"6700", 628=>x"8100",
---- 629=>x"7e00", 630=>x"7a00", 631=>x"6500", 632=>x"8200",
---- 633=>x"7c00", 634=>x"7400", 635=>x"5900", 636=>x"7f00",
---- 637=>x"7b00", 638=>x"6f00", 639=>x"4100", 640=>x"7d00",
---- 641=>x"7a00", 642=>x"5800", 643=>x"3100", 644=>x"7d00",
---- 645=>x"7000", 646=>x"3d00", 647=>x"2800", 648=>x"7f00",
---- 649=>x"5b00", 650=>x"2e00", 651=>x"2d00", 652=>x"7600",
---- 653=>x"bc00", 654=>x"d200", 655=>x"3200", 656=>x"6200",
---- 657=>x"3000", 658=>x"2e00", 659=>x"3400", 660=>x"4600",
---- 661=>x"2d00", 662=>x"2e00", 663=>x"3000", 664=>x"3300",
---- 665=>x"3300", 666=>x"2f00", 667=>x"2d00", 668=>x"2e00",
---- 669=>x"3300", 670=>x"3100", 671=>x"3100", 672=>x"3000",
---- 673=>x"3200", 674=>x"2f00", 675=>x"2f00", 676=>x"3000",
---- 677=>x"3200", 678=>x"3000", 679=>x"3200", 680=>x"2e00",
---- 681=>x"2e00", 682=>x"3000", 683=>x"3200", 684=>x"2d00",
---- 685=>x"3500", 686=>x"ca00", 687=>x"2f00", 688=>x"2e00",
---- 689=>x"3b00", 690=>x"3700", 691=>x"2d00", 692=>x"3200",
---- 693=>x"3500", 694=>x"3100", 695=>x"3100", 696=>x"3500",
---- 697=>x"2f00", 698=>x"3100", 699=>x"3100", 700=>x"3800",
---- 701=>x"3000", 702=>x"2e00", 703=>x"3100", 704=>x"3500",
---- 705=>x"2c00", 706=>x"2b00", 707=>x"3300", 708=>x"3300",
---- 709=>x"2e00", 710=>x"2f00", 711=>x"3400", 712=>x"3000",
---- 713=>x"2a00", 714=>x"2c00", 715=>x"3600", 716=>x"2e00",
---- 717=>x"2900", 718=>x"2c00", 719=>x"3300", 720=>x"3100",
---- 721=>x"2e00", 722=>x"3200", 723=>x"3100", 724=>x"3900",
---- 725=>x"3100", 726=>x"3700", 727=>x"3400", 728=>x"3900",
---- 729=>x"3700", 730=>x"3500", 731=>x"3500", 732=>x"3a00",
---- 733=>x"4400", 734=>x"3500", 735=>x"3600", 736=>x"3900",
---- 737=>x"3f00", 738=>x"3400", 739=>x"3400", 740=>x"3700",
---- 741=>x"3d00", 742=>x"3500", 743=>x"3600", 744=>x"3e00",
---- 745=>x"3f00", 746=>x"3200", 747=>x"3600", 748=>x"3f00",
---- 749=>x"3400", 750=>x"3700", 751=>x"4100", 752=>x"3e00",
---- 753=>x"2d00", 754=>x"3d00", 755=>x"4000", 756=>x"3600",
---- 757=>x"2d00", 758=>x"c700", 759=>x"3700", 760=>x"3200",
---- 761=>x"3200", 762=>x"3500", 763=>x"3400", 764=>x"3600",
---- 765=>x"3a00", 766=>x"3500", 767=>x"3400", 768=>x"3300",
---- 769=>x"3a00", 770=>x"3800", 771=>x"3300", 772=>x"3600",
---- 773=>x"3600", 774=>x"3200", 775=>x"3400", 776=>x"3900",
---- 777=>x"3700", 778=>x"3200", 779=>x"3600", 780=>x"3500",
---- 781=>x"3100", 782=>x"d200", 783=>x"3900", 784=>x"3200",
---- 785=>x"2e00", 786=>x"2c00", 787=>x"3700", 788=>x"3800",
---- 789=>x"3100", 790=>x"3200", 791=>x"3300", 792=>x"3400",
---- 793=>x"2a00", 794=>x"2c00", 795=>x"2800", 796=>x"2a00",
---- 797=>x"2600", 798=>x"2700", 799=>x"2200", 800=>x"5d00",
---- 801=>x"2b00", 802=>x"2500", 803=>x"2400", 804=>x"c400",
---- 805=>x"8200", 806=>x"3700", 807=>x"2300", 808=>x"d500",
---- 809=>x"d300", 810=>x"9c00", 811=>x"4800", 812=>x"d100",
---- 813=>x"d400", 814=>x"2800", 815=>x"ae00", 816=>x"d300",
---- 817=>x"d200", 818=>x"d400", 819=>x"d800", 820=>x"d100",
---- 821=>x"d300", 822=>x"d500", 823=>x"d600", 824=>x"d100",
---- 825=>x"d300", 826=>x"d400", 827=>x"d500", 828=>x"d100",
---- 829=>x"d100", 830=>x"d400", 831=>x"d600", 832=>x"d100",
---- 833=>x"d300", 834=>x"d300", 835=>x"d500", 836=>x"ce00",
---- 837=>x"d100", 838=>x"d200", 839=>x"d400", 840=>x"cc00",
---- 841=>x"d000", 842=>x"d000", 843=>x"d100", 844=>x"cd00",
---- 845=>x"d000", 846=>x"cf00", 847=>x"d200", 848=>x"ce00",
---- 849=>x"d000", 850=>x"d000", 851=>x"d100", 852=>x"ce00",
---- 853=>x"d100", 854=>x"d200", 855=>x"d300", 856=>x"ce00",
---- 857=>x"d100", 858=>x"d000", 859=>x"d400", 860=>x"ce00",
---- 861=>x"d000", 862=>x"cf00", 863=>x"d200", 864=>x"cd00",
---- 865=>x"d000", 866=>x"d100", 867=>x"d300", 868=>x"ce00",
---- 869=>x"ce00", 870=>x"d300", 871=>x"d200", 872=>x"cb00",
---- 873=>x"cf00", 874=>x"cf00", 875=>x"cf00", 876=>x"ca00",
---- 877=>x"cf00", 878=>x"d100", 879=>x"ce00", 880=>x"ca00",
---- 881=>x"d000", 882=>x"ce00", 883=>x"cf00", 884=>x"ca00",
---- 885=>x"cc00", 886=>x"cd00", 887=>x"cf00", 888=>x"c900",
---- 889=>x"cc00", 890=>x"cd00", 891=>x"ce00", 892=>x"c600",
---- 893=>x"ca00", 894=>x"cc00", 895=>x"cd00", 896=>x"c500",
---- 897=>x"c900", 898=>x"cc00", 899=>x"d000", 900=>x"c700",
---- 901=>x"c800", 902=>x"c900", 903=>x"cd00", 904=>x"c600",
---- 905=>x"c800", 906=>x"c900", 907=>x"cb00", 908=>x"c300",
---- 909=>x"c800", 910=>x"c800", 911=>x"cb00", 912=>x"c300",
---- 913=>x"c600", 914=>x"c700", 915=>x"c900", 916=>x"c200",
---- 917=>x"3a00", 918=>x"c600", 919=>x"ca00", 920=>x"c200",
---- 921=>x"c400", 922=>x"c600", 923=>x"ca00", 924=>x"bf00",
---- 925=>x"c200", 926=>x"c300", 927=>x"3700", 928=>x"bf00",
---- 929=>x"c000", 930=>x"c100", 931=>x"c800", 932=>x"be00",
---- 933=>x"bf00", 934=>x"c400", 935=>x"c800", 936=>x"bc00",
---- 937=>x"bf00", 938=>x"c500", 939=>x"c700", 940=>x"bc00",
---- 941=>x"bd00", 942=>x"c200", 943=>x"c800", 944=>x"b800",
---- 945=>x"ba00", 946=>x"bf00", 947=>x"c500", 948=>x"b800",
---- 949=>x"bb00", 950=>x"c000", 951=>x"3c00", 952=>x"b700",
---- 953=>x"ba00", 954=>x"bf00", 955=>x"c200", 956=>x"b300",
---- 957=>x"ba00", 958=>x"4100", 959=>x"c100", 960=>x"b300",
---- 961=>x"b900", 962=>x"bb00", 963=>x"c000", 964=>x"b100",
---- 965=>x"b500", 966=>x"b700", 967=>x"bd00", 968=>x"ad00",
---- 969=>x"b000", 970=>x"b600", 971=>x"ba00", 972=>x"ac00",
---- 973=>x"b100", 974=>x"b300", 975=>x"b800", 976=>x"ad00",
---- 977=>x"af00", 978=>x"b200", 979=>x"b700", 980=>x"af00",
---- 981=>x"af00", 982=>x"b100", 983=>x"b400", 984=>x"b000",
---- 985=>x"b100", 986=>x"b200", 987=>x"b500", 988=>x"a900",
---- 989=>x"b000", 990=>x"b300", 991=>x"b700", 992=>x"a900",
---- 993=>x"af00", 994=>x"ae00", 995=>x"b300", 996=>x"a700",
---- 997=>x"aa00", 998=>x"ab00", 999=>x"b100", 1000=>x"a800",
---- 1001=>x"a900", 1002=>x"ad00", 1003=>x"b200", 1004=>x"aa00",
---- 1005=>x"a900", 1006=>x"ac00", 1007=>x"b000", 1008=>x"a800",
---- 1009=>x"a500", 1010=>x"ad00", 1011=>x"b200", 1012=>x"a200",
---- 1013=>x"a600", 1014=>x"aa00", 1015=>x"af00", 1016=>x"a400",
---- 1017=>x"a400", 1018=>x"a900", 1019=>x"ab00", 1020=>x"a500",
---- 1021=>x"a400", 1022=>x"a900", 1023=>x"a800"),
----
---- 43 => (0=>x"9600", 1=>x"9700", 2=>x"9800", 3=>x"9800", 4=>x"9600",
---- 5=>x"9700", 6=>x"9700", 7=>x"9800", 8=>x"9600",
---- 9=>x"9800", 10=>x"9800", 11=>x"9800", 12=>x"9a00",
---- 13=>x"9800", 14=>x"9800", 15=>x"9900", 16=>x"9c00",
---- 17=>x"9900", 18=>x"9900", 19=>x"9800", 20=>x"9c00",
---- 21=>x"9b00", 22=>x"9a00", 23=>x"9b00", 24=>x"9f00",
---- 25=>x"9d00", 26=>x"9a00", 27=>x"9d00", 28=>x"a200",
---- 29=>x"a100", 30=>x"a000", 31=>x"9f00", 32=>x"a000",
---- 33=>x"a300", 34=>x"a200", 35=>x"a100", 36=>x"a100",
---- 37=>x"a400", 38=>x"a100", 39=>x"a200", 40=>x"a000",
---- 41=>x"a400", 42=>x"a300", 43=>x"a300", 44=>x"a000",
---- 45=>x"a100", 46=>x"a300", 47=>x"a400", 48=>x"9f00",
---- 49=>x"5c00", 50=>x"a300", 51=>x"a200", 52=>x"a100",
---- 53=>x"a100", 54=>x"a200", 55=>x"a200", 56=>x"9f00",
---- 57=>x"a000", 58=>x"a200", 59=>x"a100", 60=>x"9e00",
---- 61=>x"9c00", 62=>x"9e00", 63=>x"a300", 64=>x"9c00",
---- 65=>x"9d00", 66=>x"9e00", 67=>x"a000", 68=>x"9900",
---- 69=>x"9b00", 70=>x"9e00", 71=>x"9f00", 72=>x"9800",
---- 73=>x"9a00", 74=>x"9c00", 75=>x"9c00", 76=>x"9600",
---- 77=>x"9800", 78=>x"9b00", 79=>x"9900", 80=>x"9400",
---- 81=>x"9600", 82=>x"9a00", 83=>x"9b00", 84=>x"9300",
---- 85=>x"9500", 86=>x"9700", 87=>x"9900", 88=>x"9200",
---- 89=>x"9300", 90=>x"9400", 91=>x"9700", 92=>x"9100",
---- 93=>x"9200", 94=>x"9200", 95=>x"9600", 96=>x"9000",
---- 97=>x"8e00", 98=>x"9100", 99=>x"9200", 100=>x"9100",
---- 101=>x"7000", 102=>x"9000", 103=>x"9100", 104=>x"9000",
---- 105=>x"9000", 106=>x"8f00", 107=>x"9200", 108=>x"9200",
---- 109=>x"8f00", 110=>x"9100", 111=>x"9000", 112=>x"9200",
---- 113=>x"9100", 114=>x"8f00", 115=>x"9000", 116=>x"9200",
---- 117=>x"9200", 118=>x"9000", 119=>x"9200", 120=>x"9200",
---- 121=>x"9200", 122=>x"9000", 123=>x"9100", 124=>x"9500",
---- 125=>x"9200", 126=>x"9100", 127=>x"9100", 128=>x"9700",
---- 129=>x"9300", 130=>x"9200", 131=>x"9100", 132=>x"9700",
---- 133=>x"9700", 134=>x"9500", 135=>x"9200", 136=>x"9900",
---- 137=>x"9600", 138=>x"9600", 139=>x"9400", 140=>x"9900",
---- 141=>x"9800", 142=>x"9600", 143=>x"9700", 144=>x"9900",
---- 145=>x"9900", 146=>x"9900", 147=>x"9600", 148=>x"9700",
---- 149=>x"9c00", 150=>x"9d00", 151=>x"9b00", 152=>x"9b00",
---- 153=>x"9b00", 154=>x"9f00", 155=>x"9c00", 156=>x"9e00",
---- 157=>x"9b00", 158=>x"9d00", 159=>x"9b00", 160=>x"9b00",
---- 161=>x"9a00", 162=>x"9c00", 163=>x"9a00", 164=>x"9b00",
---- 165=>x"9900", 166=>x"9b00", 167=>x"9a00", 168=>x"9d00",
---- 169=>x"9900", 170=>x"9800", 171=>x"9900", 172=>x"9d00",
---- 173=>x"9900", 174=>x"9800", 175=>x"9900", 176=>x"9a00",
---- 177=>x"9a00", 178=>x"9900", 179=>x"9900", 180=>x"9c00",
---- 181=>x"9c00", 182=>x"9d00", 183=>x"9a00", 184=>x"9d00",
---- 185=>x"9b00", 186=>x"9a00", 187=>x"9b00", 188=>x"9d00",
---- 189=>x"9a00", 190=>x"9b00", 191=>x"9800", 192=>x"9b00",
---- 193=>x"9a00", 194=>x"9c00", 195=>x"9800", 196=>x"9b00",
---- 197=>x"9a00", 198=>x"9b00", 199=>x"9c00", 200=>x"9c00",
---- 201=>x"9a00", 202=>x"9a00", 203=>x"9900", 204=>x"9c00",
---- 205=>x"9a00", 206=>x"9b00", 207=>x"9900", 208=>x"9a00",
---- 209=>x"9900", 210=>x"9900", 211=>x"9a00", 212=>x"9a00",
---- 213=>x"9a00", 214=>x"9900", 215=>x"9b00", 216=>x"9a00",
---- 217=>x"9a00", 218=>x"9b00", 219=>x"9a00", 220=>x"9900",
---- 221=>x"9800", 222=>x"9b00", 223=>x"9c00", 224=>x"9700",
---- 225=>x"9800", 226=>x"9900", 227=>x"9800", 228=>x"6900",
---- 229=>x"9700", 230=>x"9900", 231=>x"9900", 232=>x"9800",
---- 233=>x"9a00", 234=>x"9a00", 235=>x"9900", 236=>x"9700",
---- 237=>x"9900", 238=>x"9c00", 239=>x"9a00", 240=>x"9900",
---- 241=>x"9800", 242=>x"9900", 243=>x"9b00", 244=>x"9c00",
---- 245=>x"9a00", 246=>x"9d00", 247=>x"9c00", 248=>x"a000",
---- 249=>x"9a00", 250=>x"9e00", 251=>x"9d00", 252=>x"9b00",
---- 253=>x"9900", 254=>x"9d00", 255=>x"9d00", 256=>x"9900",
---- 257=>x"9b00", 258=>x"9c00", 259=>x"9c00", 260=>x"9800",
---- 261=>x"9900", 262=>x"9b00", 263=>x"9c00", 264=>x"9600",
---- 265=>x"9700", 266=>x"9900", 267=>x"9900", 268=>x"9a00",
---- 269=>x"9a00", 270=>x"9800", 271=>x"9700", 272=>x"9a00",
---- 273=>x"9a00", 274=>x"9700", 275=>x"9500", 276=>x"9600",
---- 277=>x"9a00", 278=>x"9600", 279=>x"9400", 280=>x"9200",
---- 281=>x"9900", 282=>x"9700", 283=>x"9100", 284=>x"9200",
---- 285=>x"9200", 286=>x"9600", 287=>x"a900", 288=>x"a800",
---- 289=>x"9800", 290=>x"b800", 291=>x"d300", 292=>x"c000",
---- 293=>x"c500", 294=>x"d300", 295=>x"cb00", 296=>x"cb00",
---- 297=>x"c500", 298=>x"be00", 299=>x"c000", 300=>x"b900",
---- 301=>x"ad00", 302=>x"b700", 303=>x"c700", 304=>x"b900",
---- 305=>x"c100", 306=>x"c700", 307=>x"c800", 308=>x"c200",
---- 309=>x"c800", 310=>x"ca00", 311=>x"d000", 312=>x"ca00",
---- 313=>x"ca00", 314=>x"cd00", 315=>x"cb00", 316=>x"cd00",
---- 317=>x"c700", 318=>x"c700", 319=>x"c700", 320=>x"c900",
---- 321=>x"c600", 322=>x"be00", 323=>x"bf00", 324=>x"c200",
---- 325=>x"c000", 326=>x"bf00", 327=>x"c200", 328=>x"bd00",
---- 329=>x"c100", 330=>x"c300", 331=>x"c300", 332=>x"be00",
---- 333=>x"c200", 334=>x"c300", 335=>x"c600", 336=>x"c200",
---- 337=>x"c300", 338=>x"c200", 339=>x"c700", 340=>x"c300",
---- 341=>x"c300", 342=>x"c600", 343=>x"c700", 344=>x"c600",
---- 345=>x"c600", 346=>x"c800", 347=>x"c600", 348=>x"c800",
---- 349=>x"c900", 350=>x"c900", 351=>x"c900", 352=>x"c700",
---- 353=>x"c900", 354=>x"c900", 355=>x"ca00", 356=>x"c700",
---- 357=>x"c800", 358=>x"c800", 359=>x"c900", 360=>x"c900",
---- 361=>x"c900", 362=>x"c700", 363=>x"c800", 364=>x"c800",
---- 365=>x"c800", 366=>x"c800", 367=>x"c300", 368=>x"c700",
---- 369=>x"c900", 370=>x"cb00", 371=>x"c800", 372=>x"c800",
---- 373=>x"cc00", 374=>x"ca00", 375=>x"c900", 376=>x"c600",
---- 377=>x"c600", 378=>x"c400", 379=>x"cd00", 380=>x"c700",
---- 381=>x"cb00", 382=>x"c900", 383=>x"af00", 384=>x"ce00",
---- 385=>x"bc00", 386=>x"8100", 387=>x"5500", 388=>x"8100",
---- 389=>x"5900", 390=>x"5500", 391=>x"5000", 392=>x"2d00",
---- 393=>x"bf00", 394=>x"7900", 395=>x"6700", 396=>x"5b00",
---- 397=>x"3f00", 398=>x"8100", 399=>x"8400", 400=>x"7700",
---- 401=>x"4d00", 402=>x"5c00", 403=>x"9300", 404=>x"6000",
---- 405=>x"7100", 406=>x"5600", 407=>x"7100", 408=>x"4f00",
---- 409=>x"5b00", 410=>x"6300", 411=>x"5600", 412=>x"7300",
---- 413=>x"6300", 414=>x"6400", 415=>x"6400", 416=>x"5800",
---- 417=>x"8400", 418=>x"6c00", 419=>x"5f00", 420=>x"4800",
---- 421=>x"4b00", 422=>x"7400", 423=>x"5500", 424=>x"4d00",
---- 425=>x"3700", 426=>x"4a00", 427=>x"6f00", 428=>x"5400",
---- 429=>x"4200", 430=>x"2700", 431=>x"4500", 432=>x"5200",
---- 433=>x"4300", 434=>x"3000", 435=>x"2b00", 436=>x"5500",
---- 437=>x"4000", 438=>x"2f00", 439=>x"2c00", 440=>x"5a00",
---- 441=>x"4600", 442=>x"2800", 443=>x"2b00", 444=>x"5e00",
---- 445=>x"4d00", 446=>x"2c00", 447=>x"2a00", 448=>x"6500",
---- 449=>x"5400", 450=>x"3300", 451=>x"2400", 452=>x"6b00",
---- 453=>x"5600", 454=>x"3b00", 455=>x"2e00", 456=>x"7100",
---- 457=>x"5500", 458=>x"4100", 459=>x"2f00", 460=>x"7700",
---- 461=>x"5a00", 462=>x"4a00", 463=>x"2e00", 464=>x"7e00",
---- 465=>x"6300", 466=>x"4e00", 467=>x"3500", 468=>x"8a00",
---- 469=>x"6700", 470=>x"5600", 471=>x"3d00", 472=>x"9300",
---- 473=>x"6f00", 474=>x"a400", 475=>x"4b00", 476=>x"9c00",
---- 477=>x"7500", 478=>x"5f00", 479=>x"5000", 480=>x"a200",
---- 481=>x"7700", 482=>x"6000", 483=>x"af00", 484=>x"a700",
---- 485=>x"7f00", 486=>x"5b00", 487=>x"4400", 488=>x"a300",
---- 489=>x"7800", 490=>x"b600", 491=>x"3600", 492=>x"8400",
---- 493=>x"6200", 494=>x"4000", 495=>x"3500", 496=>x"6400",
---- 497=>x"4e00", 498=>x"3b00", 499=>x"3600", 500=>x"5d00",
---- 501=>x"5a00", 502=>x"5500", 503=>x"5300", 504=>x"8600",
---- 505=>x"7700", 506=>x"6c00", 507=>x"6200", 508=>x"7500",
---- 509=>x"5f00", 510=>x"5300", 511=>x"5000", 512=>x"4400",
---- 513=>x"4400", 514=>x"4700", 515=>x"4400", 516=>x"3600",
---- 517=>x"3800", 518=>x"3d00", 519=>x"4200", 520=>x"3900",
---- 521=>x"3c00", 522=>x"3600", 523=>x"3d00", 524=>x"3200",
---- 525=>x"3700", 526=>x"c700", 527=>x"3800", 528=>x"2800",
---- 529=>x"3200", 530=>x"3700", 531=>x"3800", 532=>x"2e00",
---- 533=>x"3500", 534=>x"2f00", 535=>x"3400", 536=>x"2f00",
---- 537=>x"2c00", 538=>x"d600", 539=>x"2e00", 540=>x"3300",
---- 541=>x"2f00", 542=>x"2b00", 543=>x"2f00", 544=>x"cc00",
---- 545=>x"3200", 546=>x"2f00", 547=>x"3300", 548=>x"3600",
---- 549=>x"4100", 550=>x"c900", 551=>x"3700", 552=>x"4d00",
---- 553=>x"4f00", 554=>x"3a00", 555=>x"3800", 556=>x"5500",
---- 557=>x"5200", 558=>x"3800", 559=>x"3600", 560=>x"5a00",
---- 561=>x"5400", 562=>x"3900", 563=>x"3700", 564=>x"6200",
---- 565=>x"5a00", 566=>x"3f00", 567=>x"3c00", 568=>x"6c00",
---- 569=>x"5c00", 570=>x"4300", 571=>x"3f00", 572=>x"6e00",
---- 573=>x"6100", 574=>x"4500", 575=>x"3e00", 576=>x"6e00",
---- 577=>x"6400", 578=>x"4800", 579=>x"3900", 580=>x"7400",
---- 581=>x"6800", 582=>x"4c00", 583=>x"3900", 584=>x"7600",
---- 585=>x"6900", 586=>x"4700", 587=>x"3a00", 588=>x"7900",
---- 589=>x"6900", 590=>x"4500", 591=>x"3a00", 592=>x"7700",
---- 593=>x"6400", 594=>x"3f00", 595=>x"3700", 596=>x"7400",
---- 597=>x"5e00", 598=>x"3e00", 599=>x"3a00", 600=>x"7400",
---- 601=>x"5600", 602=>x"3e00", 603=>x"3700", 604=>x"6f00",
---- 605=>x"5000", 606=>x"3a00", 607=>x"2a00", 608=>x"6d00",
---- 609=>x"4a00", 610=>x"3500", 611=>x"2c00", 612=>x"6500",
---- 613=>x"4200", 614=>x"2f00", 615=>x"2a00", 616=>x"5b00",
---- 617=>x"4000", 618=>x"2b00", 619=>x"2e00", 620=>x"5700",
---- 621=>x"3300", 622=>x"2600", 623=>x"3200", 624=>x"4c00",
---- 625=>x"2d00", 626=>x"2b00", 627=>x"3000", 628=>x"3a00",
---- 629=>x"2800", 630=>x"2b00", 631=>x"3000", 632=>x"2f00",
---- 633=>x"2b00", 634=>x"2c00", 635=>x"3500", 636=>x"2700",
---- 637=>x"2b00", 638=>x"2a00", 639=>x"ce00", 640=>x"2700",
---- 641=>x"2b00", 642=>x"2d00", 643=>x"3400", 644=>x"2c00",
---- 645=>x"2d00", 646=>x"2f00", 647=>x"3700", 648=>x"2f00",
---- 649=>x"2b00", 650=>x"3100", 651=>x"3600", 652=>x"3400",
---- 653=>x"2a00", 654=>x"3100", 655=>x"3700", 656=>x"3200",
---- 657=>x"2d00", 658=>x"3200", 659=>x"3900", 660=>x"2f00",
---- 661=>x"2e00", 662=>x"3500", 663=>x"3900", 664=>x"2e00",
---- 665=>x"3000", 666=>x"3200", 667=>x"3f00", 668=>x"2f00",
---- 669=>x"2f00", 670=>x"3b00", 671=>x"4600", 672=>x"2e00",
---- 673=>x"2f00", 674=>x"3e00", 675=>x"4500", 676=>x"2d00",
---- 677=>x"3100", 678=>x"3f00", 679=>x"4000", 680=>x"2f00",
---- 681=>x"3200", 682=>x"4100", 683=>x"3c00", 684=>x"2f00",
---- 685=>x"3900", 686=>x"3a00", 687=>x"bf00", 688=>x"3200",
---- 689=>x"3600", 690=>x"3c00", 691=>x"4500", 692=>x"3500",
---- 693=>x"3500", 694=>x"4300", 695=>x"4300", 696=>x"3500",
---- 697=>x"3300", 698=>x"4900", 699=>x"3e00", 700=>x"3600",
---- 701=>x"3c00", 702=>x"4900", 703=>x"3b00", 704=>x"3500",
---- 705=>x"4300", 706=>x"4100", 707=>x"3600", 708=>x"3b00",
---- 709=>x"4400", 710=>x"3800", 711=>x"3c00", 712=>x"3600",
---- 713=>x"3500", 714=>x"3300", 715=>x"4100", 716=>x"4100",
---- 717=>x"3000", 718=>x"2d00", 719=>x"4100", 720=>x"4000",
---- 721=>x"3100", 722=>x"2f00", 723=>x"4500", 724=>x"3f00",
---- 725=>x"3400", 726=>x"3000", 727=>x"4800", 728=>x"3900",
---- 729=>x"3400", 730=>x"2f00", 731=>x"5300", 732=>x"3500",
---- 733=>x"3800", 734=>x"2c00", 735=>x"5700", 736=>x"3200",
---- 737=>x"3500", 738=>x"2a00", 739=>x"5300", 740=>x"3100",
---- 741=>x"3400", 742=>x"2c00", 743=>x"5800", 744=>x"3100",
---- 745=>x"3300", 746=>x"2f00", 747=>x"6000", 748=>x"2f00",
---- 749=>x"3200", 750=>x"3600", 751=>x"6000", 752=>x"2e00",
---- 753=>x"3300", 754=>x"3b00", 755=>x"6400", 756=>x"3000",
---- 757=>x"cc00", 758=>x"3800", 759=>x"6200", 760=>x"3300",
---- 761=>x"3400", 762=>x"4000", 763=>x"6800", 764=>x"3700",
---- 765=>x"3400", 766=>x"4300", 767=>x"6700", 768=>x"3400",
---- 769=>x"3900", 770=>x"4300", 771=>x"6500", 772=>x"3100",
---- 773=>x"3e00", 774=>x"4100", 775=>x"6300", 776=>x"3000",
---- 777=>x"3e00", 778=>x"3d00", 779=>x"6100", 780=>x"3200",
---- 781=>x"3f00", 782=>x"3e00", 783=>x"5f00", 784=>x"3200",
---- 785=>x"3e00", 786=>x"4900", 787=>x"5900", 788=>x"3500",
---- 789=>x"4000", 790=>x"5400", 791=>x"6100", 792=>x"2e00",
---- 793=>x"3900", 794=>x"5000", 795=>x"5600", 796=>x"2900",
---- 797=>x"3700", 798=>x"4d00", 799=>x"5000", 800=>x"2800",
---- 801=>x"3900", 802=>x"4b00", 803=>x"5400", 804=>x"2600",
---- 805=>x"3c00", 806=>x"4100", 807=>x"4a00", 808=>x"2700",
---- 809=>x"3400", 810=>x"3500", 811=>x"3f00", 812=>x"4f00",
---- 813=>x"2e00", 814=>x"d000", 815=>x"3500", 816=>x"b400",
---- 817=>x"5500", 818=>x"2900", 819=>x"3300", 820=>x"db00",
---- 821=>x"b800", 822=>x"4f00", 823=>x"3000", 824=>x"d800",
---- 825=>x"dc00", 826=>x"ab00", 827=>x"4200", 828=>x"d800",
---- 829=>x"d800", 830=>x"dd00", 831=>x"9c00", 832=>x"d800",
---- 833=>x"d900", 834=>x"db00", 835=>x"da00", 836=>x"2900",
---- 837=>x"d900", 838=>x"da00", 839=>x"df00", 840=>x"d700",
---- 841=>x"d800", 842=>x"db00", 843=>x"dd00", 844=>x"d500",
---- 845=>x"d500", 846=>x"db00", 847=>x"de00", 848=>x"d500",
---- 849=>x"d700", 850=>x"da00", 851=>x"2400", 852=>x"d500",
---- 853=>x"d600", 854=>x"d700", 855=>x"dc00", 856=>x"d500",
---- 857=>x"d300", 858=>x"d800", 859=>x"db00", 860=>x"d500",
---- 861=>x"d400", 862=>x"d600", 863=>x"d900", 864=>x"d400",
---- 865=>x"d400", 866=>x"d500", 867=>x"d900", 868=>x"d100",
---- 869=>x"d600", 870=>x"d600", 871=>x"d900", 872=>x"d100",
---- 873=>x"d500", 874=>x"d400", 875=>x"d600", 876=>x"d100",
---- 877=>x"d300", 878=>x"d400", 879=>x"d500", 880=>x"d100",
---- 881=>x"d300", 882=>x"d400", 883=>x"d400", 884=>x"d000",
---- 885=>x"d200", 886=>x"2b00", 887=>x"d400", 888=>x"cf00",
---- 889=>x"d300", 890=>x"d400", 891=>x"d400", 892=>x"cf00",
---- 893=>x"d100", 894=>x"d200", 895=>x"d300", 896=>x"cf00",
---- 897=>x"d100", 898=>x"d100", 899=>x"d300", 900=>x"cf00",
---- 901=>x"cd00", 902=>x"d000", 903=>x"d200", 904=>x"cd00",
---- 905=>x"ce00", 906=>x"d000", 907=>x"d200", 908=>x"cf00",
---- 909=>x"cf00", 910=>x"cf00", 911=>x"d200", 912=>x"cd00",
---- 913=>x"2f00", 914=>x"d000", 915=>x"d300", 916=>x"cc00",
---- 917=>x"cf00", 918=>x"2d00", 919=>x"d100", 920=>x"cb00",
---- 921=>x"cd00", 922=>x"d000", 923=>x"d300", 924=>x"ca00",
---- 925=>x"cd00", 926=>x"d100", 927=>x"d200", 928=>x"cc00",
---- 929=>x"ce00", 930=>x"d000", 931=>x"d000", 932=>x"ca00",
---- 933=>x"cc00", 934=>x"cf00", 935=>x"d000", 936=>x"cb00",
---- 937=>x"cb00", 938=>x"ce00", 939=>x"cf00", 940=>x"c800",
---- 941=>x"c900", 942=>x"cf00", 943=>x"ce00", 944=>x"c500",
---- 945=>x"c900", 946=>x"cb00", 947=>x"cd00", 948=>x"c400",
---- 949=>x"c700", 950=>x"ca00", 951=>x"ce00", 952=>x"c400",
---- 953=>x"c600", 954=>x"c900", 955=>x"cb00", 956=>x"c500",
---- 957=>x"c700", 958=>x"c700", 959=>x"cb00", 960=>x"c200",
---- 961=>x"c400", 962=>x"c800", 963=>x"cb00", 964=>x"c000",
---- 965=>x"c200", 966=>x"c600", 967=>x"c900", 968=>x"bf00",
---- 969=>x"c000", 970=>x"c300", 971=>x"c700", 972=>x"bd00",
---- 973=>x"be00", 974=>x"c200", 975=>x"c500", 976=>x"b900",
---- 977=>x"be00", 978=>x"c100", 979=>x"c400", 980=>x"b900",
---- 981=>x"bd00", 982=>x"c000", 983=>x"c200", 984=>x"b700",
---- 985=>x"ba00", 986=>x"be00", 987=>x"bf00", 988=>x"b900",
---- 989=>x"bb00", 990=>x"bd00", 991=>x"bf00", 992=>x"b600",
---- 993=>x"ba00", 994=>x"bc00", 995=>x"bd00", 996=>x"b300",
---- 997=>x"b300", 998=>x"ba00", 999=>x"bb00", 1000=>x"b400",
---- 1001=>x"b300", 1002=>x"b800", 1003=>x"bb00", 1004=>x"b400",
---- 1005=>x"b500", 1006=>x"b600", 1007=>x"ba00", 1008=>x"b100",
---- 1009=>x"b200", 1010=>x"b600", 1011=>x"b900", 1012=>x"ae00",
---- 1013=>x"b200", 1014=>x"b800", 1015=>x"4400", 1016=>x"ad00",
---- 1017=>x"b100", 1018=>x"b500", 1019=>x"b900", 1020=>x"ae00",
---- 1021=>x"5100", 1022=>x"b100", 1023=>x"b600"),
----
---- 44 => (0=>x"9a00", 1=>x"9a00", 2=>x"9c00", 3=>x"9a00", 4=>x"9900",
---- 5=>x"9c00", 6=>x"9b00", 7=>x"9a00", 8=>x"9900",
---- 9=>x"9a00", 10=>x"9b00", 11=>x"9b00", 12=>x"9500",
---- 13=>x"9900", 14=>x"9900", 15=>x"9800", 16=>x"9900",
---- 17=>x"9c00", 18=>x"9b00", 19=>x"9a00", 20=>x"9a00",
---- 21=>x"9d00", 22=>x"9e00", 23=>x"9d00", 24=>x"9b00",
---- 25=>x"9d00", 26=>x"a000", 27=>x"9e00", 28=>x"9e00",
---- 29=>x"a100", 30=>x"a000", 31=>x"a200", 32=>x"9e00",
---- 33=>x"a000", 34=>x"a100", 35=>x"a200", 36=>x"a200",
---- 37=>x"9f00", 38=>x"a100", 39=>x"a300", 40=>x"a300",
---- 41=>x"9f00", 42=>x"a100", 43=>x"a300", 44=>x"a100",
---- 45=>x"a100", 46=>x"a000", 47=>x"a100", 48=>x"a200",
---- 49=>x"a500", 50=>x"a000", 51=>x"9e00", 52=>x"a200",
---- 53=>x"a300", 54=>x"a000", 55=>x"9e00", 56=>x"a200",
---- 57=>x"a100", 58=>x"a100", 59=>x"a000", 60=>x"a000",
---- 61=>x"a000", 62=>x"9f00", 63=>x"9c00", 64=>x"a000",
---- 65=>x"a200", 66=>x"9e00", 67=>x"9d00", 68=>x"9f00",
---- 69=>x"a100", 70=>x"9f00", 71=>x"9e00", 72=>x"6300",
---- 73=>x"9e00", 74=>x"9d00", 75=>x"9d00", 76=>x"9c00",
---- 77=>x"9e00", 78=>x"9d00", 79=>x"a000", 80=>x"9900",
---- 81=>x"9e00", 82=>x"9a00", 83=>x"9e00", 84=>x"9a00",
---- 85=>x"9a00", 86=>x"9b00", 87=>x"9d00", 88=>x"9800",
---- 89=>x"9700", 90=>x"9a00", 91=>x"9c00", 92=>x"9600",
---- 93=>x"9500", 94=>x"9900", 95=>x"9c00", 96=>x"9500",
---- 97=>x"9600", 98=>x"9800", 99=>x"9a00", 100=>x"9000",
---- 101=>x"9600", 102=>x"9500", 103=>x"9700", 104=>x"9200",
---- 105=>x"9400", 106=>x"9400", 107=>x"9700", 108=>x"9300",
---- 109=>x"9400", 110=>x"9400", 111=>x"9600", 112=>x"9100",
---- 113=>x"9500", 114=>x"9400", 115=>x"9400", 116=>x"9100",
---- 117=>x"9300", 118=>x"9300", 119=>x"9400", 120=>x"8f00",
---- 121=>x"9200", 122=>x"9400", 123=>x"9400", 124=>x"8f00",
---- 125=>x"9200", 126=>x"9400", 127=>x"9300", 128=>x"9100",
---- 129=>x"9200", 130=>x"9100", 131=>x"9200", 132=>x"9100",
---- 133=>x"9000", 134=>x"9000", 135=>x"9000", 136=>x"9200",
---- 137=>x"9000", 138=>x"8f00", 139=>x"8f00", 140=>x"9600",
---- 141=>x"9300", 142=>x"9300", 143=>x"8d00", 144=>x"9700",
---- 145=>x"9400", 146=>x"9200", 147=>x"8e00", 148=>x"9700",
---- 149=>x"9400", 150=>x"9500", 151=>x"8f00", 152=>x"9700",
---- 153=>x"9800", 154=>x"9700", 155=>x"8e00", 156=>x"9800",
---- 157=>x"9800", 158=>x"9900", 159=>x"9200", 160=>x"9900",
---- 161=>x"9800", 162=>x"9900", 163=>x"9200", 164=>x"6600",
---- 165=>x"9a00", 166=>x"9a00", 167=>x"9200", 168=>x"9700",
---- 169=>x"9900", 170=>x"9800", 171=>x"9100", 172=>x"9900",
---- 173=>x"9b00", 174=>x"9800", 175=>x"9200", 176=>x"9800",
---- 177=>x"9800", 178=>x"9800", 179=>x"9300", 180=>x"9700",
---- 181=>x"9800", 182=>x"9800", 183=>x"9700", 184=>x"9b00",
---- 185=>x"9a00", 186=>x"9a00", 187=>x"9500", 188=>x"9a00",
---- 189=>x"9b00", 190=>x"9a00", 191=>x"9500", 192=>x"9800",
---- 193=>x"9a00", 194=>x"9800", 195=>x"9600", 196=>x"9900",
---- 197=>x"9900", 198=>x"9900", 199=>x"9700", 200=>x"9800",
---- 201=>x"9900", 202=>x"9b00", 203=>x"a100", 204=>x"9800",
---- 205=>x"9a00", 206=>x"9c00", 207=>x"9800", 208=>x"9900",
---- 209=>x"9900", 210=>x"9b00", 211=>x"9900", 212=>x"9a00",
---- 213=>x"9900", 214=>x"9900", 215=>x"9700", 216=>x"9a00",
---- 217=>x"9a00", 218=>x"9900", 219=>x"9600", 220=>x"9b00",
---- 221=>x"9a00", 222=>x"9900", 223=>x"9600", 224=>x"6600",
---- 225=>x"9900", 226=>x"9b00", 227=>x"9b00", 228=>x"9a00",
---- 229=>x"9900", 230=>x"9800", 231=>x"9a00", 232=>x"9a00",
---- 233=>x"9c00", 234=>x"9800", 235=>x"9a00", 236=>x"9800",
---- 237=>x"9b00", 238=>x"9900", 239=>x"9800", 240=>x"9900",
---- 241=>x"9a00", 242=>x"9a00", 243=>x"9800", 244=>x"9b00",
---- 245=>x"9b00", 246=>x"9800", 247=>x"9800", 248=>x"9d00",
---- 249=>x"9c00", 250=>x"9b00", 251=>x"9700", 252=>x"9d00",
---- 253=>x"9b00", 254=>x"9b00", 255=>x"9500", 256=>x"9a00",
---- 257=>x"9c00", 258=>x"9900", 259=>x"9200", 260=>x"9b00",
---- 261=>x"9a00", 262=>x"9400", 263=>x"9200", 264=>x"9a00",
---- 265=>x"9700", 266=>x"9400", 267=>x"8f00", 268=>x"9600",
---- 269=>x"9600", 270=>x"9000", 271=>x"8700", 272=>x"9600",
---- 273=>x"9400", 274=>x"8b00", 275=>x"8700", 276=>x"8e00",
---- 277=>x"8d00", 278=>x"9a00", 279=>x"bb00", 280=>x"9300",
---- 281=>x"ab00", 282=>x"c900", 283=>x"d600", 284=>x"c100",
---- 285=>x"d200", 286=>x"cd00", 287=>x"c400", 288=>x"d100",
---- 289=>x"be00", 290=>x"b800", 291=>x"bf00", 292=>x"c000",
---- 293=>x"bb00", 294=>x"be00", 295=>x"be00", 296=>x"c300",
---- 297=>x"c300", 298=>x"c600", 299=>x"ce00", 300=>x"c400",
---- 301=>x"c600", 302=>x"cf00", 303=>x"d300", 304=>x"cb00",
---- 305=>x"cf00", 306=>x"cf00", 307=>x"ce00", 308=>x"cf00",
---- 309=>x"cb00", 310=>x"cb00", 311=>x"ca00", 312=>x"c600",
---- 313=>x"c400", 314=>x"c400", 315=>x"c300", 316=>x"c000",
---- 317=>x"bc00", 318=>x"c000", 319=>x"c000", 320=>x"c300",
---- 321=>x"c100", 322=>x"be00", 323=>x"c200", 324=>x"c200",
---- 325=>x"c000", 326=>x"bf00", 327=>x"c500", 328=>x"c200",
---- 329=>x"c300", 330=>x"c300", 331=>x"c700", 332=>x"c300",
---- 333=>x"3b00", 334=>x"c700", 335=>x"c900", 336=>x"c400",
---- 337=>x"c600", 338=>x"ca00", 339=>x"cb00", 340=>x"c700",
---- 341=>x"c900", 342=>x"cd00", 343=>x"ca00", 344=>x"c700",
---- 345=>x"ca00", 346=>x"c900", 347=>x"cd00", 348=>x"c900",
---- 349=>x"cb00", 350=>x"cb00", 351=>x"cd00", 352=>x"c900",
---- 353=>x"ca00", 354=>x"cc00", 355=>x"ce00", 356=>x"c700",
---- 357=>x"cb00", 358=>x"ce00", 359=>x"cd00", 360=>x"c600",
---- 361=>x"cd00", 362=>x"d000", 363=>x"cc00", 364=>x"c300",
---- 365=>x"d000", 366=>x"cc00", 367=>x"cc00", 368=>x"cb00",
---- 369=>x"cf00", 370=>x"d000", 371=>x"d500", 372=>x"ce00",
---- 373=>x"d500", 374=>x"cf00", 375=>x"a600", 376=>x"c900",
---- 377=>x"ad00", 378=>x"9600", 379=>x"7700", 380=>x"7f00",
---- 381=>x"5d00", 382=>x"8100", 383=>x"8600", 384=>x"6600",
---- 385=>x"6900", 386=>x"8400", 387=>x"8c00", 388=>x"6a00",
---- 389=>x"6700", 390=>x"7a00", 391=>x"8d00", 392=>x"6500",
---- 393=>x"6a00", 394=>x"6c00", 395=>x"8d00", 396=>x"6800",
---- 397=>x"7700", 398=>x"6a00", 399=>x"8600", 400=>x"7200",
---- 401=>x"7800", 402=>x"7800", 403=>x"7600", 404=>x"8c00",
---- 405=>x"7200", 406=>x"7f00", 407=>x"6b00", 408=>x"7f00",
---- 409=>x"8100", 410=>x"7500", 411=>x"6a00", 412=>x"7400",
---- 413=>x"8b00", 414=>x"7b00", 415=>x"7800", 416=>x"5900",
---- 417=>x"8000", 418=>x"8900", 419=>x"8300", 420=>x"4900",
---- 421=>x"5300", 422=>x"8b00", 423=>x"8700", 424=>x"5b00",
---- 425=>x"4500", 426=>x"6e00", 427=>x"8a00", 428=>x"6300",
---- 429=>x"4a00", 430=>x"5100", 431=>x"8300", 432=>x"5e00",
---- 433=>x"5600", 434=>x"b300", 435=>x"7700", 436=>x"c600",
---- 437=>x"5600", 438=>x"b800", 439=>x"6300", 440=>x"2900",
---- 441=>x"5100", 442=>x"4900", 443=>x"5100", 444=>x"2e00",
---- 445=>x"3f00", 446=>x"4c00", 447=>x"4700", 448=>x"2a00",
---- 449=>x"3200", 450=>x"4a00", 451=>x"4300", 452=>x"2800",
---- 453=>x"2900", 454=>x"3a00", 455=>x"4500", 456=>x"2400",
---- 457=>x"2500", 458=>x"2e00", 459=>x"4800", 460=>x"2200",
---- 461=>x"2400", 462=>x"2800", 463=>x"4700", 464=>x"2700",
---- 465=>x"2600", 466=>x"2900", 467=>x"3800", 468=>x"2d00",
---- 469=>x"2b00", 470=>x"2900", 471=>x"3000", 472=>x"3100",
---- 473=>x"2c00", 474=>x"2800", 475=>x"2700", 476=>x"3300",
---- 477=>x"2700", 478=>x"2900", 479=>x"2700", 480=>x"3100",
---- 481=>x"2600", 482=>x"2b00", 483=>x"2900", 484=>x"3000",
---- 485=>x"2700", 486=>x"2800", 487=>x"d600", 488=>x"2f00",
---- 489=>x"2a00", 490=>x"2700", 491=>x"2700", 492=>x"2d00",
---- 493=>x"2700", 494=>x"2600", 495=>x"2600", 496=>x"2c00",
---- 497=>x"2700", 498=>x"2900", 499=>x"2900", 500=>x"3700",
---- 501=>x"2c00", 502=>x"2d00", 503=>x"2a00", 504=>x"4000",
---- 505=>x"3400", 506=>x"2d00", 507=>x"2700", 508=>x"3d00",
---- 509=>x"4200", 510=>x"3000", 511=>x"2c00", 512=>x"4500",
---- 513=>x"4000", 514=>x"2b00", 515=>x"2700", 516=>x"4600",
---- 517=>x"2f00", 518=>x"2c00", 519=>x"2700", 520=>x"3900",
---- 521=>x"2c00", 522=>x"2d00", 523=>x"2800", 524=>x"2e00",
---- 525=>x"3100", 526=>x"3100", 527=>x"2800", 528=>x"3000",
---- 529=>x"3000", 530=>x"3100", 531=>x"2500", 532=>x"3100",
---- 533=>x"2f00", 534=>x"3200", 535=>x"2f00", 536=>x"2f00",
---- 537=>x"2c00", 538=>x"3100", 539=>x"2f00", 540=>x"2a00",
---- 541=>x"2d00", 542=>x"2800", 543=>x"2600", 544=>x"cc00",
---- 545=>x"2c00", 546=>x"3000", 547=>x"2d00", 548=>x"3600",
---- 549=>x"3000", 550=>x"3800", 551=>x"3100", 552=>x"3600",
---- 553=>x"2d00", 554=>x"3c00", 555=>x"3300", 556=>x"3400",
---- 557=>x"2900", 558=>x"3300", 559=>x"3400", 560=>x"2f00",
---- 561=>x"2900", 562=>x"3400", 563=>x"3100", 564=>x"2e00",
---- 565=>x"2b00", 566=>x"3400", 567=>x"3400", 568=>x"3000",
---- 569=>x"2d00", 570=>x"3500", 571=>x"3600", 572=>x"3300",
---- 573=>x"2e00", 574=>x"3500", 575=>x"3c00", 576=>x"3200",
---- 577=>x"d200", 578=>x"3700", 579=>x"3900", 580=>x"3300",
---- 581=>x"3100", 582=>x"3b00", 583=>x"3700", 584=>x"3200",
---- 585=>x"3400", 586=>x"4000", 587=>x"3900", 588=>x"3200",
---- 589=>x"3500", 590=>x"3e00", 591=>x"3900", 592=>x"3100",
---- 593=>x"3700", 594=>x"3600", 595=>x"c600", 596=>x"2e00",
---- 597=>x"3800", 598=>x"3300", 599=>x"3b00", 600=>x"2c00",
---- 601=>x"3600", 602=>x"3000", 603=>x"3a00", 604=>x"3000",
---- 605=>x"3300", 606=>x"3100", 607=>x"3c00", 608=>x"3500",
---- 609=>x"3600", 610=>x"3800", 611=>x"4000", 612=>x"3600",
---- 613=>x"3c00", 614=>x"3a00", 615=>x"3d00", 616=>x"3200",
---- 617=>x"3b00", 618=>x"4300", 619=>x"4600", 620=>x"2f00",
---- 621=>x"3800", 622=>x"4200", 623=>x"4700", 624=>x"3400",
---- 625=>x"4000", 626=>x"4100", 627=>x"4300", 628=>x"3000",
---- 629=>x"3b00", 630=>x"4500", 631=>x"4a00", 632=>x"2e00",
---- 633=>x"3c00", 634=>x"4700", 635=>x"4a00", 636=>x"3200",
---- 637=>x"3e00", 638=>x"4500", 639=>x"4800", 640=>x"3200",
---- 641=>x"3b00", 642=>x"4600", 643=>x"4300", 644=>x"3600",
---- 645=>x"3e00", 646=>x"4a00", 647=>x"3e00", 648=>x"3300",
---- 649=>x"4400", 650=>x"b600", 651=>x"3f00", 652=>x"c800",
---- 653=>x"4500", 654=>x"4b00", 655=>x"3c00", 656=>x"3700",
---- 657=>x"4b00", 658=>x"5300", 659=>x"4000", 660=>x"3b00",
---- 661=>x"5100", 662=>x"5200", 663=>x"4800", 664=>x"3900",
---- 665=>x"5c00", 666=>x"4900", 667=>x"4b00", 668=>x"3900",
---- 669=>x"5b00", 670=>x"4900", 671=>x"4700", 672=>x"3e00",
---- 673=>x"5b00", 674=>x"4400", 675=>x"4600", 676=>x"4200",
---- 677=>x"5700", 678=>x"4600", 679=>x"4600", 680=>x"4a00",
---- 681=>x"5500", 682=>x"4800", 683=>x"4800", 684=>x"4a00",
---- 685=>x"5000", 686=>x"4800", 687=>x"4800", 688=>x"b300",
---- 689=>x"5300", 690=>x"4700", 691=>x"4700", 692=>x"4600",
---- 693=>x"5500", 694=>x"4c00", 695=>x"4b00", 696=>x"4500",
---- 697=>x"4d00", 698=>x"4900", 699=>x"5200", 700=>x"4d00",
---- 701=>x"4800", 702=>x"4600", 703=>x"5200", 704=>x"4f00",
---- 705=>x"4c00", 706=>x"4800", 707=>x"5200", 708=>x"5400",
---- 709=>x"4800", 710=>x"4c00", 711=>x"5200", 712=>x"5900",
---- 713=>x"4600", 714=>x"4b00", 715=>x"4f00", 716=>x"6000",
---- 717=>x"4700", 718=>x"5300", 719=>x"5400", 720=>x"5d00",
---- 721=>x"4100", 722=>x"4f00", 723=>x"5900", 724=>x"5900",
---- 725=>x"3f00", 726=>x"5000", 727=>x"5400", 728=>x"5700",
---- 729=>x"4600", 730=>x"5000", 731=>x"5300", 732=>x"5e00",
---- 733=>x"4400", 734=>x"5000", 735=>x"5d00", 736=>x"5e00",
---- 737=>x"4900", 738=>x"5000", 739=>x"5900", 740=>x"6100",
---- 741=>x"4400", 742=>x"4e00", 743=>x"5700", 744=>x"6200",
---- 745=>x"4600", 746=>x"5400", 747=>x"5400", 748=>x"6200",
---- 749=>x"4900", 750=>x"5700", 751=>x"5c00", 752=>x"6800",
---- 753=>x"4a00", 754=>x"5500", 755=>x"5b00", 756=>x"6900",
---- 757=>x"4900", 758=>x"5900", 759=>x"5800", 760=>x"6300",
---- 761=>x"4700", 762=>x"5900", 763=>x"5400", 764=>x"6400",
---- 765=>x"5000", 766=>x"5700", 767=>x"5500", 768=>x"6500",
---- 769=>x"5300", 770=>x"5600", 771=>x"5700", 772=>x"6800",
---- 773=>x"5400", 774=>x"5a00", 775=>x"5700", 776=>x"6800",
---- 777=>x"5100", 778=>x"5c00", 779=>x"5900", 780=>x"6a00",
---- 781=>x"4f00", 782=>x"5a00", 783=>x"5a00", 784=>x"6a00",
---- 785=>x"4e00", 786=>x"5600", 787=>x"5800", 788=>x"6b00",
---- 789=>x"4f00", 790=>x"5300", 791=>x"5900", 792=>x"6900",
---- 793=>x"4e00", 794=>x"5100", 795=>x"5400", 796=>x"6600",
---- 797=>x"4b00", 798=>x"4f00", 799=>x"5500", 800=>x"9b00",
---- 801=>x"4d00", 802=>x"4d00", 803=>x"5200", 804=>x"6500",
---- 805=>x"4b00", 806=>x"4800", 807=>x"4e00", 808=>x"6600",
---- 809=>x"4a00", 810=>x"4600", 811=>x"4e00", 812=>x"5d00",
---- 813=>x"4600", 814=>x"4100", 815=>x"4800", 816=>x"5300",
---- 817=>x"4000", 818=>x"3700", 819=>x"4400", 820=>x"af00",
---- 821=>x"4500", 822=>x"3b00", 823=>x"3d00", 824=>x"3800",
---- 825=>x"4000", 826=>x"3000", 827=>x"3800", 828=>x"3400",
---- 829=>x"3400", 830=>x"2c00", 831=>x"2f00", 832=>x"7d00",
---- 833=>x"3300", 834=>x"2d00", 835=>x"2b00", 836=>x"ca00",
---- 837=>x"5d00", 838=>x"2b00", 839=>x"2d00", 840=>x"df00",
---- 841=>x"aa00", 842=>x"3400", 843=>x"2500", 844=>x"dd00",
---- 845=>x"d900", 846=>x"6c00", 847=>x"2300", 848=>x"db00",
---- 849=>x"e200", 850=>x"b300", 851=>x"3500", 852=>x"dc00",
---- 853=>x"dc00", 854=>x"db00", 855=>x"6700", 856=>x"dc00",
---- 857=>x"dd00", 858=>x"e300", 859=>x"a700", 860=>x"db00",
---- 861=>x"dd00", 862=>x"df00", 863=>x"d500", 864=>x"d800",
---- 865=>x"dd00", 866=>x"dc00", 867=>x"e200", 868=>x"d700",
---- 869=>x"db00", 870=>x"dd00", 871=>x"e200", 872=>x"d800",
---- 873=>x"da00", 874=>x"dc00", 875=>x"de00", 876=>x"d700",
---- 877=>x"d800", 878=>x"da00", 879=>x"dc00", 880=>x"d500",
---- 881=>x"d700", 882=>x"da00", 883=>x"da00", 884=>x"d700",
---- 885=>x"d800", 886=>x"d800", 887=>x"da00", 888=>x"d500",
---- 889=>x"d700", 890=>x"d800", 891=>x"d900", 892=>x"d300",
---- 893=>x"d600", 894=>x"d600", 895=>x"da00", 896=>x"d500",
---- 897=>x"d500", 898=>x"d600", 899=>x"d600", 900=>x"d500",
---- 901=>x"d400", 902=>x"d700", 903=>x"d500", 904=>x"d200",
---- 905=>x"d600", 906=>x"d500", 907=>x"d600", 908=>x"d200",
---- 909=>x"d400", 910=>x"d400", 911=>x"d400", 912=>x"d600",
---- 913=>x"d300", 914=>x"d500", 915=>x"d300", 916=>x"d200",
---- 917=>x"d400", 918=>x"d500", 919=>x"d600", 920=>x"d300",
---- 921=>x"d300", 922=>x"d400", 923=>x"d600", 924=>x"d200",
---- 925=>x"d500", 926=>x"d600", 927=>x"d600", 928=>x"d200",
---- 929=>x"d500", 930=>x"2b00", 931=>x"d500", 932=>x"d100",
---- 933=>x"d400", 934=>x"d500", 935=>x"d400", 936=>x"d100",
---- 937=>x"d300", 938=>x"d300", 939=>x"d300", 940=>x"d000",
---- 941=>x"d100", 942=>x"d200", 943=>x"d400", 944=>x"ce00",
---- 945=>x"d000", 946=>x"d100", 947=>x"d400", 948=>x"d000",
---- 949=>x"d100", 950=>x"d000", 951=>x"d300", 952=>x"3100",
---- 953=>x"d000", 954=>x"d200", 955=>x"d300", 956=>x"cd00",
---- 957=>x"ce00", 958=>x"d000", 959=>x"d100", 960=>x"ce00",
---- 961=>x"d100", 962=>x"cf00", 963=>x"d000", 964=>x"cc00",
---- 965=>x"ce00", 966=>x"ce00", 967=>x"d100", 968=>x"c900",
---- 969=>x"cc00", 970=>x"cf00", 971=>x"d000", 972=>x"c800",
---- 973=>x"cb00", 974=>x"cd00", 975=>x"ce00", 976=>x"c800",
---- 977=>x"c800", 978=>x"cd00", 979=>x"ce00", 980=>x"c700",
---- 981=>x"c900", 982=>x"cc00", 983=>x"cc00", 984=>x"c400",
---- 985=>x"c800", 986=>x"cb00", 987=>x"ce00", 988=>x"c300",
---- 989=>x"c500", 990=>x"c900", 991=>x"cb00", 992=>x"c000",
---- 993=>x"c400", 994=>x"c600", 995=>x"c800", 996=>x"bd00",
---- 997=>x"c300", 998=>x"c300", 999=>x"c500", 1000=>x"bb00",
---- 1001=>x"c100", 1002=>x"c500", 1003=>x"c700", 1004=>x"ba00",
---- 1005=>x"bd00", 1006=>x"c600", 1007=>x"c700", 1008=>x"bc00",
---- 1009=>x"bd00", 1010=>x"c400", 1011=>x"c500", 1012=>x"b800",
---- 1013=>x"bc00", 1014=>x"c100", 1015=>x"c300", 1016=>x"bb00",
---- 1017=>x"bf00", 1018=>x"c100", 1019=>x"c400", 1020=>x"b900",
---- 1021=>x"bf00", 1022=>x"c000", 1023=>x"c200"),
----
---- 45 => (0=>x"9e00", 1=>x"9c00", 2=>x"9a00", 3=>x"9800", 4=>x"9e00",
---- 5=>x"9e00", 6=>x"9a00", 7=>x"9900", 8=>x"9c00",
---- 9=>x"9c00", 10=>x"9b00", 11=>x"9900", 12=>x"9900",
---- 13=>x"9b00", 14=>x"9b00", 15=>x"9900", 16=>x"9b00",
---- 17=>x"9b00", 18=>x"9a00", 19=>x"9c00", 20=>x"9f00",
---- 21=>x"9c00", 22=>x"9a00", 23=>x"6300", 24=>x"a000",
---- 25=>x"9f00", 26=>x"9f00", 27=>x"9e00", 28=>x"a200",
---- 29=>x"a200", 30=>x"a200", 31=>x"9e00", 32=>x"a100",
---- 33=>x"a200", 34=>x"a200", 35=>x"9f00", 36=>x"a400",
---- 37=>x"a000", 38=>x"a200", 39=>x"a300", 40=>x"a400",
---- 41=>x"a400", 42=>x"a200", 43=>x"a200", 44=>x"a000",
---- 45=>x"a200", 46=>x"a100", 47=>x"a100", 48=>x"a000",
---- 49=>x"a100", 50=>x"a000", 51=>x"a000", 52=>x"9e00",
---- 53=>x"9f00", 54=>x"9f00", 55=>x"9f00", 56=>x"9d00",
---- 57=>x"9e00", 58=>x"a000", 59=>x"9c00", 60=>x"a000",
---- 61=>x"9d00", 62=>x"a100", 63=>x"9e00", 64=>x"9f00",
---- 65=>x"9e00", 66=>x"a000", 67=>x"a000", 68=>x"9e00",
---- 69=>x"9d00", 70=>x"9f00", 71=>x"9e00", 72=>x"9c00",
---- 73=>x"9d00", 74=>x"9d00", 75=>x"9d00", 76=>x"9c00",
---- 77=>x"9d00", 78=>x"9d00", 79=>x"9d00", 80=>x"9d00",
---- 81=>x"9c00", 82=>x"9d00", 83=>x"9c00", 84=>x"9e00",
---- 85=>x"9900", 86=>x"9c00", 87=>x"9c00", 88=>x"9c00",
---- 89=>x"9c00", 90=>x"9b00", 91=>x"9800", 92=>x"9a00",
---- 93=>x"9b00", 94=>x"9a00", 95=>x"9a00", 96=>x"9a00",
---- 97=>x"9b00", 98=>x"9b00", 99=>x"9c00", 100=>x"9a00",
---- 101=>x"9a00", 102=>x"9a00", 103=>x"9b00", 104=>x"9700",
---- 105=>x"9a00", 106=>x"9a00", 107=>x"9a00", 108=>x"9700",
---- 109=>x"9800", 110=>x"9a00", 111=>x"9800", 112=>x"9900",
---- 113=>x"9800", 114=>x"9900", 115=>x"9700", 116=>x"9300",
---- 117=>x"9500", 118=>x"9700", 119=>x"9800", 120=>x"9000",
---- 121=>x"9200", 122=>x"9700", 123=>x"9a00", 124=>x"9300",
---- 125=>x"9200", 126=>x"9400", 127=>x"9500", 128=>x"9200",
---- 129=>x"9100", 130=>x"9200", 131=>x"9300", 132=>x"8f00",
---- 133=>x"9000", 134=>x"9000", 135=>x"8e00", 136=>x"8e00",
---- 137=>x"9000", 138=>x"8e00", 139=>x"8c00", 140=>x"8a00",
---- 141=>x"8c00", 142=>x"8c00", 143=>x"8b00", 144=>x"8800",
---- 145=>x"8500", 146=>x"8600", 147=>x"8600", 148=>x"8800",
---- 149=>x"8400", 150=>x"8100", 151=>x"7f00", 152=>x"8700",
---- 153=>x"8000", 154=>x"7a00", 155=>x"7600", 156=>x"8900",
---- 157=>x"7d00", 158=>x"7700", 159=>x"6c00", 160=>x"8b00",
---- 161=>x"7f00", 162=>x"7100", 163=>x"6400", 164=>x"8f00",
---- 165=>x"8300", 166=>x"7300", 167=>x"5e00", 168=>x"8d00",
---- 169=>x"8300", 170=>x"7500", 171=>x"5d00", 172=>x"8d00",
---- 173=>x"8500", 174=>x"7700", 175=>x"5c00", 176=>x"8f00",
---- 177=>x"8500", 178=>x"7a00", 179=>x"6400", 180=>x"9100",
---- 181=>x"8600", 182=>x"7a00", 183=>x"6600", 184=>x"9200",
---- 185=>x"8d00", 186=>x"7e00", 187=>x"6a00", 188=>x"8f00",
---- 189=>x"8700", 190=>x"7b00", 191=>x"6500", 192=>x"9200",
---- 193=>x"8900", 194=>x"7b00", 195=>x"6400", 196=>x"9300",
---- 197=>x"8900", 198=>x"7c00", 199=>x"6400", 200=>x"9100",
---- 201=>x"8700", 202=>x"7a00", 203=>x"6500", 204=>x"8f00",
---- 205=>x"8700", 206=>x"7700", 207=>x"6600", 208=>x"9000",
---- 209=>x"8800", 210=>x"7900", 211=>x"6700", 212=>x"9100",
---- 213=>x"8700", 214=>x"7d00", 215=>x"6c00", 216=>x"9000",
---- 217=>x"8600", 218=>x"7b00", 219=>x"6900", 220=>x"9000",
---- 221=>x"8600", 222=>x"7a00", 223=>x"6700", 224=>x"6d00",
---- 225=>x"8600", 226=>x"7b00", 227=>x"6b00", 228=>x"9400",
---- 229=>x"8700", 230=>x"8100", 231=>x"6700", 232=>x"9400",
---- 233=>x"8700", 234=>x"7900", 235=>x"6c00", 236=>x"9200",
---- 237=>x"8800", 238=>x"7800", 239=>x"6600", 240=>x"9300",
---- 241=>x"8800", 242=>x"7700", 243=>x"6500", 244=>x"9200",
---- 245=>x"8600", 246=>x"7a00", 247=>x"6500", 248=>x"9100",
---- 249=>x"8600", 250=>x"7500", 251=>x"6000", 252=>x"8f00",
---- 253=>x"8100", 254=>x"6e00", 255=>x"5f00", 256=>x"8c00",
---- 257=>x"7a00", 258=>x"6800", 259=>x"5300", 260=>x"8800",
---- 261=>x"7700", 262=>x"6000", 263=>x"4700", 264=>x"8400",
---- 265=>x"6e00", 266=>x"5500", 267=>x"6000", 268=>x"7c00",
---- 269=>x"7300", 270=>x"9100", 271=>x"c600", 272=>x"6200",
---- 273=>x"bb00", 274=>x"da00", 275=>x"d600", 276=>x"d700",
---- 277=>x"d700", 278=>x"c700", 279=>x"bc00", 280=>x"c900",
---- 281=>x"be00", 282=>x"ba00", 283=>x"ba00", 284=>x"c100",
---- 285=>x"bf00", 286=>x"bd00", 287=>x"bf00", 288=>x"bf00",
---- 289=>x"c400", 290=>x"c900", 291=>x"d000", 292=>x"c500",
---- 293=>x"cf00", 294=>x"d000", 295=>x"cd00", 296=>x"d200",
---- 297=>x"d100", 298=>x"cc00", 299=>x"c800", 300=>x"d100",
---- 301=>x"ce00", 302=>x"3b00", 303=>x"c100", 304=>x"cd00",
---- 305=>x"c600", 306=>x"c100", 307=>x"c700", 308=>x"c600",
---- 309=>x"c400", 310=>x"3a00", 311=>x"c900", 312=>x"c400",
---- 313=>x"c500", 314=>x"c400", 315=>x"c900", 316=>x"c400",
---- 317=>x"c300", 318=>x"c600", 319=>x"c800", 320=>x"c500",
---- 321=>x"c500", 322=>x"c900", 323=>x"c900", 324=>x"c600",
---- 325=>x"c800", 326=>x"c900", 327=>x"c900", 328=>x"c800",
---- 329=>x"ca00", 330=>x"c900", 331=>x"cc00", 332=>x"ca00",
---- 333=>x"cb00", 334=>x"cc00", 335=>x"cc00", 336=>x"cc00",
---- 337=>x"cc00", 338=>x"cb00", 339=>x"cb00", 340=>x"cc00",
---- 341=>x"ca00", 342=>x"cb00", 343=>x"cc00", 344=>x"cd00",
---- 345=>x"ca00", 346=>x"cc00", 347=>x"cc00", 348=>x"cb00",
---- 349=>x"3500", 350=>x"cc00", 351=>x"cc00", 352=>x"ca00",
---- 353=>x"ca00", 354=>x"cb00", 355=>x"cb00", 356=>x"cb00",
---- 357=>x"ce00", 358=>x"cc00", 359=>x"cb00", 360=>x"cc00",
---- 361=>x"cf00", 362=>x"d200", 363=>x"d200", 364=>x"d300",
---- 365=>x"d300", 366=>x"c000", 367=>x"9800", 368=>x"bf00",
---- 369=>x"8900", 370=>x"6900", 371=>x"5400", 372=>x"6800",
---- 373=>x"5300", 374=>x"5b00", 375=>x"5c00", 376=>x"5e00",
---- 377=>x"5e00", 378=>x"6100", 379=>x"5c00", 380=>x"7300",
---- 381=>x"6000", 382=>x"6000", 383=>x"5900", 384=>x"8100",
---- 385=>x"8c00", 386=>x"7200", 387=>x"7b00", 388=>x"9200",
---- 389=>x"9c00", 390=>x"9e00", 391=>x"a200", 392=>x"9900",
---- 393=>x"a700", 394=>x"a300", 395=>x"a500", 396=>x"9800",
---- 397=>x"a400", 398=>x"a000", 399=>x"a800", 400=>x"9500",
---- 401=>x"9700", 402=>x"9d00", 403=>x"ab00", 404=>x"8800",
---- 405=>x"9800", 406=>x"9a00", 407=>x"a700", 408=>x"7900",
---- 409=>x"9700", 410=>x"9800", 411=>x"a600", 412=>x"7a00",
---- 413=>x"9400", 414=>x"9c00", 415=>x"b000", 416=>x"7f00",
---- 417=>x"9000", 418=>x"a400", 419=>x"bb00", 420=>x"8200",
---- 421=>x"8a00", 422=>x"a200", 423=>x"9f00", 424=>x"8700",
---- 425=>x"8f00", 426=>x"9a00", 427=>x"8700", 428=>x"8500",
---- 429=>x"9300", 430=>x"9a00", 431=>x"8e00", 432=>x"8600",
---- 433=>x"8900", 434=>x"9700", 435=>x"9200", 436=>x"8e00",
---- 437=>x"8900", 438=>x"9900", 439=>x"9800", 440=>x"9200",
---- 441=>x"9200", 442=>x"a200", 443=>x"9c00", 444=>x"8b00",
---- 445=>x"9b00", 446=>x"a700", 447=>x"9900", 448=>x"6f00",
---- 449=>x"9f00", 450=>x"ac00", 451=>x"9c00", 452=>x"4f00",
---- 453=>x"9800", 454=>x"a400", 455=>x"a500", 456=>x"4400",
---- 457=>x"8d00", 458=>x"a600", 459=>x"a200", 460=>x"4400",
---- 461=>x"8200", 462=>x"ae00", 463=>x"6100", 464=>x"4700",
---- 465=>x"9500", 466=>x"b200", 467=>x"a000", 468=>x"4700",
---- 469=>x"5700", 470=>x"a800", 471=>x"aa00", 472=>x"4b00",
---- 473=>x"5500", 474=>x"9700", 475=>x"b100", 476=>x"4200",
---- 477=>x"5100", 478=>x"8d00", 479=>x"b500", 480=>x"3d00",
---- 481=>x"4a00", 482=>x"7b00", 483=>x"b600", 484=>x"3800",
---- 485=>x"4100", 486=>x"7100", 487=>x"b800", 488=>x"3200",
---- 489=>x"4300", 490=>x"6000", 491=>x"b800", 492=>x"3500",
---- 493=>x"4b00", 494=>x"4e00", 495=>x"b700", 496=>x"3400",
---- 497=>x"4200", 498=>x"3f00", 499=>x"ab00", 500=>x"3100",
---- 501=>x"3b00", 502=>x"4000", 503=>x"a800", 504=>x"2a00",
---- 505=>x"3d00", 506=>x"4000", 507=>x"a200", 508=>x"2d00",
---- 509=>x"4100", 510=>x"3a00", 511=>x"9700", 512=>x"2c00",
---- 513=>x"4500", 514=>x"3d00", 515=>x"9500", 516=>x"2500",
---- 517=>x"4700", 518=>x"3900", 519=>x"8d00", 520=>x"2900",
---- 521=>x"4200", 522=>x"3600", 523=>x"8600", 524=>x"2c00",
---- 525=>x"4400", 526=>x"3400", 527=>x"8100", 528=>x"2b00",
---- 529=>x"4700", 530=>x"3000", 531=>x"7b00", 532=>x"2e00",
---- 533=>x"4f00", 534=>x"2d00", 535=>x"7a00", 536=>x"3100",
---- 537=>x"5200", 538=>x"2a00", 539=>x"7400", 540=>x"3900",
---- 541=>x"5600", 542=>x"2900", 543=>x"6e00", 544=>x"3c00",
---- 545=>x"5100", 546=>x"2d00", 547=>x"6300", 548=>x"4000",
---- 549=>x"5200", 550=>x"2d00", 551=>x"6000", 552=>x"4200",
---- 553=>x"4a00", 554=>x"2800", 555=>x"5b00", 556=>x"4b00",
---- 557=>x"4c00", 558=>x"2c00", 559=>x"5800", 560=>x"4800",
---- 561=>x"b600", 562=>x"2a00", 563=>x"5700", 564=>x"4000",
---- 565=>x"4600", 566=>x"2a00", 567=>x"5400", 568=>x"4200",
---- 569=>x"4900", 570=>x"2c00", 571=>x"5100", 572=>x"4100",
---- 573=>x"4100", 574=>x"2900", 575=>x"4b00", 576=>x"4100",
---- 577=>x"4400", 578=>x"2200", 579=>x"4400", 580=>x"4700",
---- 581=>x"4200", 582=>x"2000", 583=>x"4100", 584=>x"4800",
---- 585=>x"3d00", 586=>x"2700", 587=>x"3800", 588=>x"4d00",
---- 589=>x"3d00", 590=>x"2600", 591=>x"3400", 592=>x"5500",
---- 593=>x"3b00", 594=>x"2700", 595=>x"3100", 596=>x"5600",
---- 597=>x"3600", 598=>x"2400", 599=>x"2d00", 600=>x"5600",
---- 601=>x"3500", 602=>x"2400", 603=>x"2900", 604=>x"5600",
---- 605=>x"3400", 606=>x"2600", 607=>x"2400", 608=>x"5700",
---- 609=>x"3100", 610=>x"2300", 611=>x"2200", 612=>x"5900",
---- 613=>x"3600", 614=>x"2300", 615=>x"2600", 616=>x"5500",
---- 617=>x"3800", 618=>x"2300", 619=>x"2600", 620=>x"4f00",
---- 621=>x"3800", 622=>x"1e00", 623=>x"2300", 624=>x"4e00",
---- 625=>x"3800", 626=>x"2200", 627=>x"2200", 628=>x"4400",
---- 629=>x"3d00", 630=>x"2500", 631=>x"2400", 632=>x"4700",
---- 633=>x"3800", 634=>x"2500", 635=>x"2500", 636=>x"4700",
---- 637=>x"3500", 638=>x"2a00", 639=>x"2700", 640=>x"4700",
---- 641=>x"3100", 642=>x"2e00", 643=>x"2b00", 644=>x"ba00",
---- 645=>x"3200", 646=>x"3000", 647=>x"2b00", 648=>x"4a00",
---- 649=>x"3200", 650=>x"3100", 651=>x"3300", 652=>x"4b00",
---- 653=>x"3200", 654=>x"2f00", 655=>x"3900", 656=>x"4c00",
---- 657=>x"3100", 658=>x"2e00", 659=>x"3300", 660=>x"4800",
---- 661=>x"3800", 662=>x"3700", 663=>x"3500", 664=>x"4c00",
---- 665=>x"3400", 666=>x"4000", 667=>x"3600", 668=>x"4800",
---- 669=>x"3900", 670=>x"3f00", 671=>x"3900", 672=>x"4600",
---- 673=>x"3900", 674=>x"3e00", 675=>x"3100", 676=>x"4700",
---- 677=>x"3f00", 678=>x"3d00", 679=>x"2f00", 680=>x"3e00",
---- 681=>x"3d00", 682=>x"3a00", 683=>x"3400", 684=>x"3b00",
---- 685=>x"3c00", 686=>x"3c00", 687=>x"3200", 688=>x"4b00",
---- 689=>x"4100", 690=>x"4300", 691=>x"3400", 692=>x"4e00",
---- 693=>x"3d00", 694=>x"4400", 695=>x"3800", 696=>x"4800",
---- 697=>x"3800", 698=>x"3e00", 699=>x"3d00", 700=>x"4700",
---- 701=>x"2f00", 702=>x"3e00", 703=>x"4900", 704=>x"4500",
---- 705=>x"2c00", 706=>x"4000", 707=>x"5300", 708=>x"4c00",
---- 709=>x"3400", 710=>x"3f00", 711=>x"5800", 712=>x"3e00",
---- 713=>x"3300", 714=>x"4100", 715=>x"5500", 716=>x"4100",
---- 717=>x"3b00", 718=>x"4200", 719=>x"5500", 720=>x"4200",
---- 721=>x"4400", 722=>x"3c00", 723=>x"5300", 724=>x"4900",
---- 725=>x"4300", 726=>x"3600", 727=>x"5a00", 728=>x"4800",
---- 729=>x"3f00", 730=>x"3800", 731=>x"5400", 732=>x"4700",
---- 733=>x"3f00", 734=>x"3f00", 735=>x"5100", 736=>x"4500",
---- 737=>x"4000", 738=>x"3c00", 739=>x"5000", 740=>x"4b00",
---- 741=>x"4600", 742=>x"4500", 743=>x"5000", 744=>x"4b00",
---- 745=>x"4600", 746=>x"4a00", 747=>x"5300", 748=>x"4a00",
---- 749=>x"4100", 750=>x"4b00", 751=>x"5200", 752=>x"4800",
---- 753=>x"4600", 754=>x"4a00", 755=>x"4b00", 756=>x"4800",
---- 757=>x"4d00", 758=>x"af00", 759=>x"4c00", 760=>x"4400",
---- 761=>x"4e00", 762=>x"4f00", 763=>x"4b00", 764=>x"4b00",
---- 765=>x"ae00", 766=>x"5400", 767=>x"5200", 768=>x"4c00",
---- 769=>x"5400", 770=>x"5900", 771=>x"aa00", 772=>x"4d00",
---- 773=>x"5000", 774=>x"5500", 775=>x"5800", 776=>x"4e00",
---- 777=>x"af00", 778=>x"5700", 779=>x"5200", 780=>x"4e00",
---- 781=>x"4f00", 782=>x"5600", 783=>x"5a00", 784=>x"5400",
---- 785=>x"4c00", 786=>x"5000", 787=>x"5900", 788=>x"4f00",
---- 789=>x"4e00", 790=>x"5400", 791=>x"5900", 792=>x"4c00",
---- 793=>x"4900", 794=>x"5300", 795=>x"5700", 796=>x"4f00",
---- 797=>x"4c00", 798=>x"5000", 799=>x"5000", 800=>x"4e00",
---- 801=>x"4600", 802=>x"4d00", 803=>x"b400", 804=>x"4900",
---- 805=>x"4300", 806=>x"4b00", 807=>x"4a00", 808=>x"4800",
---- 809=>x"4900", 810=>x"5200", 811=>x"4a00", 812=>x"4200",
---- 813=>x"4200", 814=>x"4e00", 815=>x"4900", 816=>x"3b00",
---- 817=>x"4400", 818=>x"4e00", 819=>x"4500", 820=>x"3e00",
---- 821=>x"4d00", 822=>x"4f00", 823=>x"4700", 824=>x"3700",
---- 825=>x"4900", 826=>x"4700", 827=>x"4600", 828=>x"3600",
---- 829=>x"4900", 830=>x"3f00", 831=>x"4400", 832=>x"3400",
---- 833=>x"4400", 834=>x"3a00", 835=>x"3e00", 836=>x"3200",
---- 837=>x"3c00", 838=>x"3200", 839=>x"3b00", 840=>x"3000",
---- 841=>x"4200", 842=>x"2e00", 843=>x"3700", 844=>x"2c00",
---- 845=>x"3d00", 846=>x"2c00", 847=>x"3600", 848=>x"2700",
---- 849=>x"2f00", 850=>x"2c00", 851=>x"2e00", 852=>x"2100",
---- 853=>x"3100", 854=>x"2800", 855=>x"2a00", 856=>x"2a00",
---- 857=>x"2500", 858=>x"2300", 859=>x"2800", 860=>x"5400",
---- 861=>x"1f00", 862=>x"2700", 863=>x"2500", 864=>x"9000",
---- 865=>x"2700", 866=>x"2400", 867=>x"2400", 868=>x"be00",
---- 869=>x"3100", 870=>x"1800", 871=>x"2100", 872=>x"d800",
---- 873=>x"5a00", 874=>x"1800", 875=>x"df00", 876=>x"e000",
---- 877=>x"8b00", 878=>x"1900", 879=>x"1f00", 880=>x"e100",
---- 881=>x"b600", 882=>x"2800", 883=>x"1a00", 884=>x"de00",
---- 885=>x"d000", 886=>x"4b00", 887=>x"1500", 888=>x"d900",
---- 889=>x"dd00", 890=>x"7500", 891=>x"1600", 892=>x"d600",
---- 893=>x"df00", 894=>x"a000", 895=>x"1a00", 896=>x"d600",
---- 897=>x"dc00", 898=>x"c000", 899=>x"2d00", 900=>x"d700",
---- 901=>x"d900", 902=>x"d500", 903=>x"4f00", 904=>x"d600",
---- 905=>x"d500", 906=>x"dd00", 907=>x"8200", 908=>x"d500",
---- 909=>x"d500", 910=>x"dc00", 911=>x"ae00", 912=>x"d500",
---- 913=>x"d500", 914=>x"d800", 915=>x"c900", 916=>x"d500",
---- 917=>x"d500", 918=>x"d600", 919=>x"d900", 920=>x"d600",
---- 921=>x"d400", 922=>x"d600", 923=>x"dc00", 924=>x"d600",
---- 925=>x"d600", 926=>x"d700", 927=>x"dc00", 928=>x"d600",
---- 929=>x"d800", 930=>x"da00", 931=>x"db00", 932=>x"d500",
---- 933=>x"d700", 934=>x"d900", 935=>x"d900", 936=>x"d500",
---- 937=>x"d700", 938=>x"d900", 939=>x"d800", 940=>x"d400",
---- 941=>x"d500", 942=>x"d800", 943=>x"d900", 944=>x"d500",
---- 945=>x"d600", 946=>x"d900", 947=>x"d800", 948=>x"d500",
---- 949=>x"d500", 950=>x"d700", 951=>x"d800", 952=>x"d100",
---- 953=>x"d400", 954=>x"d600", 955=>x"d700", 956=>x"d100",
---- 957=>x"d400", 958=>x"d500", 959=>x"2800", 960=>x"d100",
---- 961=>x"d400", 962=>x"d600", 963=>x"d300", 964=>x"d300",
---- 965=>x"d400", 966=>x"d400", 967=>x"d300", 968=>x"d200",
---- 969=>x"d100", 970=>x"d500", 971=>x"d400", 972=>x"d200",
---- 973=>x"d300", 974=>x"d500", 975=>x"d400", 976=>x"d100",
---- 977=>x"d300", 978=>x"d500", 979=>x"d400", 980=>x"d100",
---- 981=>x"d000", 982=>x"d200", 983=>x"d200", 984=>x"cf00",
---- 985=>x"d000", 986=>x"d300", 987=>x"d400", 988=>x"cd00",
---- 989=>x"cf00", 990=>x"d300", 991=>x"d500", 992=>x"cc00",
---- 993=>x"cd00", 994=>x"d200", 995=>x"d400", 996=>x"ca00",
---- 997=>x"cb00", 998=>x"d100", 999=>x"d300", 1000=>x"ca00",
---- 1001=>x"cb00", 1002=>x"ce00", 1003=>x"d100", 1004=>x"c900",
---- 1005=>x"cb00", 1006=>x"cd00", 1007=>x"cd00", 1008=>x"c900",
---- 1009=>x"ca00", 1010=>x"cd00", 1011=>x"ce00", 1012=>x"c700",
---- 1013=>x"c900", 1014=>x"cb00", 1015=>x"ce00", 1016=>x"c500",
---- 1017=>x"c800", 1018=>x"ca00", 1019=>x"cc00", 1020=>x"c200",
---- 1021=>x"c500", 1022=>x"c800", 1023=>x"ca00"),
----
---- 46 => (0=>x"9a00", 1=>x"9800", 2=>x"9a00", 3=>x"9900", 4=>x"9a00",
---- 5=>x"9800", 6=>x"9a00", 7=>x"9900", 8=>x"9900",
---- 9=>x"9900", 10=>x"9900", 11=>x"9900", 12=>x"9900",
---- 13=>x"9800", 14=>x"9700", 15=>x"9a00", 16=>x"9c00",
---- 17=>x"9c00", 18=>x"6400", 19=>x"9800", 20=>x"9d00",
---- 21=>x"9d00", 22=>x"9a00", 23=>x"9b00", 24=>x"9d00",
---- 25=>x"9c00", 26=>x"9c00", 27=>x"9b00", 28=>x"9d00",
---- 29=>x"9c00", 30=>x"9c00", 31=>x"9b00", 32=>x"9e00",
---- 33=>x"9e00", 34=>x"9e00", 35=>x"9e00", 36=>x"9f00",
---- 37=>x"9e00", 38=>x"9e00", 39=>x"a000", 40=>x"a000",
---- 41=>x"9d00", 42=>x"9c00", 43=>x"9f00", 44=>x"a100",
---- 45=>x"a100", 46=>x"9c00", 47=>x"9a00", 48=>x"a100",
---- 49=>x"a100", 50=>x"9e00", 51=>x"9a00", 52=>x"9e00",
---- 53=>x"9f00", 54=>x"a000", 55=>x"9b00", 56=>x"9f00",
---- 57=>x"9f00", 58=>x"9e00", 59=>x"9c00", 60=>x"9e00",
---- 61=>x"9e00", 62=>x"9d00", 63=>x"9e00", 64=>x"9d00",
---- 65=>x"9e00", 66=>x"9e00", 67=>x"9a00", 68=>x"9f00",
---- 69=>x"9d00", 70=>x"9e00", 71=>x"9c00", 72=>x"9f00",
---- 73=>x"9b00", 74=>x"9b00", 75=>x"9a00", 76=>x"9d00",
---- 77=>x"9e00", 78=>x"9b00", 79=>x"9b00", 80=>x"9c00",
---- 81=>x"9b00", 82=>x"9b00", 83=>x"9b00", 84=>x"9900",
---- 85=>x"9b00", 86=>x"9b00", 87=>x"9a00", 88=>x"9a00",
---- 89=>x"9b00", 90=>x"9a00", 91=>x"9a00", 92=>x"9900",
---- 93=>x"9900", 94=>x"9900", 95=>x"9900", 96=>x"9800",
---- 97=>x"9700", 98=>x"9900", 99=>x"9a00", 100=>x"9800",
---- 101=>x"9900", 102=>x"9a00", 103=>x"9900", 104=>x"9900",
---- 105=>x"9900", 106=>x"9800", 107=>x"9700", 108=>x"9a00",
---- 109=>x"9800", 110=>x"9500", 111=>x"9600", 112=>x"9800",
---- 113=>x"9800", 114=>x"9600", 115=>x"9400", 116=>x"9600",
---- 117=>x"9a00", 118=>x"9600", 119=>x"9200", 120=>x"9700",
---- 121=>x"9800", 122=>x"9800", 123=>x"9500", 124=>x"9500",
---- 125=>x"9600", 126=>x"9900", 127=>x"9800", 128=>x"9300",
---- 129=>x"9400", 130=>x"9800", 131=>x"9800", 132=>x"9000",
---- 133=>x"9200", 134=>x"9600", 135=>x"9600", 136=>x"8d00",
---- 137=>x"8e00", 138=>x"9000", 139=>x"9500", 140=>x"7600",
---- 141=>x"8b00", 142=>x"8d00", 143=>x"9300", 144=>x"8200",
---- 145=>x"8500", 146=>x"8800", 147=>x"8d00", 148=>x"7c00",
---- 149=>x"7f00", 150=>x"8300", 151=>x"8a00", 152=>x"7400",
---- 153=>x"7800", 154=>x"8000", 155=>x"8700", 156=>x"6b00",
---- 157=>x"6e00", 158=>x"7500", 159=>x"7f00", 160=>x"5f00",
---- 161=>x"5f00", 162=>x"6900", 163=>x"7800", 164=>x"5500",
---- 165=>x"5400", 166=>x"5900", 167=>x"6900", 168=>x"4d00",
---- 169=>x"4400", 170=>x"4900", 171=>x"5e00", 172=>x"4100",
---- 173=>x"3700", 174=>x"3900", 175=>x"5300", 176=>x"4700",
---- 177=>x"3400", 178=>x"3200", 179=>x"4300", 180=>x"4c00",
---- 181=>x"3000", 182=>x"2a00", 183=>x"3500", 184=>x"4c00",
---- 185=>x"2f00", 186=>x"2900", 187=>x"2e00", 188=>x"4c00",
---- 189=>x"2f00", 190=>x"2400", 191=>x"2c00", 192=>x"4a00",
---- 193=>x"2e00", 194=>x"2b00", 195=>x"3100", 196=>x"4c00",
---- 197=>x"3100", 198=>x"2900", 199=>x"2e00", 200=>x"4f00",
---- 201=>x"3300", 202=>x"2d00", 203=>x"2a00", 204=>x"4e00",
---- 205=>x"3600", 206=>x"3100", 207=>x"2c00", 208=>x"5200",
---- 209=>x"3500", 210=>x"2d00", 211=>x"2a00", 212=>x"5300",
---- 213=>x"3800", 214=>x"2c00", 215=>x"2c00", 216=>x"5000",
---- 217=>x"3a00", 218=>x"2e00", 219=>x"2d00", 220=>x"5300",
---- 221=>x"3c00", 222=>x"3000", 223=>x"2d00", 224=>x"5200",
---- 225=>x"c200", 226=>x"3000", 227=>x"2c00", 228=>x"5100",
---- 229=>x"3900", 230=>x"2f00", 231=>x"2b00", 232=>x"5500",
---- 233=>x"3900", 234=>x"2e00", 235=>x"2d00", 236=>x"5100",
---- 237=>x"3900", 238=>x"2c00", 239=>x"2900", 240=>x"5100",
---- 241=>x"3500", 242=>x"2c00", 243=>x"2800", 244=>x"4a00",
---- 245=>x"2e00", 246=>x"2800", 247=>x"2500", 248=>x"4200",
---- 249=>x"2900", 250=>x"db00", 251=>x"2200", 252=>x"3f00",
---- 253=>x"2700", 254=>x"1e00", 255=>x"d300", 256=>x"3200",
---- 257=>x"2500", 258=>x"4500", 259=>x"9300", 260=>x"3d00",
---- 261=>x"7300", 262=>x"ba00", 263=>x"dc00", 264=>x"9e00",
---- 265=>x"d700", 266=>x"d700", 267=>x"c800", 268=>x"de00",
---- 269=>x"cf00", 270=>x"be00", 271=>x"b900", 272=>x"c500",
---- 273=>x"bc00", 274=>x"b800", 275=>x"bc00", 276=>x"bd00",
---- 277=>x"b600", 278=>x"be00", 279=>x"cc00", 280=>x"b900",
---- 281=>x"c800", 282=>x"d400", 283=>x"d300", 284=>x"cd00",
---- 285=>x"d500", 286=>x"d100", 287=>x"ce00", 288=>x"d300",
---- 289=>x"d000", 290=>x"cc00", 291=>x"cc00", 292=>x"cd00",
---- 293=>x"cc00", 294=>x"ca00", 295=>x"c900", 296=>x"c900",
---- 297=>x"ca00", 298=>x"c900", 299=>x"c800", 300=>x"c800",
---- 301=>x"c800", 302=>x"c800", 303=>x"c900", 304=>x"c800",
---- 305=>x"c900", 306=>x"c700", 307=>x"c700", 308=>x"c800",
---- 309=>x"c800", 310=>x"c600", 311=>x"c700", 312=>x"c800",
---- 313=>x"c700", 314=>x"c600", 315=>x"c900", 316=>x"c700",
---- 317=>x"c900", 318=>x"c500", 319=>x"c900", 320=>x"c900",
---- 321=>x"ca00", 322=>x"c800", 323=>x"cb00", 324=>x"c800",
---- 325=>x"c700", 326=>x"ca00", 327=>x"ca00", 328=>x"c800",
---- 329=>x"cb00", 330=>x"cb00", 331=>x"cb00", 332=>x"ca00",
---- 333=>x"ca00", 334=>x"cb00", 335=>x"cc00", 336=>x"c900",
---- 337=>x"cb00", 338=>x"3400", 339=>x"ce00", 340=>x"ca00",
---- 341=>x"cd00", 342=>x"cc00", 343=>x"d000", 344=>x"c900",
---- 345=>x"ce00", 346=>x"cd00", 347=>x"d100", 348=>x"cc00",
---- 349=>x"cf00", 350=>x"d000", 351=>x"d200", 352=>x"cc00",
---- 353=>x"ce00", 354=>x"d300", 355=>x"d500", 356=>x"ce00",
---- 357=>x"d300", 358=>x"ce00", 359=>x"b800", 360=>x"ca00",
---- 361=>x"ad00", 362=>x"8800", 363=>x"6e00", 364=>x"7700",
---- 365=>x"5d00", 366=>x"5500", 367=>x"5500", 368=>x"5300",
---- 369=>x"5600", 370=>x"5600", 371=>x"5900", 372=>x"5c00",
---- 373=>x"5a00", 374=>x"5600", 375=>x"5900", 376=>x"5900",
---- 377=>x"5700", 378=>x"5800", 379=>x"5f00", 380=>x"5b00",
---- 381=>x"6900", 382=>x"7500", 383=>x"8700", 384=>x"8800",
---- 385=>x"9b00", 386=>x"a300", 387=>x"a800", 388=>x"a700",
---- 389=>x"a700", 390=>x"a700", 391=>x"a600", 392=>x"a600",
---- 393=>x"a700", 394=>x"a600", 395=>x"a600", 396=>x"aa00",
---- 397=>x"aa00", 398=>x"aa00", 399=>x"ac00", 400=>x"ab00",
---- 401=>x"ac00", 402=>x"b000", 403=>x"b100", 404=>x"a700",
---- 405=>x"ac00", 406=>x"ae00", 407=>x"be00", 408=>x"ae00",
---- 409=>x"b500", 410=>x"c300", 411=>x"ce00", 412=>x"c000",
---- 413=>x"ce00", 414=>x"4900", 415=>x"7100", 416=>x"bd00",
---- 417=>x"9100", 418=>x"4b00", 419=>x"2a00", 420=>x"8300",
---- 421=>x"5000", 422=>x"2800", 423=>x"2c00", 424=>x"7400",
---- 425=>x"5800", 426=>x"2b00", 427=>x"2500", 428=>x"7600",
---- 429=>x"4a00", 430=>x"2f00", 431=>x"2900", 432=>x"7600",
---- 433=>x"3e00", 434=>x"2c00", 435=>x"2b00", 436=>x"6400",
---- 437=>x"3500", 438=>x"3400", 439=>x"3000", 440=>x"5500",
---- 441=>x"2e00", 442=>x"3200", 443=>x"2f00", 444=>x"4d00",
---- 445=>x"2a00", 446=>x"3000", 447=>x"2b00", 448=>x"4e00",
---- 449=>x"2d00", 450=>x"3400", 451=>x"2f00", 452=>x"5f00",
---- 453=>x"3400", 454=>x"3c00", 455=>x"3000", 456=>x"6a00",
---- 457=>x"3500", 458=>x"3200", 459=>x"3900", 460=>x"6600",
---- 461=>x"3e00", 462=>x"3300", 463=>x"3800", 464=>x"6d00",
---- 465=>x"b300", 466=>x"2e00", 467=>x"2f00", 468=>x"7400",
---- 469=>x"4600", 470=>x"2900", 471=>x"3200", 472=>x"7500",
---- 473=>x"bf00", 474=>x"3b00", 475=>x"3000", 476=>x"8400",
---- 477=>x"4600", 478=>x"3500", 479=>x"3100", 480=>x"8f00",
---- 481=>x"4f00", 482=>x"3500", 483=>x"3800", 484=>x"9600",
---- 485=>x"5100", 486=>x"4400", 487=>x"3b00", 488=>x"9e00",
---- 489=>x"5a00", 490=>x"3f00", 491=>x"3a00", 492=>x"a300",
---- 493=>x"6e00", 494=>x"3800", 495=>x"3600", 496=>x"ac00",
---- 497=>x"7c00", 498=>x"3d00", 499=>x"3000", 500=>x"a900",
---- 501=>x"8400", 502=>x"4800", 503=>x"3500", 504=>x"a800",
---- 505=>x"8400", 506=>x"5400", 507=>x"3400", 508=>x"ad00",
---- 509=>x"8000", 510=>x"5f00", 511=>x"3600", 512=>x"b100",
---- 513=>x"7900", 514=>x"6a00", 515=>x"3b00", 516=>x"b300",
---- 517=>x"8200", 518=>x"6700", 519=>x"4c00", 520=>x"b400",
---- 521=>x"8200", 522=>x"6100", 523=>x"4e00", 524=>x"b800",
---- 525=>x"8900", 526=>x"5a00", 527=>x"4b00", 528=>x"b700",
---- 529=>x"8900", 530=>x"5c00", 531=>x"5800", 532=>x"b600",
---- 533=>x"8f00", 534=>x"5b00", 535=>x"5d00", 536=>x"b800",
---- 537=>x"9c00", 538=>x"5600", 539=>x"5d00", 540=>x"b700",
---- 541=>x"a000", 542=>x"5900", 543=>x"5200", 544=>x"b300",
---- 545=>x"a500", 546=>x"5e00", 547=>x"4c00", 548=>x"b100",
---- 549=>x"ad00", 550=>x"6a00", 551=>x"4f00", 552=>x"a700",
---- 553=>x"b100", 554=>x"7700", 555=>x"4d00", 556=>x"a700",
---- 557=>x"b400", 558=>x"8500", 559=>x"4f00", 560=>x"a100",
---- 561=>x"b700", 562=>x"6d00", 563=>x"5600", 564=>x"a000",
---- 565=>x"b400", 566=>x"9300", 567=>x"5b00", 568=>x"a000",
---- 569=>x"b500", 570=>x"9500", 571=>x"6000", 572=>x"9e00",
---- 573=>x"b300", 574=>x"a100", 575=>x"6100", 576=>x"9c00",
---- 577=>x"b400", 578=>x"aa00", 579=>x"6700", 580=>x"9a00",
---- 581=>x"ad00", 582=>x"a800", 583=>x"9100", 584=>x"9300",
---- 585=>x"af00", 586=>x"a500", 587=>x"8100", 588=>x"8e00",
---- 589=>x"ac00", 590=>x"9d00", 591=>x"9400", 592=>x"8800",
---- 593=>x"ac00", 594=>x"8d00", 595=>x"9b00", 596=>x"8000",
---- 597=>x"ad00", 598=>x"8a00", 599=>x"a200", 600=>x"7f00",
---- 601=>x"b300", 602=>x"9100", 603=>x"a100", 604=>x"7300",
---- 605=>x"4800", 606=>x"9400", 607=>x"9800", 608=>x"6a00",
---- 609=>x"ad00", 610=>x"9600", 611=>x"9100", 612=>x"6000",
---- 613=>x"a700", 614=>x"9400", 615=>x"8e00", 616=>x"5700",
---- 617=>x"a300", 618=>x"9a00", 619=>x"9100", 620=>x"4e00",
---- 621=>x"9900", 622=>x"a300", 623=>x"9100", 624=>x"4900",
---- 625=>x"9200", 626=>x"a400", 627=>x"8e00", 628=>x"4000",
---- 629=>x"8300", 630=>x"a400", 631=>x"9000", 632=>x"3200",
---- 633=>x"7a00", 634=>x"a700", 635=>x"9800", 636=>x"2d00",
---- 637=>x"6e00", 638=>x"a800", 639=>x"9d00", 640=>x"2900",
---- 641=>x"6000", 642=>x"a500", 643=>x"a400", 644=>x"2300",
---- 645=>x"5500", 646=>x"a200", 647=>x"a800", 648=>x"2100",
---- 649=>x"4600", 650=>x"9a00", 651=>x"ab00", 652=>x"2100",
---- 653=>x"3700", 654=>x"9100", 655=>x"ac00", 656=>x"dc00",
---- 657=>x"2d00", 658=>x"8800", 659=>x"af00", 660=>x"2900",
---- 661=>x"2800", 662=>x"7a00", 663=>x"ae00", 664=>x"2900",
---- 665=>x"2300", 666=>x"6900", 667=>x"ac00", 668=>x"3000",
---- 669=>x"2400", 670=>x"5900", 671=>x"a800", 672=>x"2b00",
---- 673=>x"2300", 674=>x"4a00", 675=>x"9d00", 676=>x"2800",
---- 677=>x"2300", 678=>x"4300", 679=>x"9500", 680=>x"2c00",
---- 681=>x"2600", 682=>x"4500", 683=>x"8e00", 684=>x"2b00",
---- 685=>x"2300", 686=>x"c100", 687=>x"8800", 688=>x"2800",
---- 689=>x"2300", 690=>x"3300", 691=>x"8000", 692=>x"2700",
---- 693=>x"2700", 694=>x"2d00", 695=>x"7800", 696=>x"2600",
---- 697=>x"2700", 698=>x"2a00", 699=>x"6c00", 700=>x"2e00",
---- 701=>x"2800", 702=>x"2a00", 703=>x"5e00", 704=>x"2f00",
---- 705=>x"2a00", 706=>x"2c00", 707=>x"5300", 708=>x"3100",
---- 709=>x"2d00", 710=>x"2b00", 711=>x"4b00", 712=>x"3600",
---- 713=>x"2800", 714=>x"2d00", 715=>x"4a00", 716=>x"3e00",
---- 717=>x"d300", 718=>x"2e00", 719=>x"4900", 720=>x"3e00",
---- 721=>x"2f00", 722=>x"3000", 723=>x"4800", 724=>x"4300",
---- 725=>x"3000", 726=>x"2f00", 727=>x"4300", 728=>x"4400",
---- 729=>x"2e00", 730=>x"2f00", 731=>x"4000", 732=>x"4300",
---- 733=>x"3700", 734=>x"3700", 735=>x"3f00", 736=>x"4d00",
---- 737=>x"3100", 738=>x"3200", 739=>x"3700", 740=>x"4a00",
---- 741=>x"3100", 742=>x"3800", 743=>x"3500", 744=>x"4800",
---- 745=>x"3800", 746=>x"3900", 747=>x"3600", 748=>x"4000",
---- 749=>x"4500", 750=>x"3800", 751=>x"3500", 752=>x"3d00",
---- 753=>x"4e00", 754=>x"3300", 755=>x"3000", 756=>x"3e00",
---- 757=>x"4f00", 758=>x"3d00", 759=>x"3000", 760=>x"3f00",
---- 761=>x"5100", 762=>x"3c00", 763=>x"3000", 764=>x"4400",
---- 765=>x"5600", 766=>x"3c00", 767=>x"3000", 768=>x"4400",
---- 769=>x"5400", 770=>x"3f00", 771=>x"3600", 772=>x"4200",
---- 773=>x"4e00", 774=>x"4600", 775=>x"3a00", 776=>x"4100",
---- 777=>x"4b00", 778=>x"4600", 779=>x"4100", 780=>x"4600",
---- 781=>x"4c00", 782=>x"4400", 783=>x"4500", 784=>x"4b00",
---- 785=>x"4e00", 786=>x"4200", 787=>x"4600", 788=>x"4900",
---- 789=>x"5200", 790=>x"4a00", 791=>x"b200", 792=>x"4400",
---- 793=>x"4e00", 794=>x"4500", 795=>x"5000", 796=>x"4500",
---- 797=>x"4600", 798=>x"3c00", 799=>x"5700", 800=>x"4700",
---- 801=>x"4b00", 802=>x"3e00", 803=>x"a200", 804=>x"4b00",
---- 805=>x"4700", 806=>x"3900", 807=>x"6500", 808=>x"4600",
---- 809=>x"4000", 810=>x"3700", 811=>x"7500", 812=>x"4600",
---- 813=>x"3900", 814=>x"3600", 815=>x"7c00", 816=>x"ba00",
---- 817=>x"3200", 818=>x"3100", 819=>x"8100", 820=>x"4300",
---- 821=>x"3300", 822=>x"3800", 823=>x"8d00", 824=>x"4d00",
---- 825=>x"2f00", 826=>x"3c00", 827=>x"6600", 828=>x"4600",
---- 829=>x"2c00", 830=>x"4500", 831=>x"9d00", 832=>x"c500",
---- 833=>x"2400", 834=>x"4d00", 835=>x"a500", 836=>x"3b00",
---- 837=>x"2400", 838=>x"5b00", 839=>x"a400", 840=>x"3800",
---- 841=>x"2300", 842=>x"6900", 843=>x"a200", 844=>x"2d00",
---- 845=>x"2200", 846=>x"7000", 847=>x"9e00", 848=>x"2500",
---- 849=>x"2a00", 850=>x"7d00", 851=>x"a100", 852=>x"2200",
---- 853=>x"2d00", 854=>x"8600", 855=>x"9d00", 856=>x"1e00",
---- 857=>x"3400", 858=>x"8b00", 859=>x"9c00", 860=>x"1f00",
---- 861=>x"3f00", 862=>x"8e00", 863=>x"9600", 864=>x"1b00",
---- 865=>x"4900", 866=>x"9600", 867=>x"8d00", 868=>x"1b00",
---- 869=>x"5900", 870=>x"9300", 871=>x"8e00", 872=>x"1d00",
---- 873=>x"6300", 874=>x"8f00", 875=>x"8e00", 876=>x"2300",
---- 877=>x"6e00", 878=>x"8c00", 879=>x"8d00", 880=>x"2500",
---- 881=>x"7400", 882=>x"8b00", 883=>x"8b00", 884=>x"2b00",
---- 885=>x"7700", 886=>x"8c00", 887=>x"8c00", 888=>x"3300",
---- 889=>x"7d00", 890=>x"8a00", 891=>x"8e00", 892=>x"3b00",
---- 893=>x"8500", 894=>x"8b00", 895=>x"8f00", 896=>x"3e00",
---- 897=>x"8400", 898=>x"8b00", 899=>x"8e00", 900=>x"3f00",
---- 901=>x"8500", 902=>x"8d00", 903=>x"9200", 904=>x"4700",
---- 905=>x"8500", 906=>x"8f00", 907=>x"8f00", 908=>x"5f00",
---- 909=>x"8700", 910=>x"9000", 911=>x"8c00", 912=>x"7b00",
---- 913=>x"8600", 914=>x"9300", 915=>x"8300", 916=>x"9a00",
---- 917=>x"8800", 918=>x"8f00", 919=>x"7100", 920=>x"b600",
---- 921=>x"8700", 922=>x"7900", 923=>x"6100", 924=>x"cd00",
---- 925=>x"7800", 926=>x"5b00", 927=>x"4f00", 928=>x"da00",
---- 929=>x"8900", 930=>x"4800", 931=>x"4f00", 932=>x"df00",
---- 933=>x"9f00", 934=>x"4800", 935=>x"5500", 936=>x"df00",
---- 937=>x"b900", 938=>x"5000", 939=>x"5000", 940=>x"db00",
---- 941=>x"d200", 942=>x"6200", 943=>x"4900", 944=>x"d800",
---- 945=>x"dc00", 946=>x"8a00", 947=>x"4a00", 948=>x"d700",
---- 949=>x"dd00", 950=>x"ae00", 951=>x"5100", 952=>x"d700",
---- 953=>x"dc00", 954=>x"c700", 955=>x"6400", 956=>x"d700",
---- 957=>x"d900", 958=>x"d900", 959=>x"7c00", 960=>x"d500",
---- 961=>x"d700", 962=>x"dc00", 963=>x"9c00", 964=>x"d400",
---- 965=>x"d800", 966=>x"db00", 967=>x"bc00", 968=>x"d400",
---- 969=>x"d800", 970=>x"d800", 971=>x"d200", 972=>x"d500",
---- 973=>x"d800", 974=>x"d700", 975=>x"d900", 976=>x"2a00",
---- 977=>x"d700", 978=>x"d600", 979=>x"da00", 980=>x"d300",
---- 981=>x"d700", 982=>x"d500", 983=>x"d700", 984=>x"d400",
---- 985=>x"d700", 986=>x"d700", 987=>x"d600", 988=>x"d400",
---- 989=>x"d400", 990=>x"d600", 991=>x"d600", 992=>x"d300",
---- 993=>x"d400", 994=>x"d500", 995=>x"d500", 996=>x"d200",
---- 997=>x"d200", 998=>x"d400", 999=>x"d500", 1000=>x"d200",
---- 1001=>x"d000", 1002=>x"d100", 1003=>x"d300", 1004=>x"d000",
---- 1005=>x"d100", 1006=>x"d100", 1007=>x"d200", 1008=>x"cf00",
---- 1009=>x"d200", 1010=>x"d300", 1011=>x"d300", 1012=>x"cd00",
---- 1013=>x"d000", 1014=>x"d300", 1015=>x"d300", 1016=>x"cd00",
---- 1017=>x"d000", 1018=>x"d200", 1019=>x"d000", 1020=>x"cc00",
---- 1021=>x"cf00", 1022=>x"d100", 1023=>x"d100"),
----
---- 47 => (0=>x"9800", 1=>x"9900", 2=>x"9c00", 3=>x"9900", 4=>x"9800",
---- 5=>x"9900", 6=>x"9c00", 7=>x"9800", 8=>x"9800",
---- 9=>x"9900", 10=>x"9d00", 11=>x"9a00", 12=>x"9c00",
---- 13=>x"9a00", 14=>x"9b00", 15=>x"9800", 16=>x"9a00",
---- 17=>x"9900", 18=>x"9900", 19=>x"9900", 20=>x"9a00",
---- 21=>x"9d00", 22=>x"9b00", 23=>x"6600", 24=>x"9c00",
---- 25=>x"9c00", 26=>x"9b00", 27=>x"9900", 28=>x"9d00",
---- 29=>x"9b00", 30=>x"9800", 31=>x"9a00", 32=>x"9d00",
---- 33=>x"9a00", 34=>x"9900", 35=>x"9a00", 36=>x"9f00",
---- 37=>x"9d00", 38=>x"9b00", 39=>x"9a00", 40=>x"9e00",
---- 41=>x"9f00", 42=>x"9a00", 43=>x"9c00", 44=>x"9d00",
---- 45=>x"9b00", 46=>x"9b00", 47=>x"9b00", 48=>x"9b00",
---- 49=>x"9d00", 50=>x"9c00", 51=>x"9b00", 52=>x"9c00",
---- 53=>x"9e00", 54=>x"9b00", 55=>x"9b00", 56=>x"9d00",
---- 57=>x"9b00", 58=>x"9c00", 59=>x"9e00", 60=>x"9e00",
---- 61=>x"9b00", 62=>x"9a00", 63=>x"9c00", 64=>x"9d00",
---- 65=>x"9b00", 66=>x"9d00", 67=>x"9c00", 68=>x"9d00",
---- 69=>x"9d00", 70=>x"9c00", 71=>x"9c00", 72=>x"a000",
---- 73=>x"9e00", 74=>x"9a00", 75=>x"9f00", 76=>x"9d00",
---- 77=>x"9d00", 78=>x"9900", 79=>x"9900", 80=>x"9b00",
---- 81=>x"9a00", 82=>x"9800", 83=>x"9800", 84=>x"9b00",
---- 85=>x"9900", 86=>x"9900", 87=>x"9a00", 88=>x"9b00",
---- 89=>x"9900", 90=>x"9b00", 91=>x"9c00", 92=>x"9a00",
---- 93=>x"9a00", 94=>x"9b00", 95=>x"9a00", 96=>x"6600",
---- 97=>x"6600", 98=>x"9c00", 99=>x"9a00", 100=>x"9900",
---- 101=>x"9900", 102=>x"9a00", 103=>x"9900", 104=>x"9a00",
---- 105=>x"9800", 106=>x"9700", 107=>x"9800", 108=>x"9800",
---- 109=>x"9700", 110=>x"9400", 111=>x"9200", 112=>x"9600",
---- 113=>x"9600", 114=>x"9300", 115=>x"9300", 116=>x"6c00",
---- 117=>x"9200", 118=>x"9400", 119=>x"9300", 120=>x"9300",
---- 121=>x"8e00", 122=>x"9200", 123=>x"9100", 124=>x"9500",
---- 125=>x"9200", 126=>x"9000", 127=>x"8d00", 128=>x"9500",
---- 129=>x"9200", 130=>x"8e00", 131=>x"8e00", 132=>x"9700",
---- 133=>x"9000", 134=>x"8e00", 135=>x"8b00", 136=>x"9900",
---- 137=>x"9200", 138=>x"8f00", 139=>x"8f00", 140=>x"9600",
---- 141=>x"9400", 142=>x"9100", 143=>x"9100", 144=>x"9500",
---- 145=>x"9600", 146=>x"9300", 147=>x"6e00", 148=>x"9200",
---- 149=>x"9700", 150=>x"9500", 151=>x"9100", 152=>x"8e00",
---- 153=>x"9300", 154=>x"9600", 155=>x"6c00", 156=>x"8b00",
---- 157=>x"8f00", 158=>x"9400", 159=>x"9500", 160=>x"8300",
---- 161=>x"8a00", 162=>x"9200", 163=>x"9700", 164=>x"7b00",
---- 165=>x"8800", 166=>x"8e00", 167=>x"9300", 168=>x"7300",
---- 169=>x"8200", 170=>x"8800", 171=>x"9000", 172=>x"6b00",
---- 173=>x"7b00", 174=>x"8500", 175=>x"8a00", 176=>x"a500",
---- 177=>x"7100", 178=>x"7d00", 179=>x"8800", 180=>x"4e00",
---- 181=>x"6600", 182=>x"7300", 183=>x"7f00", 184=>x"4500",
---- 185=>x"6000", 186=>x"6b00", 187=>x"7800", 188=>x"3b00",
---- 189=>x"5600", 190=>x"6800", 191=>x"7400", 192=>x"3400",
---- 193=>x"4d00", 194=>x"6100", 195=>x"6b00", 196=>x"3700",
---- 197=>x"3400", 198=>x"4e00", 199=>x"6100", 200=>x"2700",
---- 201=>x"2d00", 202=>x"3b00", 203=>x"5200", 204=>x"2500",
---- 205=>x"2d00", 206=>x"3100", 207=>x"4600", 208=>x"2800",
---- 209=>x"2900", 210=>x"2b00", 211=>x"3600", 212=>x"2f00",
---- 213=>x"2900", 214=>x"2900", 215=>x"2c00", 216=>x"2d00",
---- 217=>x"2b00", 218=>x"2800", 219=>x"2700", 220=>x"2e00",
---- 221=>x"2d00", 222=>x"2900", 223=>x"2800", 224=>x"2c00",
---- 225=>x"2e00", 226=>x"2b00", 227=>x"2a00", 228=>x"2f00",
---- 229=>x"2c00", 230=>x"2c00", 231=>x"2700", 232=>x"2e00",
---- 233=>x"2b00", 234=>x"2700", 235=>x"2600", 236=>x"2a00",
---- 237=>x"2600", 238=>x"2600", 239=>x"2400", 240=>x"2800",
---- 241=>x"2700", 242=>x"2100", 243=>x"3300", 244=>x"2400",
---- 245=>x"2200", 246=>x"4600", 247=>x"a200", 248=>x"2300",
---- 249=>x"5c00", 250=>x"b700", 251=>x"d900", 252=>x"7300",
---- 253=>x"c800", 254=>x"de00", 255=>x"d100", 256=>x"d500",
---- 257=>x"db00", 258=>x"ce00", 259=>x"a900", 260=>x"d200",
---- 261=>x"c000", 262=>x"ac00", 263=>x"b600", 264=>x"b900",
---- 265=>x"ad00", 266=>x"bc00", 267=>x"d400", 268=>x"b900",
---- 269=>x"c400", 270=>x"d300", 271=>x"d500", 272=>x"c900",
---- 273=>x"d300", 274=>x"d500", 275=>x"d200", 276=>x"d400",
---- 277=>x"d300", 278=>x"d000", 279=>x"cf00", 280=>x"d100",
---- 281=>x"ce00", 282=>x"cb00", 283=>x"ca00", 284=>x"cc00",
---- 285=>x"c800", 286=>x"c700", 287=>x"c900", 288=>x"c800",
---- 289=>x"c800", 290=>x"c900", 291=>x"c900", 292=>x"c900",
---- 293=>x"c700", 294=>x"c500", 295=>x"c800", 296=>x"ca00",
---- 297=>x"c600", 298=>x"c600", 299=>x"c900", 300=>x"c600",
---- 301=>x"c600", 302=>x"3800", 303=>x"ca00", 304=>x"c500",
---- 305=>x"c600", 306=>x"c900", 307=>x"cc00", 308=>x"c900",
---- 309=>x"c900", 310=>x"cb00", 311=>x"cc00", 312=>x"ca00",
---- 313=>x"c900", 314=>x"cb00", 315=>x"3200", 316=>x"ca00",
---- 317=>x"ca00", 318=>x"cc00", 319=>x"cc00", 320=>x"c700",
---- 321=>x"cd00", 322=>x"cf00", 323=>x"ce00", 324=>x"ca00",
---- 325=>x"3100", 326=>x"d000", 327=>x"cf00", 328=>x"cd00",
---- 329=>x"ce00", 330=>x"d100", 331=>x"d200", 332=>x"d000",
---- 333=>x"d200", 334=>x"d100", 335=>x"d300", 336=>x"d100",
---- 337=>x"d100", 338=>x"d500", 339=>x"ca00", 340=>x"d300",
---- 341=>x"d100", 342=>x"d600", 343=>x"ac00", 344=>x"d300",
---- 345=>x"d600", 346=>x"c200", 347=>x"9b00", 348=>x"d900",
---- 349=>x"cb00", 350=>x"a900", 351=>x"a600", 352=>x"c900",
---- 353=>x"af00", 354=>x"9700", 355=>x"8400", 356=>x"9a00",
---- 357=>x"7e00", 358=>x"6500", 359=>x"5000", 360=>x"6200",
---- 361=>x"5b00", 362=>x"5600", 363=>x"5500", 364=>x"5b00",
---- 365=>x"5d00", 366=>x"5b00", 367=>x"5800", 368=>x"9f00",
---- 369=>x"5a00", 370=>x"5c00", 371=>x"6000", 372=>x"6000",
---- 373=>x"6600", 374=>x"6e00", 375=>x"7900", 376=>x"7200",
---- 377=>x"8300", 378=>x"9500", 379=>x"9d00", 380=>x"9b00",
---- 381=>x"9f00", 382=>x"a800", 383=>x"aa00", 384=>x"a900",
---- 385=>x"a500", 386=>x"a500", 387=>x"ad00", 388=>x"aa00",
---- 389=>x"a800", 390=>x"a800", 391=>x"b200", 392=>x"a900",
---- 393=>x"b000", 394=>x"b700", 395=>x"c900", 396=>x"b200",
---- 397=>x"b900", 398=>x"c900", 399=>x"d500", 400=>x"b900",
---- 401=>x"ce00", 402=>x"b600", 403=>x"6900", 404=>x"d000",
---- 405=>x"a300", 406=>x"3f00", 407=>x"2100", 408=>x"8a00",
---- 409=>x"3300", 410=>x"2500", 411=>x"2f00", 412=>x"2e00",
---- 413=>x"2a00", 414=>x"2a00", 415=>x"2c00", 416=>x"2b00",
---- 417=>x"2f00", 418=>x"2d00", 419=>x"2d00", 420=>x"2900",
---- 421=>x"2e00", 422=>x"2c00", 423=>x"3100", 424=>x"2c00",
---- 425=>x"2e00", 426=>x"2a00", 427=>x"2c00", 428=>x"2900",
---- 429=>x"2600", 430=>x"2c00", 431=>x"2e00", 432=>x"2a00",
---- 433=>x"2a00", 434=>x"2f00", 435=>x"2e00", 436=>x"3000",
---- 437=>x"3000", 438=>x"2e00", 439=>x"2f00", 440=>x"2c00",
---- 441=>x"2d00", 442=>x"2f00", 443=>x"3100", 444=>x"2d00",
---- 445=>x"3000", 446=>x"2e00", 447=>x"3300", 448=>x"3400",
---- 449=>x"3800", 450=>x"3600", 451=>x"3700", 452=>x"3100",
---- 453=>x"3200", 454=>x"3400", 455=>x"3800", 456=>x"3000",
---- 457=>x"3300", 458=>x"3300", 459=>x"3700", 460=>x"3500",
---- 461=>x"3900", 462=>x"3500", 463=>x"3700", 464=>x"3000",
---- 465=>x"3900", 466=>x"3a00", 467=>x"3600", 468=>x"3400",
---- 469=>x"3800", 470=>x"3700", 471=>x"3b00", 472=>x"3000",
---- 473=>x"3a00", 474=>x"3800", 475=>x"3b00", 476=>x"2f00",
---- 477=>x"3900", 478=>x"3700", 479=>x"3800", 480=>x"3a00",
---- 481=>x"4100", 482=>x"3a00", 483=>x"3c00", 484=>x"3d00",
---- 485=>x"4900", 486=>x"3b00", 487=>x"3800", 488=>x"3d00",
---- 489=>x"3c00", 490=>x"3f00", 491=>x"3c00", 492=>x"4500",
---- 493=>x"3f00", 494=>x"3700", 495=>x"3b00", 496=>x"3d00",
---- 497=>x"4500", 498=>x"3e00", 499=>x"3d00", 500=>x"3600",
---- 501=>x"4400", 502=>x"4600", 503=>x"4300", 504=>x"3400",
---- 505=>x"b900", 506=>x"3f00", 507=>x"3c00", 508=>x"2e00",
---- 509=>x"3e00", 510=>x"3e00", 511=>x"3e00", 512=>x"2c00",
---- 513=>x"4300", 514=>x"4500", 515=>x"4000", 516=>x"3100",
---- 517=>x"c200", 518=>x"4700", 519=>x"3c00", 520=>x"3c00",
---- 521=>x"3a00", 522=>x"4400", 523=>x"3a00", 524=>x"3900",
---- 525=>x"4300", 526=>x"4b00", 527=>x"3c00", 528=>x"3d00",
---- 529=>x"4700", 530=>x"4a00", 531=>x"3c00", 532=>x"4400",
---- 533=>x"4c00", 534=>x"4400", 535=>x"3b00", 536=>x"4c00",
---- 537=>x"5300", 538=>x"4100", 539=>x"3c00", 540=>x"ad00",
---- 541=>x"5300", 542=>x"3f00", 543=>x"3700", 544=>x"5900",
---- 545=>x"5700", 546=>x"4200", 547=>x"3100", 548=>x"5f00",
---- 549=>x"4d00", 550=>x"3d00", 551=>x"3700", 552=>x"5c00",
---- 553=>x"4c00", 554=>x"3d00", 555=>x"3700", 556=>x"5600",
---- 557=>x"5300", 558=>x"3500", 559=>x"3000", 560=>x"4f00",
---- 561=>x"4f00", 562=>x"3200", 563=>x"3500", 564=>x"4200",
---- 565=>x"4c00", 566=>x"3300", 567=>x"3200", 568=>x"4500",
---- 569=>x"4e00", 570=>x"3000", 571=>x"3400", 572=>x"4000",
---- 573=>x"4b00", 574=>x"2b00", 575=>x"3700", 576=>x"3b00",
---- 577=>x"4400", 578=>x"2600", 579=>x"3700", 580=>x"3900",
---- 581=>x"3a00", 582=>x"2400", 583=>x"3c00", 584=>x"3c00",
---- 585=>x"3900", 586=>x"2600", 587=>x"3700", 588=>x"4200",
---- 589=>x"3100", 590=>x"2900", 591=>x"2d00", 592=>x"4d00",
---- 593=>x"2800", 594=>x"2400", 595=>x"2b00", 596=>x"5d00",
---- 597=>x"2400", 598=>x"2a00", 599=>x"2d00", 600=>x"6d00",
---- 601=>x"2500", 602=>x"2800", 603=>x"2b00", 604=>x"8200",
---- 605=>x"3000", 606=>x"2700", 607=>x"2500", 608=>x"8400",
---- 609=>x"4300", 610=>x"2b00", 611=>x"2a00", 612=>x"8900",
---- 613=>x"4c00", 614=>x"2300", 615=>x"2d00", 616=>x"9300",
---- 617=>x"5200", 618=>x"1b00", 619=>x"2b00", 620=>x"9700",
---- 621=>x"5600", 622=>x"1c00", 623=>x"3000", 624=>x"9900",
---- 625=>x"6000", 626=>x"2400", 627=>x"2f00", 628=>x"9a00",
---- 629=>x"7300", 630=>x"3300", 631=>x"2b00", 632=>x"9c00",
---- 633=>x"8200", 634=>x"3c00", 635=>x"2d00", 636=>x"9600",
---- 637=>x"8500", 638=>x"4600", 639=>x"2c00", 640=>x"9400",
---- 641=>x"8200", 642=>x"5000", 643=>x"2a00", 644=>x"8f00",
---- 645=>x"8900", 646=>x"5700", 647=>x"2800", 648=>x"8500",
---- 649=>x"8d00", 650=>x"5f00", 651=>x"2700", 652=>x"8a00",
---- 653=>x"8f00", 654=>x"6a00", 655=>x"2b00", 656=>x"8b00",
---- 657=>x"8d00", 658=>x"7100", 659=>x"3600", 660=>x"8b00",
---- 661=>x"8600", 662=>x"6c00", 663=>x"3f00", 664=>x"9000",
---- 665=>x"8200", 666=>x"6800", 667=>x"4600", 668=>x"9700",
---- 669=>x"8700", 670=>x"6700", 671=>x"4f00", 672=>x"9f00",
---- 673=>x"8900", 674=>x"6600", 675=>x"5e00", 676=>x"9b00",
---- 677=>x"8500", 678=>x"6600", 679=>x"6200", 680=>x"9f00",
---- 681=>x"8000", 682=>x"6700", 683=>x"6b00", 684=>x"a300",
---- 685=>x"8400", 686=>x"6d00", 687=>x"6600", 688=>x"a600",
---- 689=>x"8500", 690=>x"7100", 691=>x"6f00", 692=>x"a700",
---- 693=>x"8100", 694=>x"7400", 695=>x"7900", 696=>x"a500",
---- 697=>x"7e00", 698=>x"7700", 699=>x"8200", 700=>x"a000",
---- 701=>x"8700", 702=>x"8600", 703=>x"8800", 704=>x"9c00",
---- 705=>x"8d00", 706=>x"8a00", 707=>x"9000", 708=>x"9500",
---- 709=>x"9400", 710=>x"8a00", 711=>x"9500", 712=>x"9700",
---- 713=>x"9d00", 714=>x"8e00", 715=>x"9500", 716=>x"9100",
---- 717=>x"a000", 718=>x"9000", 719=>x"9700", 720=>x"8e00",
---- 721=>x"a300", 722=>x"9600", 723=>x"9a00", 724=>x"9000",
---- 725=>x"a400", 726=>x"9700", 727=>x"9900", 728=>x"8800",
---- 729=>x"a600", 730=>x"9300", 731=>x"9900", 732=>x"8900",
---- 733=>x"ae00", 734=>x"9600", 735=>x"9c00", 736=>x"8600",
---- 737=>x"ac00", 738=>x"6700", 739=>x"9c00", 740=>x"8300",
---- 741=>x"ad00", 742=>x"9e00", 743=>x"9e00", 744=>x"8000",
---- 745=>x"b000", 746=>x"9f00", 747=>x"a300", 748=>x"8400",
---- 749=>x"ae00", 750=>x"9c00", 751=>x"a200", 752=>x"8200",
---- 753=>x"af00", 754=>x"9e00", 755=>x"a000", 756=>x"7d00",
---- 757=>x"b500", 758=>x"9f00", 759=>x"a100", 760=>x"8000",
---- 761=>x"b100", 762=>x"9d00", 763=>x"a300", 764=>x"8200",
---- 765=>x"ae00", 766=>x"9a00", 767=>x"9f00", 768=>x"8d00",
---- 769=>x"ad00", 770=>x"9900", 771=>x"9d00", 772=>x"8c00",
---- 773=>x"ae00", 774=>x"9900", 775=>x"9900", 776=>x"9300",
---- 777=>x"ac00", 778=>x"9700", 779=>x"9200", 780=>x"9900",
---- 781=>x"a300", 782=>x"9a00", 783=>x"8900", 784=>x"9c00",
---- 785=>x"a100", 786=>x"9900", 787=>x"8300", 788=>x"a400",
---- 789=>x"9d00", 790=>x"6b00", 791=>x"8000", 792=>x"aa00",
---- 793=>x"9b00", 794=>x"9000", 795=>x"7e00", 796=>x"a700",
---- 797=>x"9700", 798=>x"8f00", 799=>x"8000", 800=>x"a600",
---- 801=>x"9600", 802=>x"8f00", 803=>x"8800", 804=>x"a500",
---- 805=>x"9500", 806=>x"7500", 807=>x"8b00", 808=>x"a700",
---- 809=>x"9200", 810=>x"8600", 811=>x"8e00", 812=>x"a300",
---- 813=>x"8f00", 814=>x"8900", 815=>x"9500", 816=>x"a100",
---- 817=>x"9000", 818=>x"8600", 819=>x"9500", 820=>x"a000",
---- 821=>x"9000", 822=>x"8800", 823=>x"9400", 824=>x"9900",
---- 825=>x"8e00", 826=>x"8a00", 827=>x"9300", 828=>x"9400",
---- 829=>x"8a00", 830=>x"8d00", 831=>x"9300", 832=>x"9000",
---- 833=>x"8b00", 834=>x"9100", 835=>x"9400", 836=>x"8b00",
---- 837=>x"8800", 838=>x"9000", 839=>x"9100", 840=>x"8600",
---- 841=>x"8900", 842=>x"8f00", 843=>x"9300", 844=>x"8600",
---- 845=>x"8800", 846=>x"9400", 847=>x"9600", 848=>x"8900",
---- 849=>x"8900", 850=>x"9500", 851=>x"9600", 852=>x"8c00",
---- 853=>x"8900", 854=>x"9800", 855=>x"6a00", 856=>x"8d00",
---- 857=>x"8d00", 858=>x"9600", 859=>x"9600", 860=>x"8d00",
---- 861=>x"8f00", 862=>x"9600", 863=>x"9300", 864=>x"8e00",
---- 865=>x"9400", 866=>x"9500", 867=>x"9400", 868=>x"8e00",
---- 869=>x"9700", 870=>x"9400", 871=>x"9500", 872=>x"8f00",
---- 873=>x"9b00", 874=>x"9300", 875=>x"9400", 876=>x"8f00",
---- 877=>x"9900", 878=>x"9600", 879=>x"9000", 880=>x"9100",
---- 881=>x"9400", 882=>x"9700", 883=>x"8f00", 884=>x"9200",
---- 885=>x"9700", 886=>x"9b00", 887=>x"8f00", 888=>x"9100",
---- 889=>x"9000", 890=>x"6700", 891=>x"9500", 892=>x"8f00",
---- 893=>x"9100", 894=>x"9500", 895=>x"9800", 896=>x"9200",
---- 897=>x"9500", 898=>x"9400", 899=>x"9700", 900=>x"9400",
---- 901=>x"9700", 902=>x"9300", 903=>x"9200", 904=>x"8e00",
---- 905=>x"9600", 906=>x"9500", 907=>x"9100", 908=>x"7f00",
---- 909=>x"8900", 910=>x"8c00", 911=>x"8d00", 912=>x"7100",
---- 913=>x"7900", 914=>x"7f00", 915=>x"8000", 916=>x"6000",
---- 917=>x"6b00", 918=>x"6d00", 919=>x"7200", 920=>x"4f00",
---- 921=>x"5f00", 922=>x"5f00", 923=>x"5d00", 924=>x"4500",
---- 925=>x"5200", 926=>x"5000", 927=>x"5000", 928=>x"4800",
---- 929=>x"5000", 930=>x"4500", 931=>x"4700", 932=>x"5300",
---- 933=>x"5c00", 934=>x"4d00", 935=>x"4d00", 936=>x"5800",
---- 937=>x"5d00", 938=>x"5900", 939=>x"5900", 940=>x"5d00",
---- 941=>x"5f00", 942=>x"6200", 943=>x"5d00", 944=>x"5d00",
---- 945=>x"6200", 946=>x"6700", 947=>x"6500", 948=>x"5b00",
---- 949=>x"6200", 950=>x"6a00", 951=>x"6900", 952=>x"5500",
---- 953=>x"6200", 954=>x"6500", 955=>x"6a00", 956=>x"4b00",
---- 957=>x"5d00", 958=>x"6500", 959=>x"6a00", 960=>x"4b00",
---- 961=>x"5900", 962=>x"6300", 963=>x"6b00", 964=>x"5a00",
---- 965=>x"5300", 966=>x"5d00", 967=>x"6300", 968=>x"7300",
---- 969=>x"4d00", 970=>x"5c00", 971=>x"6100", 972=>x"8b00",
---- 973=>x"4a00", 974=>x"5b00", 975=>x"6100", 976=>x"ab00",
---- 977=>x"4e00", 978=>x"5300", 979=>x"5f00", 980=>x"c700",
---- 981=>x"6100", 982=>x"4e00", 983=>x"5a00", 984=>x"d400",
---- 985=>x"7700", 986=>x"4900", 987=>x"5700", 988=>x"db00",
---- 989=>x"9700", 990=>x"4900", 991=>x"5300", 992=>x"d800",
---- 993=>x"b500", 994=>x"5400", 995=>x"4c00", 996=>x"d700",
---- 997=>x"c600", 998=>x"6100", 999=>x"4400", 1000=>x"d500",
---- 1001=>x"d300", 1002=>x"7900", 1003=>x"4000", 1004=>x"d600",
---- 1005=>x"d800", 1006=>x"9800", 1007=>x"4500", 1008=>x"d300",
---- 1009=>x"d900", 1010=>x"b500", 1011=>x"4d00", 1012=>x"d300",
---- 1013=>x"d500", 1014=>x"c900", 1015=>x"6400", 1016=>x"d400",
---- 1017=>x"d500", 1018=>x"2800", 1019=>x"8200", 1020=>x"d300",
---- 1021=>x"d300", 1022=>x"d700", 1023=>x"9b00"),
----
---- 48 => (0=>x"9b00", 1=>x"9c00", 2=>x"9e00", 3=>x"9b00", 4=>x"9a00",
---- 5=>x"9c00", 6=>x"9e00", 7=>x"9b00", 8=>x"9a00",
---- 9=>x"9c00", 10=>x"9e00", 11=>x"9b00", 12=>x"9700",
---- 13=>x"9a00", 14=>x"9b00", 15=>x"9a00", 16=>x"9b00",
---- 17=>x"9b00", 18=>x"9a00", 19=>x"9a00", 20=>x"6500",
---- 21=>x"9c00", 22=>x"9800", 23=>x"9a00", 24=>x"9900",
---- 25=>x"9900", 26=>x"9800", 27=>x"9900", 28=>x"9b00",
---- 29=>x"9b00", 30=>x"9800", 31=>x"9800", 32=>x"9900",
---- 33=>x"9b00", 34=>x"9b00", 35=>x"9700", 36=>x"6700",
---- 37=>x"9b00", 38=>x"9b00", 39=>x"9900", 40=>x"9d00",
---- 41=>x"9c00", 42=>x"9900", 43=>x"9800", 44=>x"9a00",
---- 45=>x"9a00", 46=>x"9700", 47=>x"9a00", 48=>x"9b00",
---- 49=>x"9a00", 50=>x"9900", 51=>x"9700", 52=>x"9b00",
---- 53=>x"9a00", 54=>x"9900", 55=>x"9900", 56=>x"9d00",
---- 57=>x"9a00", 58=>x"9c00", 59=>x"9a00", 60=>x"9d00",
---- 61=>x"6400", 62=>x"9b00", 63=>x"9c00", 64=>x"9e00",
---- 65=>x"9d00", 66=>x"9b00", 67=>x"9c00", 68=>x"9d00",
---- 69=>x"9d00", 70=>x"9c00", 71=>x"9a00", 72=>x"9d00",
---- 73=>x"9c00", 74=>x"9c00", 75=>x"9b00", 76=>x"9c00",
---- 77=>x"9e00", 78=>x"9e00", 79=>x"9d00", 80=>x"9a00",
---- 81=>x"9c00", 82=>x"9f00", 83=>x"9d00", 84=>x"9900",
---- 85=>x"9800", 86=>x"9900", 87=>x"9c00", 88=>x"9b00",
---- 89=>x"9a00", 90=>x"9700", 91=>x"9c00", 92=>x"9b00",
---- 93=>x"9b00", 94=>x"9900", 95=>x"9900", 96=>x"9900",
---- 97=>x"9b00", 98=>x"9700", 99=>x"9600", 100=>x"9a00",
---- 101=>x"9b00", 102=>x"9600", 103=>x"9800", 104=>x"9700",
---- 105=>x"9800", 106=>x"9700", 107=>x"9700", 108=>x"9300",
---- 109=>x"9500", 110=>x"9400", 111=>x"9400", 112=>x"9100",
---- 113=>x"9400", 114=>x"9200", 115=>x"9200", 116=>x"9100",
---- 117=>x"9100", 118=>x"9200", 119=>x"9100", 120=>x"9100",
---- 121=>x"8f00", 122=>x"9100", 123=>x"9200", 124=>x"8e00",
---- 125=>x"8f00", 126=>x"9000", 127=>x"9100", 128=>x"8c00",
---- 129=>x"8e00", 130=>x"8e00", 131=>x"8f00", 132=>x"8b00",
---- 133=>x"8f00", 134=>x"8d00", 135=>x"8e00", 136=>x"8d00",
---- 137=>x"8d00", 138=>x"8e00", 139=>x"9000", 140=>x"8e00",
---- 141=>x"8f00", 142=>x"9100", 143=>x"9000", 144=>x"8f00",
---- 145=>x"8e00", 146=>x"9000", 147=>x"8f00", 148=>x"9000",
---- 149=>x"8e00", 150=>x"9000", 151=>x"9300", 152=>x"9100",
---- 153=>x"8f00", 154=>x"9100", 155=>x"9300", 156=>x"9200",
---- 157=>x"9100", 158=>x"9100", 159=>x"9100", 160=>x"9400",
---- 161=>x"9300", 162=>x"8e00", 163=>x"9100", 164=>x"9600",
---- 165=>x"9300", 166=>x"9000", 167=>x"8d00", 168=>x"9400",
---- 169=>x"9300", 170=>x"9400", 171=>x"9000", 172=>x"9200",
---- 173=>x"9400", 174=>x"9400", 175=>x"9000", 176=>x"8f00",
---- 177=>x"9500", 178=>x"9600", 179=>x"9400", 180=>x"8c00",
---- 181=>x"9300", 182=>x"9400", 183=>x"9600", 184=>x"8600",
---- 185=>x"9000", 186=>x"9300", 187=>x"9600", 188=>x"8200",
---- 189=>x"8c00", 190=>x"6f00", 191=>x"9500", 192=>x"7b00",
---- 193=>x"8600", 194=>x"8b00", 195=>x"9300", 196=>x"7300",
---- 197=>x"7e00", 198=>x"8600", 199=>x"8f00", 200=>x"6500",
---- 201=>x"7800", 202=>x"8100", 203=>x"8700", 204=>x"5d00",
---- 205=>x"6b00", 206=>x"7d00", 207=>x"8600", 208=>x"4b00",
---- 209=>x"5e00", 210=>x"8800", 211=>x"7f00", 212=>x"c500",
---- 213=>x"5300", 214=>x"6500", 215=>x"7800", 216=>x"2f00",
---- 217=>x"4100", 218=>x"5800", 219=>x"6d00", 220=>x"2900",
---- 221=>x"2f00", 222=>x"4400", 223=>x"5a00", 224=>x"2700",
---- 225=>x"2600", 226=>x"2f00", 227=>x"4000", 228=>x"2500",
---- 229=>x"2400", 230=>x"2200", 231=>x"4d00", 232=>x"2700",
---- 233=>x"2000", 234=>x"5100", 235=>x"b400", 236=>x"2800",
---- 237=>x"6a00", 238=>x"3f00", 239=>x"df00", 240=>x"8400",
---- 241=>x"ce00", 242=>x"de00", 243=>x"d600", 244=>x"d500",
---- 245=>x"d900", 246=>x"c900", 247=>x"a600", 248=>x"d900",
---- 249=>x"bc00", 250=>x"9f00", 251=>x"b200", 252=>x"af00",
---- 253=>x"9b00", 254=>x"c100", 255=>x"d600", 256=>x"a200",
---- 257=>x"c300", 258=>x"d700", 259=>x"d700", 260=>x"d000",
---- 261=>x"d900", 262=>x"d800", 263=>x"d500", 264=>x"2900",
---- 265=>x"d800", 266=>x"2e00", 267=>x"cf00", 268=>x"d400",
---- 269=>x"d200", 270=>x"ce00", 271=>x"cb00", 272=>x"d100",
---- 273=>x"ce00", 274=>x"cb00", 275=>x"cc00", 276=>x"cd00",
---- 277=>x"c800", 278=>x"ca00", 279=>x"c900", 280=>x"c800",
---- 281=>x"c900", 282=>x"c800", 283=>x"cb00", 284=>x"c900",
---- 285=>x"c800", 286=>x"c900", 287=>x"cb00", 288=>x"c800",
---- 289=>x"ca00", 290=>x"cd00", 291=>x"ce00", 292=>x"c800",
---- 293=>x"cb00", 294=>x"cd00", 295=>x"cd00", 296=>x"ca00",
---- 297=>x"cb00", 298=>x"ca00", 299=>x"cd00", 300=>x"ca00",
---- 301=>x"cd00", 302=>x"cc00", 303=>x"cc00", 304=>x"cc00",
---- 305=>x"cb00", 306=>x"cd00", 307=>x"d100", 308=>x"ca00",
---- 309=>x"ce00", 310=>x"cd00", 311=>x"c700", 312=>x"cf00",
---- 313=>x"cc00", 314=>x"cd00", 315=>x"b500", 316=>x"ce00",
---- 317=>x"cd00", 318=>x"c400", 319=>x"a200", 320=>x"ce00",
---- 321=>x"d000", 322=>x"aa00", 323=>x"9900", 324=>x"d200",
---- 325=>x"bd00", 326=>x"9800", 327=>x"9e00", 328=>x"cf00",
---- 329=>x"a300", 330=>x"9600", 331=>x"a700", 332=>x"b300",
---- 333=>x"9200", 334=>x"9f00", 335=>x"af00", 336=>x"9600",
---- 337=>x"9e00", 338=>x"ac00", 339=>x"9700", 340=>x"9800",
---- 341=>x"a700", 342=>x"9800", 343=>x"9700", 344=>x"a500",
---- 345=>x"9c00", 346=>x"8d00", 347=>x"6a00", 348=>x"9200",
---- 349=>x"7300", 350=>x"5100", 351=>x"5000", 352=>x"5b00",
---- 353=>x"4d00", 354=>x"5700", 355=>x"5f00", 356=>x"5200",
---- 357=>x"5700", 358=>x"5c00", 359=>x"5e00", 360=>x"5700",
---- 361=>x"5c00", 362=>x"5900", 363=>x"9b00", 364=>x"5a00",
---- 365=>x"6600", 366=>x"7200", 367=>x"8900", 368=>x"6700",
---- 369=>x"8100", 370=>x"9800", 371=>x"ad00", 372=>x"8d00",
---- 373=>x"a600", 374=>x"b800", 375=>x"c200", 376=>x"a700",
---- 377=>x"b500", 378=>x"bf00", 379=>x"3500", 380=>x"b000",
---- 381=>x"b400", 382=>x"c500", 383=>x"c800", 384=>x"b000",
---- 385=>x"c300", 386=>x"3400", 387=>x"6100", 388=>x"c400",
---- 389=>x"d300", 390=>x"6a00", 391=>x"1f00", 392=>x"d200",
---- 393=>x"7700", 394=>x"2500", 395=>x"2900", 396=>x"7900",
---- 397=>x"2000", 398=>x"2b00", 399=>x"2900", 400=>x"2b00",
---- 401=>x"2600", 402=>x"2b00", 403=>x"2b00", 404=>x"2d00",
---- 405=>x"2600", 406=>x"2800", 407=>x"2e00", 408=>x"2e00",
---- 409=>x"2900", 410=>x"2c00", 411=>x"2f00", 412=>x"2d00",
---- 413=>x"2b00", 414=>x"3100", 415=>x"3500", 416=>x"2a00",
---- 417=>x"2e00", 418=>x"3600", 419=>x"3700", 420=>x"2f00",
---- 421=>x"2f00", 422=>x"3300", 423=>x"3800", 424=>x"3100",
---- 425=>x"3500", 426=>x"3500", 427=>x"3700", 428=>x"3600",
---- 429=>x"3b00", 430=>x"3700", 431=>x"3600", 432=>x"2f00",
---- 433=>x"3700", 434=>x"3700", 435=>x"3900", 436=>x"3400",
---- 437=>x"ca00", 438=>x"3900", 439=>x"3b00", 440=>x"3300",
---- 441=>x"3700", 442=>x"3900", 443=>x"3800", 444=>x"3400",
---- 445=>x"3700", 446=>x"3700", 447=>x"3800", 448=>x"3700",
---- 449=>x"3700", 450=>x"3700", 451=>x"3900", 452=>x"3700",
---- 453=>x"3800", 454=>x"3900", 455=>x"3c00", 456=>x"3900",
---- 457=>x"3b00", 458=>x"c400", 459=>x"3a00", 460=>x"3b00",
---- 461=>x"3a00", 462=>x"3c00", 463=>x"3d00", 464=>x"3a00",
---- 465=>x"3b00", 466=>x"3b00", 467=>x"3b00", 468=>x"3b00",
---- 469=>x"3900", 470=>x"3900", 471=>x"3a00", 472=>x"3e00",
---- 473=>x"3d00", 474=>x"3c00", 475=>x"3f00", 476=>x"3a00",
---- 477=>x"3f00", 478=>x"4100", 479=>x"4000", 480=>x"3c00",
---- 481=>x"3c00", 482=>x"4300", 483=>x"3e00", 484=>x"3c00",
---- 485=>x"3f00", 486=>x"3e00", 487=>x"3f00", 488=>x"3e00",
---- 489=>x"4700", 490=>x"4a00", 491=>x"3b00", 492=>x"3e00",
---- 493=>x"4600", 494=>x"4300", 495=>x"3800", 496=>x"3e00",
---- 497=>x"4000", 498=>x"3900", 499=>x"3600", 500=>x"4200",
---- 501=>x"3e00", 502=>x"3800", 503=>x"2f00", 504=>x"4000",
---- 505=>x"4200", 506=>x"3700", 507=>x"3100", 508=>x"4100",
---- 509=>x"4100", 510=>x"3500", 511=>x"3100", 512=>x"4000",
---- 513=>x"3800", 514=>x"3300", 515=>x"3000", 516=>x"3f00",
---- 517=>x"3700", 518=>x"3000", 519=>x"3100", 520=>x"3d00",
---- 521=>x"3300", 522=>x"2d00", 523=>x"3000", 524=>x"3800",
---- 525=>x"3000", 526=>x"2e00", 527=>x"3200", 528=>x"3d00",
---- 529=>x"2e00", 530=>x"2e00", 531=>x"3200", 532=>x"ca00",
---- 533=>x"3000", 534=>x"3000", 535=>x"3400", 536=>x"3300",
---- 537=>x"2e00", 538=>x"3200", 539=>x"3200", 540=>x"3400",
---- 541=>x"3300", 542=>x"3500", 543=>x"3200", 544=>x"3200",
---- 545=>x"3200", 546=>x"3100", 547=>x"2f00", 548=>x"2b00",
---- 549=>x"2f00", 550=>x"2d00", 551=>x"2e00", 552=>x"2e00",
---- 553=>x"3100", 554=>x"3000", 555=>x"2d00", 556=>x"3000",
---- 557=>x"3400", 558=>x"2c00", 559=>x"3200", 560=>x"2f00",
---- 561=>x"2f00", 562=>x"2900", 563=>x"3c00", 564=>x"3400",
---- 565=>x"3000", 566=>x"2e00", 567=>x"4100", 568=>x"3300",
---- 569=>x"2d00", 570=>x"3000", 571=>x"c700", 572=>x"3100",
---- 573=>x"2500", 574=>x"3200", 575=>x"3600", 576=>x"3200",
---- 577=>x"2c00", 578=>x"3300", 579=>x"3400", 580=>x"2f00",
---- 581=>x"2a00", 582=>x"3700", 583=>x"3200", 584=>x"2e00",
---- 585=>x"2f00", 586=>x"3700", 587=>x"2f00", 588=>x"2d00",
---- 589=>x"3100", 590=>x"3500", 591=>x"2b00", 592=>x"3700",
---- 593=>x"3200", 594=>x"3300", 595=>x"2d00", 596=>x"4000",
---- 597=>x"3600", 598=>x"3200", 599=>x"2b00", 600=>x"3e00",
---- 601=>x"3b00", 602=>x"3200", 603=>x"2c00", 604=>x"3c00",
---- 605=>x"3b00", 606=>x"3300", 607=>x"3100", 608=>x"3800",
---- 609=>x"3700", 610=>x"2f00", 611=>x"2b00", 612=>x"3a00",
---- 613=>x"3500", 614=>x"2b00", 615=>x"3300", 616=>x"3600",
---- 617=>x"2e00", 618=>x"2700", 619=>x"3f00", 620=>x"3000",
---- 621=>x"2c00", 622=>x"2c00", 623=>x"4d00", 624=>x"2b00",
---- 625=>x"2b00", 626=>x"3700", 627=>x"5a00", 628=>x"2500",
---- 629=>x"2500", 630=>x"4000", 631=>x"6800", 632=>x"2400",
---- 633=>x"2700", 634=>x"4c00", 635=>x"7900", 636=>x"2200",
---- 637=>x"2400", 638=>x"5700", 639=>x"8600", 640=>x"2400",
---- 641=>x"2500", 642=>x"5c00", 643=>x"8f00", 644=>x"2a00",
---- 645=>x"3200", 646=>x"7000", 647=>x"9100", 648=>x"3300",
---- 649=>x"4500", 650=>x"7d00", 651=>x"9500", 652=>x"3000",
---- 653=>x"5d00", 654=>x"8700", 655=>x"9400", 656=>x"2d00",
---- 657=>x"6d00", 658=>x"8e00", 659=>x"9500", 660=>x"3400",
---- 661=>x"7a00", 662=>x"9200", 663=>x"9200", 664=>x"4900",
---- 665=>x"8200", 666=>x"9400", 667=>x"9100", 668=>x"5e00",
---- 669=>x"8800", 670=>x"9400", 671=>x"9000", 672=>x"6c00",
---- 673=>x"8d00", 674=>x"9500", 675=>x"8d00", 676=>x"7900",
---- 677=>x"8e00", 678=>x"9400", 679=>x"9000", 680=>x"8500",
---- 681=>x"8d00", 682=>x"9000", 683=>x"9100", 684=>x"8a00",
---- 685=>x"8c00", 686=>x"8f00", 687=>x"9300", 688=>x"8c00",
---- 689=>x"8c00", 690=>x"9000", 691=>x"9100", 692=>x"8f00",
---- 693=>x"9100", 694=>x"9000", 695=>x"9000", 696=>x"9500",
---- 697=>x"9100", 698=>x"9300", 699=>x"8e00", 700=>x"9200",
---- 701=>x"9000", 702=>x"9500", 703=>x"9300", 704=>x"9500",
---- 705=>x"9300", 706=>x"9600", 707=>x"9300", 708=>x"9500",
---- 709=>x"9300", 710=>x"9500", 711=>x"9500", 712=>x"9600",
---- 713=>x"9300", 714=>x"9500", 715=>x"9700", 716=>x"9a00",
---- 717=>x"9400", 718=>x"9600", 719=>x"9500", 720=>x"9900",
---- 721=>x"9600", 722=>x"9500", 723=>x"9700", 724=>x"9900",
---- 725=>x"9800", 726=>x"9700", 727=>x"9a00", 728=>x"9a00",
---- 729=>x"9500", 730=>x"9500", 731=>x"9a00", 732=>x"9800",
---- 733=>x"9300", 734=>x"9600", 735=>x"9b00", 736=>x"9900",
---- 737=>x"9100", 738=>x"9900", 739=>x"9900", 740=>x"9700",
---- 741=>x"8e00", 742=>x"9c00", 743=>x"9a00", 744=>x"9400",
---- 745=>x"9100", 746=>x"9b00", 747=>x"9d00", 748=>x"9200",
---- 749=>x"9300", 750=>x"9800", 751=>x"9f00", 752=>x"9200",
---- 753=>x"9400", 754=>x"9700", 755=>x"9f00", 756=>x"9500",
---- 757=>x"9100", 758=>x"9a00", 759=>x"9e00", 760=>x"9700",
---- 761=>x"9200", 762=>x"9700", 763=>x"9700", 764=>x"9400",
---- 765=>x"8d00", 766=>x"8c00", 767=>x"9000", 768=>x"8e00",
---- 769=>x"8100", 770=>x"7e00", 771=>x"8400", 772=>x"8300",
---- 773=>x"7900", 774=>x"7100", 775=>x"7600", 776=>x"7500",
---- 777=>x"7600", 778=>x"6e00", 779=>x"6e00", 780=>x"7000",
---- 781=>x"7200", 782=>x"7200", 783=>x"6900", 784=>x"7200",
---- 785=>x"7200", 786=>x"7a00", 787=>x"7200", 788=>x"7800",
---- 789=>x"7f00", 790=>x"7f00", 791=>x"8200", 792=>x"7c00",
---- 793=>x"8800", 794=>x"8100", 795=>x"8600", 796=>x"8600",
---- 797=>x"8a00", 798=>x"8400", 799=>x"8700", 800=>x"8e00",
---- 801=>x"8b00", 802=>x"8a00", 803=>x"8a00", 804=>x"9300",
---- 805=>x"8f00", 806=>x"8d00", 807=>x"8c00", 808=>x"9500",
---- 809=>x"9200", 810=>x"9100", 811=>x"9100", 812=>x"9700",
---- 813=>x"9400", 814=>x"9100", 815=>x"9200", 816=>x"9500",
---- 817=>x"9400", 818=>x"9200", 819=>x"9100", 820=>x"9500",
---- 821=>x"9700", 822=>x"9100", 823=>x"9100", 824=>x"6c00",
---- 825=>x"9600", 826=>x"9300", 827=>x"9100", 828=>x"9600",
---- 829=>x"9600", 830=>x"9400", 831=>x"9200", 832=>x"9400",
---- 833=>x"9400", 834=>x"9100", 835=>x"9000", 836=>x"9200",
---- 837=>x"9300", 838=>x"9400", 839=>x"9200", 840=>x"9300",
---- 841=>x"9000", 842=>x"9300", 843=>x"9100", 844=>x"9200",
---- 845=>x"9300", 846=>x"9100", 847=>x"9100", 848=>x"9200",
---- 849=>x"9200", 850=>x"9000", 851=>x"9100", 852=>x"9300",
---- 853=>x"9400", 854=>x"9100", 855=>x"9200", 856=>x"9500",
---- 857=>x"9900", 858=>x"9100", 859=>x"9100", 860=>x"9500",
---- 861=>x"9500", 862=>x"9200", 863=>x"9200", 864=>x"9200",
---- 865=>x"6c00", 866=>x"9100", 867=>x"9300", 868=>x"9200",
---- 869=>x"9100", 870=>x"9100", 871=>x"8e00", 872=>x"9300",
---- 873=>x"9100", 874=>x"8f00", 875=>x"9000", 876=>x"9100",
---- 877=>x"9200", 878=>x"9200", 879=>x"9000", 880=>x"6e00",
---- 881=>x"9000", 882=>x"9000", 883=>x"8f00", 884=>x"8d00",
---- 885=>x"8f00", 886=>x"8f00", 887=>x"8d00", 888=>x"9000",
---- 889=>x"8e00", 890=>x"8e00", 891=>x"8c00", 892=>x"8f00",
---- 893=>x"8f00", 894=>x"8f00", 895=>x"8f00", 896=>x"8d00",
---- 897=>x"9000", 898=>x"8f00", 899=>x"9000", 900=>x"9000",
---- 901=>x"8f00", 902=>x"8e00", 903=>x"8e00", 904=>x"9000",
---- 905=>x"8e00", 906=>x"8f00", 907=>x"8f00", 908=>x"8e00",
---- 909=>x"9100", 910=>x"9000", 911=>x"9300", 912=>x"8500",
---- 913=>x"8900", 914=>x"8900", 915=>x"8e00", 916=>x"7400",
---- 917=>x"7c00", 918=>x"7e00", 919=>x"8400", 920=>x"6600",
---- 921=>x"6a00", 922=>x"7000", 923=>x"7900", 924=>x"5700",
---- 925=>x"5d00", 926=>x"6200", 927=>x"6500", 928=>x"4800",
---- 929=>x"4e00", 930=>x"5500", 931=>x"5300", 932=>x"b300",
---- 933=>x"4a00", 934=>x"4d00", 935=>x"4c00", 936=>x"5400",
---- 937=>x"5200", 938=>x"5200", 939=>x"4c00", 940=>x"5a00",
---- 941=>x"5b00", 942=>x"5700", 943=>x"5300", 944=>x"6400",
---- 945=>x"6100", 946=>x"5e00", 947=>x"5900", 948=>x"6800",
---- 949=>x"6700", 950=>x"6500", 951=>x"5f00", 952=>x"9400",
---- 953=>x"6b00", 954=>x"6900", 955=>x"6400", 956=>x"6900",
---- 957=>x"9200", 958=>x"6b00", 959=>x"6700", 960=>x"6b00",
---- 961=>x"6b00", 962=>x"6c00", 963=>x"6900", 964=>x"6900",
---- 965=>x"7000", 966=>x"6e00", 967=>x"6800", 968=>x"6500",
---- 969=>x"6b00", 970=>x"6b00", 971=>x"6900", 972=>x"6300",
---- 973=>x"6600", 974=>x"6800", 975=>x"6500", 976=>x"6200",
---- 977=>x"6500", 978=>x"6300", 979=>x"6600", 980=>x"5e00",
---- 981=>x"6300", 982=>x"6200", 983=>x"6600", 984=>x"5800",
---- 985=>x"5f00", 986=>x"6200", 987=>x"6200", 988=>x"5600",
---- 989=>x"5c00", 990=>x"6100", 991=>x"6300", 992=>x"5600",
---- 993=>x"5800", 994=>x"5f00", 995=>x"6100", 996=>x"5500",
---- 997=>x"5a00", 998=>x"5e00", 999=>x"6300", 1000=>x"5300",
---- 1001=>x"5600", 1002=>x"5c00", 1003=>x"6400", 1004=>x"5100",
---- 1005=>x"5400", 1006=>x"5a00", 1007=>x"5f00", 1008=>x"4a00",
---- 1009=>x"5200", 1010=>x"5e00", 1011=>x"6500", 1012=>x"4600",
---- 1013=>x"5200", 1014=>x"5500", 1015=>x"5800", 1016=>x"4a00",
---- 1017=>x"5600", 1018=>x"5800", 1019=>x"5e00", 1020=>x"6800",
---- 1021=>x"6400", 1022=>x"5a00", 1023=>x"5c00"),
----
---- 49 => (0=>x"9c00", 1=>x"a000", 2=>x"9d00", 3=>x"9b00", 4=>x"9c00",
---- 5=>x"a000", 6=>x"9c00", 7=>x"9b00", 8=>x"9c00",
---- 9=>x"9e00", 10=>x"9d00", 11=>x"9b00", 12=>x"9c00",
---- 13=>x"9b00", 14=>x"9c00", 15=>x"9a00", 16=>x"9b00",
---- 17=>x"9c00", 18=>x"9900", 19=>x"9a00", 20=>x"9900",
---- 21=>x"9900", 22=>x"9900", 23=>x"9800", 24=>x"9900",
---- 25=>x"9a00", 26=>x"9a00", 27=>x"9800", 28=>x"9500",
---- 29=>x"9800", 30=>x"9900", 31=>x"9900", 32=>x"9800",
---- 33=>x"9500", 34=>x"9900", 35=>x"9800", 36=>x"9800",
---- 37=>x"9700", 38=>x"9800", 39=>x"9800", 40=>x"9700",
---- 41=>x"9700", 42=>x"9700", 43=>x"9b00", 44=>x"9700",
---- 45=>x"9800", 46=>x"9700", 47=>x"9700", 48=>x"9700",
---- 49=>x"9800", 50=>x"9700", 51=>x"9700", 52=>x"9900",
---- 53=>x"9900", 54=>x"9800", 55=>x"9800", 56=>x"9a00",
---- 57=>x"9c00", 58=>x"6300", 59=>x"9600", 60=>x"9c00",
---- 61=>x"6200", 62=>x"9b00", 63=>x"9b00", 64=>x"9d00",
---- 65=>x"9d00", 66=>x"9a00", 67=>x"9b00", 68=>x"9c00",
---- 69=>x"9a00", 70=>x"9b00", 71=>x"9e00", 72=>x"9d00",
---- 73=>x"9b00", 74=>x"9a00", 75=>x"9b00", 76=>x"9c00",
---- 77=>x"9d00", 78=>x"9b00", 79=>x"9a00", 80=>x"9b00",
---- 81=>x"9b00", 82=>x"9c00", 83=>x"9900", 84=>x"9d00",
---- 85=>x"9b00", 86=>x"9a00", 87=>x"9800", 88=>x"9b00",
---- 89=>x"9800", 90=>x"6700", 91=>x"9600", 92=>x"9800",
---- 93=>x"9800", 94=>x"9600", 95=>x"9500", 96=>x"9700",
---- 97=>x"9800", 98=>x"9600", 99=>x"9400", 100=>x"9800",
---- 101=>x"9400", 102=>x"9300", 103=>x"9400", 104=>x"9300",
---- 105=>x"9100", 106=>x"9200", 107=>x"9100", 108=>x"9200",
---- 109=>x"9100", 110=>x"8f00", 111=>x"8e00", 112=>x"9100",
---- 113=>x"9100", 114=>x"9000", 115=>x"9100", 116=>x"9300",
---- 117=>x"9000", 118=>x"8f00", 119=>x"8f00", 120=>x"9200",
---- 121=>x"9300", 122=>x"9000", 123=>x"8f00", 124=>x"9200",
---- 125=>x"9200", 126=>x"8e00", 127=>x"9000", 128=>x"8f00",
---- 129=>x"8f00", 130=>x"8f00", 131=>x"9000", 132=>x"8e00",
---- 133=>x"9300", 134=>x"9300", 135=>x"8e00", 136=>x"9100",
---- 137=>x"9200", 138=>x"9300", 139=>x"8f00", 140=>x"9100",
---- 141=>x"9100", 142=>x"9300", 143=>x"8f00", 144=>x"9100",
---- 145=>x"9200", 146=>x"9000", 147=>x"8f00", 148=>x"9300",
---- 149=>x"9500", 150=>x"9400", 151=>x"8e00", 152=>x"9400",
---- 153=>x"9500", 154=>x"9400", 155=>x"8f00", 156=>x"9200",
---- 157=>x"9300", 158=>x"9200", 159=>x"8f00", 160=>x"8f00",
---- 161=>x"9100", 162=>x"9200", 163=>x"9000", 164=>x"9000",
---- 165=>x"9200", 166=>x"9200", 167=>x"9000", 168=>x"9100",
---- 169=>x"9400", 170=>x"9300", 171=>x"9200", 172=>x"8e00",
---- 173=>x"8f00", 174=>x"9200", 175=>x"9300", 176=>x"8f00",
---- 177=>x"9000", 178=>x"9000", 179=>x"9200", 180=>x"9100",
---- 181=>x"8f00", 182=>x"9200", 183=>x"9100", 184=>x"9500",
---- 185=>x"8f00", 186=>x"9200", 187=>x"9000", 188=>x"9600",
---- 189=>x"9300", 190=>x"9000", 191=>x"9200", 192=>x"9500",
---- 193=>x"9400", 194=>x"9100", 195=>x"8f00", 196=>x"9300",
---- 197=>x"9500", 198=>x"9300", 199=>x"9100", 200=>x"9200",
---- 201=>x"9500", 202=>x"9300", 203=>x"9200", 204=>x"8d00",
---- 205=>x"9400", 206=>x"9400", 207=>x"9200", 208=>x"8700",
---- 209=>x"8f00", 210=>x"6d00", 211=>x"9400", 212=>x"8200",
---- 213=>x"8900", 214=>x"8f00", 215=>x"9300", 216=>x"7900",
---- 217=>x"8200", 218=>x"8900", 219=>x"8d00", 220=>x"6a00",
---- 221=>x"7200", 222=>x"8300", 223=>x"9500", 224=>x"5800",
---- 225=>x"8a00", 226=>x"b700", 227=>x"ca00", 228=>x"a200",
---- 229=>x"d100", 230=>x"dc00", 231=>x"dd00", 232=>x"dc00",
---- 233=>x"dd00", 234=>x"d500", 235=>x"c300", 236=>x"db00",
---- 237=>x"c400", 238=>x"b900", 239=>x"c400", 240=>x"b300",
---- 241=>x"af00", 242=>x"cd00", 243=>x"d900", 244=>x"b200",
---- 245=>x"d300", 246=>x"da00", 247=>x"2400", 248=>x"d600",
---- 249=>x"db00", 250=>x"da00", 251=>x"d600", 252=>x"db00",
---- 253=>x"da00", 254=>x"d600", 255=>x"d300", 256=>x"2900",
---- 257=>x"d400", 258=>x"d500", 259=>x"d100", 260=>x"d400",
---- 261=>x"d100", 262=>x"d000", 263=>x"ca00", 264=>x"d100",
---- 265=>x"ce00", 266=>x"cb00", 267=>x"c800", 268=>x"ce00",
---- 269=>x"ca00", 270=>x"c800", 271=>x"c800", 272=>x"cc00",
---- 273=>x"c800", 274=>x"c800", 275=>x"cb00", 276=>x"c800",
---- 277=>x"ca00", 278=>x"cb00", 279=>x"cc00", 280=>x"cc00",
---- 281=>x"cd00", 282=>x"cb00", 283=>x"cb00", 284=>x"cd00",
---- 285=>x"cc00", 286=>x"cc00", 287=>x"cc00", 288=>x"cd00",
---- 289=>x"cb00", 290=>x"cb00", 291=>x"c900", 292=>x"cb00",
---- 293=>x"cc00", 294=>x"c900", 295=>x"c300", 296=>x"cd00",
---- 297=>x"cb00", 298=>x"bf00", 299=>x"c100", 300=>x"d000",
---- 301=>x"bd00", 302=>x"b200", 303=>x"bc00", 304=>x"c000",
---- 305=>x"a900", 306=>x"a800", 307=>x"b200", 308=>x"ac00",
---- 309=>x"9f00", 310=>x"a200", 311=>x"a700", 312=>x"a200",
---- 313=>x"9c00", 314=>x"9a00", 315=>x"5600", 316=>x"9900",
---- 317=>x"9d00", 318=>x"a900", 319=>x"bc00", 320=>x"9c00",
---- 321=>x"aa00", 322=>x"bd00", 323=>x"9900", 324=>x"ab00",
---- 325=>x"b700", 326=>x"9a00", 327=>x"8000", 328=>x"b700",
---- 329=>x"9c00", 330=>x"8600", 331=>x"9d00", 332=>x"9700",
---- 333=>x"8f00", 334=>x"a900", 335=>x"ab00", 336=>x"9700",
---- 337=>x"a600", 338=>x"9700", 339=>x"7c00", 340=>x"8b00",
---- 341=>x"7500", 342=>x"5d00", 343=>x"6700", 344=>x"4f00",
---- 345=>x"5900", 346=>x"5f00", 347=>x"7a00", 348=>x"5700",
---- 349=>x"6200", 350=>x"6f00", 351=>x"6800", 352=>x"6000",
---- 353=>x"6b00", 354=>x"8900", 355=>x"b500", 356=>x"6600",
---- 357=>x"8200", 358=>x"b000", 359=>x"c700", 360=>x"8600",
---- 361=>x"a900", 362=>x"bf00", 363=>x"cc00", 364=>x"ae00",
---- 365=>x"ba00", 366=>x"c900", 367=>x"db00", 368=>x"be00",
---- 369=>x"cd00", 370=>x"b900", 371=>x"6d00", 372=>x"cd00",
---- 373=>x"ba00", 374=>x"4400", 375=>x"2100", 376=>x"d100",
---- 377=>x"5f00", 378=>x"1f00", 379=>x"3000", 380=>x"6b00",
---- 381=>x"2400", 382=>x"2e00", 383=>x"3100", 384=>x"2300",
---- 385=>x"2a00", 386=>x"2b00", 387=>x"2d00", 388=>x"2a00",
---- 389=>x"2b00", 390=>x"2e00", 391=>x"3200", 392=>x"2700",
---- 393=>x"2b00", 394=>x"3000", 395=>x"3300", 396=>x"2c00",
---- 397=>x"2f00", 398=>x"3100", 399=>x"3300", 400=>x"2f00",
---- 401=>x"3000", 402=>x"3500", 403=>x"3300", 404=>x"2e00",
---- 405=>x"3100", 406=>x"3300", 407=>x"3700", 408=>x"3500",
---- 409=>x"3300", 410=>x"3000", 411=>x"3600", 412=>x"3700",
---- 413=>x"3700", 414=>x"3200", 415=>x"3400", 416=>x"3900",
---- 417=>x"3400", 418=>x"3300", 419=>x"3600", 420=>x"3900",
---- 421=>x"3700", 422=>x"3700", 423=>x"3b00", 424=>x"3a00",
---- 425=>x"3a00", 426=>x"ca00", 427=>x"3800", 428=>x"3800",
---- 429=>x"3d00", 430=>x"3c00", 431=>x"3d00", 432=>x"3700",
---- 433=>x"3600", 434=>x"3c00", 435=>x"3c00", 436=>x"3800",
---- 437=>x"4100", 438=>x"3e00", 439=>x"3d00", 440=>x"3c00",
---- 441=>x"3f00", 442=>x"3e00", 443=>x"3c00", 444=>x"3b00",
---- 445=>x"3c00", 446=>x"4200", 447=>x"3800", 448=>x"3d00",
---- 449=>x"3f00", 450=>x"3e00", 451=>x"3300", 452=>x"4100",
---- 453=>x"4100", 454=>x"3b00", 455=>x"cb00", 456=>x"4100",
---- 457=>x"4000", 458=>x"3700", 459=>x"3200", 460=>x"4100",
---- 461=>x"3f00", 462=>x"3800", 463=>x"2f00", 464=>x"4200",
---- 465=>x"3e00", 466=>x"3800", 467=>x"2f00", 468=>x"3d00",
---- 469=>x"3900", 470=>x"3700", 471=>x"3300", 472=>x"3d00",
---- 473=>x"3400", 474=>x"3000", 475=>x"3400", 476=>x"3e00",
---- 477=>x"3300", 478=>x"2c00", 479=>x"3000", 480=>x"3a00",
---- 481=>x"3300", 482=>x"3100", 483=>x"3500", 484=>x"3500",
---- 485=>x"2e00", 486=>x"3400", 487=>x"3500", 488=>x"3400",
---- 489=>x"3000", 490=>x"3200", 491=>x"3000", 492=>x"3000",
---- 493=>x"3000", 494=>x"3200", 495=>x"3300", 496=>x"3400",
---- 497=>x"3000", 498=>x"3300", 499=>x"3300", 500=>x"3300",
---- 501=>x"3000", 502=>x"2e00", 503=>x"2f00", 504=>x"3000",
---- 505=>x"3300", 506=>x"cb00", 507=>x"3400", 508=>x"3200",
---- 509=>x"3500", 510=>x"3400", 511=>x"3500", 512=>x"3000",
---- 513=>x"3200", 514=>x"3200", 515=>x"3600", 516=>x"3300",
---- 517=>x"2f00", 518=>x"3200", 519=>x"ca00", 520=>x"3200",
---- 521=>x"3200", 522=>x"3800", 523=>x"3800", 524=>x"3100",
---- 525=>x"3200", 526=>x"3400", 527=>x"3500", 528=>x"3400",
---- 529=>x"3600", 530=>x"3200", 531=>x"2f00", 532=>x"3000",
---- 533=>x"3500", 534=>x"2f00", 535=>x"2c00", 536=>x"3400",
---- 537=>x"3300", 538=>x"3100", 539=>x"3000", 540=>x"3c00",
---- 541=>x"3600", 542=>x"2e00", 543=>x"2d00", 544=>x"3600",
---- 545=>x"3700", 546=>x"3000", 547=>x"2c00", 548=>x"3500",
---- 549=>x"3700", 550=>x"2d00", 551=>x"2d00", 552=>x"3b00",
---- 553=>x"3900", 554=>x"2e00", 555=>x"4300", 556=>x"3b00",
---- 557=>x"3400", 558=>x"3100", 559=>x"4400", 560=>x"3b00",
---- 561=>x"2e00", 562=>x"2c00", 563=>x"4800", 564=>x"3800",
---- 565=>x"2900", 566=>x"2b00", 567=>x"5000", 568=>x"3200",
---- 569=>x"2900", 570=>x"3000", 571=>x"5f00", 572=>x"2a00",
---- 573=>x"2900", 574=>x"3800", 575=>x"6b00", 576=>x"2d00",
---- 577=>x"2c00", 578=>x"4600", 579=>x"7700", 580=>x"2d00",
---- 581=>x"d100", 582=>x"5900", 583=>x"8300", 584=>x"2c00",
---- 585=>x"3500", 586=>x"6900", 587=>x"8900", 588=>x"2800",
---- 589=>x"4000", 590=>x"7400", 591=>x"8b00", 592=>x"2b00",
---- 593=>x"4b00", 594=>x"7e00", 595=>x"8f00", 596=>x"2e00",
---- 597=>x"5a00", 598=>x"8300", 599=>x"8d00", 600=>x"3800",
---- 601=>x"6c00", 602=>x"8a00", 603=>x"8c00", 604=>x"ba00",
---- 605=>x"7800", 606=>x"8c00", 607=>x"8a00", 608=>x"5600",
---- 609=>x"8300", 610=>x"8c00", 611=>x"8900", 612=>x"6600",
---- 613=>x"8800", 614=>x"8c00", 615=>x"7600", 616=>x"7400",
---- 617=>x"8d00", 618=>x"8c00", 619=>x"8700", 620=>x"7e00",
---- 621=>x"8e00", 622=>x"8900", 623=>x"8900", 624=>x"8700",
---- 625=>x"8d00", 626=>x"8a00", 627=>x"8a00", 628=>x"8d00",
---- 629=>x"8f00", 630=>x"8a00", 631=>x"8c00", 632=>x"9100",
---- 633=>x"9200", 634=>x"8e00", 635=>x"9000", 636=>x"9100",
---- 637=>x"9200", 638=>x"8b00", 639=>x"9400", 640=>x"9200",
---- 641=>x"9000", 642=>x"8d00", 643=>x"9b00", 644=>x"9400",
---- 645=>x"9000", 646=>x"9000", 647=>x"9d00", 648=>x"9500",
---- 649=>x"8f00", 650=>x"9400", 651=>x"9f00", 652=>x"9300",
---- 653=>x"9100", 654=>x"9500", 655=>x"9f00", 656=>x"9200",
---- 657=>x"8e00", 658=>x"9a00", 659=>x"9f00", 660=>x"9200",
---- 661=>x"9200", 662=>x"9c00", 663=>x"9e00", 664=>x"9200",
---- 665=>x"9500", 666=>x"9e00", 667=>x"9c00", 668=>x"9200",
---- 669=>x"9500", 670=>x"9f00", 671=>x"9d00", 672=>x"9200",
---- 673=>x"9900", 674=>x"9f00", 675=>x"9b00", 676=>x"9100",
---- 677=>x"9b00", 678=>x"9e00", 679=>x"9900", 680=>x"9400",
---- 681=>x"9d00", 682=>x"9900", 683=>x"9a00", 684=>x"9700",
---- 685=>x"9c00", 686=>x"9b00", 687=>x"9b00", 688=>x"9500",
---- 689=>x"9c00", 690=>x"9b00", 691=>x"9900", 692=>x"9700",
---- 693=>x"9d00", 694=>x"9b00", 695=>x"9b00", 696=>x"9800",
---- 697=>x"9c00", 698=>x"9a00", 699=>x"9c00", 700=>x"9a00",
---- 701=>x"9b00", 702=>x"9f00", 703=>x"9b00", 704=>x"9a00",
---- 705=>x"9d00", 706=>x"9d00", 707=>x"9a00", 708=>x"9a00",
---- 709=>x"9a00", 710=>x"9a00", 711=>x"9900", 712=>x"9b00",
---- 713=>x"9d00", 714=>x"9c00", 715=>x"9a00", 716=>x"9c00",
---- 717=>x"9e00", 718=>x"9c00", 719=>x"9d00", 720=>x"9b00",
---- 721=>x"9c00", 722=>x"9c00", 723=>x"9c00", 724=>x"9a00",
---- 725=>x"9c00", 726=>x"9a00", 727=>x"9b00", 728=>x"9b00",
---- 729=>x"9900", 730=>x"6600", 731=>x"9b00", 732=>x"9a00",
---- 733=>x"9c00", 734=>x"9800", 735=>x"9d00", 736=>x"9b00",
---- 737=>x"9d00", 738=>x"9a00", 739=>x"9b00", 740=>x"9c00",
---- 741=>x"9c00", 742=>x"9d00", 743=>x"9d00", 744=>x"9e00",
---- 745=>x"9c00", 746=>x"9c00", 747=>x"9d00", 748=>x"9e00",
---- 749=>x"9d00", 750=>x"9900", 751=>x"9c00", 752=>x"9d00",
---- 753=>x"9c00", 754=>x"9b00", 755=>x"9a00", 756=>x"9d00",
---- 757=>x"9d00", 758=>x"9c00", 759=>x"9800", 760=>x"9a00",
---- 761=>x"9d00", 762=>x"9a00", 763=>x"9800", 764=>x"9300",
---- 765=>x"9300", 766=>x"9400", 767=>x"9400", 768=>x"8900",
---- 769=>x"8b00", 770=>x"8c00", 771=>x"8d00", 772=>x"7c00",
---- 773=>x"8200", 774=>x"8300", 775=>x"8600", 776=>x"7300",
---- 777=>x"7a00", 778=>x"7c00", 779=>x"7c00", 780=>x"6f00",
---- 781=>x"6e00", 782=>x"7500", 783=>x"7600", 784=>x"6d00",
---- 785=>x"7000", 786=>x"6f00", 787=>x"7200", 788=>x"7500",
---- 789=>x"7700", 790=>x"7300", 791=>x"7300", 792=>x"8400",
---- 793=>x"7d00", 794=>x"7c00", 795=>x"7a00", 796=>x"8e00",
---- 797=>x"8100", 798=>x"8000", 799=>x"8000", 800=>x"8e00",
---- 801=>x"8a00", 802=>x"8500", 803=>x"8400", 804=>x"8d00",
---- 805=>x"8e00", 806=>x"8700", 807=>x"8600", 808=>x"8e00",
---- 809=>x"8d00", 810=>x"8900", 811=>x"8b00", 812=>x"9100",
---- 813=>x"8e00", 814=>x"8e00", 815=>x"8d00", 816=>x"9200",
---- 817=>x"8f00", 818=>x"8f00", 819=>x"8f00", 820=>x"9100",
---- 821=>x"6f00", 822=>x"9200", 823=>x"8f00", 824=>x"9100",
---- 825=>x"8c00", 826=>x"9000", 827=>x"9100", 828=>x"9000",
---- 829=>x"8d00", 830=>x"7100", 831=>x"8e00", 832=>x"9200",
---- 833=>x"8f00", 834=>x"9000", 835=>x"8c00", 836=>x"9100",
---- 837=>x"8f00", 838=>x"9100", 839=>x"9200", 840=>x"9000",
---- 841=>x"9000", 842=>x"9100", 843=>x"9000", 844=>x"9000",
---- 845=>x"8d00", 846=>x"9300", 847=>x"8e00", 848=>x"9000",
---- 849=>x"8e00", 850=>x"9100", 851=>x"8f00", 852=>x"9000",
---- 853=>x"9100", 854=>x"9100", 855=>x"8f00", 856=>x"9200",
---- 857=>x"9100", 858=>x"9000", 859=>x"9000", 860=>x"9200",
---- 861=>x"9200", 862=>x"8f00", 863=>x"8e00", 864=>x"9300",
---- 865=>x"9100", 866=>x"8f00", 867=>x"8f00", 868=>x"9200",
---- 869=>x"9100", 870=>x"8f00", 871=>x"8e00", 872=>x"9100",
---- 873=>x"9000", 874=>x"8e00", 875=>x"8d00", 876=>x"6f00",
---- 877=>x"8e00", 878=>x"8b00", 879=>x"8c00", 880=>x"8e00",
---- 881=>x"8c00", 882=>x"8d00", 883=>x"8c00", 884=>x"8d00",
---- 885=>x"8b00", 886=>x"8c00", 887=>x"8a00", 888=>x"8d00",
---- 889=>x"8c00", 890=>x"8c00", 891=>x"8900", 892=>x"8e00",
---- 893=>x"8900", 894=>x"8a00", 895=>x"8b00", 896=>x"8e00",
---- 897=>x"8b00", 898=>x"8a00", 899=>x"8c00", 900=>x"9300",
---- 901=>x"8c00", 902=>x"8c00", 903=>x"8d00", 904=>x"8d00",
---- 905=>x"9000", 906=>x"9000", 907=>x"8e00", 908=>x"9200",
---- 909=>x"9300", 910=>x"9100", 911=>x"8f00", 912=>x"9300",
---- 913=>x"9200", 914=>x"9100", 915=>x"9200", 916=>x"8900",
---- 917=>x"8c00", 918=>x"9000", 919=>x"9000", 920=>x"7c00",
---- 921=>x"8000", 922=>x"8400", 923=>x"8a00", 924=>x"6b00",
---- 925=>x"6f00", 926=>x"7400", 927=>x"7b00", 928=>x"5c00",
---- 929=>x"6000", 930=>x"6100", 931=>x"6a00", 932=>x"4f00",
---- 933=>x"5300", 934=>x"5200", 935=>x"5200", 936=>x"4600",
---- 937=>x"4600", 938=>x"4300", 939=>x"4200", 940=>x"5100",
---- 941=>x"4a00", 942=>x"4400", 943=>x"4100", 944=>x"5900",
---- 945=>x"5100", 946=>x"4b00", 947=>x"4400", 948=>x"5c00",
---- 949=>x"5700", 950=>x"5200", 951=>x"4d00", 952=>x"6100",
---- 953=>x"6000", 954=>x"5900", 955=>x"5600", 956=>x"6300",
---- 957=>x"6000", 958=>x"5900", 959=>x"5b00", 960=>x"6500",
---- 961=>x"6200", 962=>x"5d00", 963=>x"5d00", 964=>x"6700",
---- 965=>x"6200", 966=>x"6100", 967=>x"5f00", 968=>x"6900",
---- 969=>x"6100", 970=>x"5f00", 971=>x"6300", 972=>x"6a00",
---- 973=>x"6500", 974=>x"6000", 975=>x"6300", 976=>x"6800",
---- 977=>x"6700", 978=>x"6200", 979=>x"6400", 980=>x"6a00",
---- 981=>x"6900", 982=>x"6500", 983=>x"6800", 984=>x"6800",
---- 985=>x"6b00", 986=>x"6800", 987=>x"6c00", 988=>x"6600",
---- 989=>x"6b00", 990=>x"6b00", 991=>x"6e00", 992=>x"6300",
---- 993=>x"6a00", 994=>x"6d00", 995=>x"9000", 996=>x"6500",
---- 997=>x"6b00", 998=>x"6f00", 999=>x"6e00", 1000=>x"6a00",
---- 1001=>x"6a00", 1002=>x"6d00", 1003=>x"6e00", 1004=>x"5d00",
---- 1005=>x"6700", 1006=>x"6d00", 1007=>x"6900", 1008=>x"6500",
---- 1009=>x"6600", 1010=>x"6400", 1011=>x"6b00", 1012=>x"6000",
---- 1013=>x"6500", 1014=>x"6400", 1015=>x"6800", 1016=>x"5a00",
---- 1017=>x"5b00", 1018=>x"5f00", 1019=>x"6900", 1020=>x"5a00",
---- 1021=>x"5b00", 1022=>x"6000", 1023=>x"6400"),
----
---- 50 => (0=>x"9900", 1=>x"a100", 2=>x"bf00", 3=>x"cc00", 4=>x"9a00",
---- 5=>x"a100", 6=>x"c000", 7=>x"cd00", 8=>x"9800",
---- 9=>x"a000", 10=>x"be00", 11=>x"cc00", 12=>x"9800",
---- 13=>x"9800", 14=>x"ae00", 15=>x"c700", 16=>x"9a00",
---- 17=>x"9600", 18=>x"9c00", 19=>x"ba00", 20=>x"9a00",
---- 21=>x"9800", 22=>x"9500", 23=>x"a700", 24=>x"9a00",
---- 25=>x"9600", 26=>x"9500", 27=>x"9900", 28=>x"9800",
---- 29=>x"9800", 30=>x"9700", 31=>x"9400", 32=>x"9800",
---- 33=>x"9600", 34=>x"9400", 35=>x"9600", 36=>x"9700",
---- 37=>x"9800", 38=>x"9700", 39=>x"9400", 40=>x"9600",
---- 41=>x"9700", 42=>x"9800", 43=>x"9600", 44=>x"9800",
---- 45=>x"9500", 46=>x"9600", 47=>x"9500", 48=>x"9800",
---- 49=>x"9500", 50=>x"9600", 51=>x"9600", 52=>x"9800",
---- 53=>x"9700", 54=>x"9600", 55=>x"9700", 56=>x"9800",
---- 57=>x"9700", 58=>x"9800", 59=>x"9700", 60=>x"9800",
---- 61=>x"9900", 62=>x"9600", 63=>x"9600", 64=>x"9a00",
---- 65=>x"9b00", 66=>x"9800", 67=>x"9800", 68=>x"9b00",
---- 69=>x"9900", 70=>x"9800", 71=>x"9900", 72=>x"9c00",
---- 73=>x"9900", 74=>x"9700", 75=>x"9800", 76=>x"9b00",
---- 77=>x"9900", 78=>x"9500", 79=>x"9400", 80=>x"9700",
---- 81=>x"9900", 82=>x"9600", 83=>x"9400", 84=>x"6800",
---- 85=>x"9300", 86=>x"9500", 87=>x"9400", 88=>x"9500",
---- 89=>x"9400", 90=>x"9000", 91=>x"8f00", 92=>x"9300",
---- 93=>x"9500", 94=>x"9200", 95=>x"8f00", 96=>x"9300",
---- 97=>x"9100", 98=>x"9300", 99=>x"9000", 100=>x"9200",
---- 101=>x"8f00", 102=>x"8e00", 103=>x"8d00", 104=>x"9200",
---- 105=>x"8c00", 106=>x"8c00", 107=>x"8e00", 108=>x"9300",
---- 109=>x"9100", 110=>x"8c00", 111=>x"7200", 112=>x"9000",
---- 113=>x"8d00", 114=>x"8e00", 115=>x"8b00", 116=>x"8f00",
---- 117=>x"8e00", 118=>x"8d00", 119=>x"8e00", 120=>x"8e00",
---- 121=>x"8f00", 122=>x"8d00", 123=>x"8d00", 124=>x"9000",
---- 125=>x"8e00", 126=>x"9000", 127=>x"8e00", 128=>x"9000",
---- 129=>x"8f00", 130=>x"9100", 131=>x"8f00", 132=>x"8d00",
---- 133=>x"8f00", 134=>x"8e00", 135=>x"8d00", 136=>x"8e00",
---- 137=>x"9000", 138=>x"8e00", 139=>x"9000", 140=>x"8e00",
---- 141=>x"8e00", 142=>x"8e00", 143=>x"8e00", 144=>x"8f00",
---- 145=>x"8f00", 146=>x"8f00", 147=>x"8c00", 148=>x"8c00",
---- 149=>x"9100", 150=>x"8d00", 151=>x"8c00", 152=>x"8d00",
---- 153=>x"8e00", 154=>x"8f00", 155=>x"8f00", 156=>x"8f00",
---- 157=>x"9100", 158=>x"8f00", 159=>x"8f00", 160=>x"8f00",
---- 161=>x"8f00", 162=>x"8f00", 163=>x"9000", 164=>x"8c00",
---- 165=>x"8f00", 166=>x"9000", 167=>x"8f00", 168=>x"8e00",
---- 169=>x"8f00", 170=>x"9000", 171=>x"8e00", 172=>x"8e00",
---- 173=>x"8e00", 174=>x"9200", 175=>x"9200", 176=>x"9000",
---- 177=>x"8e00", 178=>x"9000", 179=>x"9000", 180=>x"9100",
---- 181=>x"8e00", 182=>x"8e00", 183=>x"8e00", 184=>x"8f00",
---- 185=>x"8f00", 186=>x"9000", 187=>x"8e00", 188=>x"8c00",
---- 189=>x"8e00", 190=>x"8e00", 191=>x"9000", 192=>x"8e00",
---- 193=>x"8e00", 194=>x"8d00", 195=>x"8d00", 196=>x"8f00",
---- 197=>x"8f00", 198=>x"8d00", 199=>x"8d00", 200=>x"9000",
---- 201=>x"8e00", 202=>x"8b00", 203=>x"8e00", 204=>x"9100",
---- 205=>x"8d00", 206=>x"8c00", 207=>x"8d00", 208=>x"9000",
---- 209=>x"8c00", 210=>x"8c00", 211=>x"8b00", 212=>x"6c00",
---- 213=>x"8e00", 214=>x"8c00", 215=>x"8a00", 216=>x"8f00",
---- 217=>x"8700", 218=>x"8700", 219=>x"8a00", 220=>x"9f00",
---- 221=>x"a300", 222=>x"9b00", 223=>x"8600", 224=>x"d700",
---- 225=>x"da00", 226=>x"ce00", 227=>x"a800", 228=>x"d200",
---- 229=>x"c900", 230=>x"c800", 231=>x"cd00", 232=>x"bd00",
---- 233=>x"c600", 234=>x"cf00", 235=>x"d800", 236=>x"d000",
---- 237=>x"da00", 238=>x"df00", 239=>x"e200", 240=>x"db00",
---- 241=>x"e100", 242=>x"e200", 243=>x"df00", 244=>x"da00",
---- 245=>x"db00", 246=>x"da00", 247=>x"d900", 248=>x"d600",
---- 249=>x"d500", 250=>x"d700", 251=>x"d700", 252=>x"d200",
---- 253=>x"d300", 254=>x"d500", 255=>x"ce00", 256=>x"c800",
---- 257=>x"cb00", 258=>x"ce00", 259=>x"cb00", 260=>x"c600",
---- 261=>x"ca00", 262=>x"ca00", 263=>x"3100", 264=>x"ca00",
---- 265=>x"cc00", 266=>x"cd00", 267=>x"d300", 268=>x"cb00",
---- 269=>x"cc00", 270=>x"cf00", 271=>x"d300", 272=>x"cb00",
---- 273=>x"cf00", 274=>x"d300", 275=>x"d500", 276=>x"ce00",
---- 277=>x"d200", 278=>x"d500", 279=>x"d700", 280=>x"cd00",
---- 281=>x"d200", 282=>x"d500", 283=>x"d500", 284=>x"cb00",
---- 285=>x"ce00", 286=>x"d200", 287=>x"d500", 288=>x"c700",
---- 289=>x"ce00", 290=>x"d100", 291=>x"d400", 292=>x"c700",
---- 293=>x"d300", 294=>x"d300", 295=>x"d400", 296=>x"c900",
---- 297=>x"d000", 298=>x"d100", 299=>x"d300", 300=>x"c800",
---- 301=>x"cd00", 302=>x"d200", 303=>x"d200", 304=>x"be00",
---- 305=>x"ca00", 306=>x"d000", 307=>x"cd00", 308=>x"bc00",
---- 309=>x"cc00", 310=>x"c100", 311=>x"c400", 312=>x"be00",
---- 313=>x"a400", 314=>x"a800", 315=>x"be00", 316=>x"9600",
---- 317=>x"7b00", 318=>x"a700", 319=>x"bd00", 320=>x"7a00",
---- 321=>x"9600", 322=>x"ad00", 323=>x"ba00", 324=>x"9100",
---- 325=>x"a600", 326=>x"b000", 327=>x"b600", 328=>x"a900",
---- 329=>x"a600", 330=>x"a900", 331=>x"c600", 332=>x"9b00",
---- 333=>x"9000", 334=>x"ad00", 335=>x"df00", 336=>x"7d00",
---- 337=>x"9d00", 338=>x"c300", 339=>x"e500", 340=>x"8200",
---- 341=>x"b100", 342=>x"d900", 343=>x"d600", 344=>x"9f00",
---- 345=>x"c700", 346=>x"e700", 347=>x"a900", 348=>x"c400",
---- 349=>x"d900", 350=>x"e000", 351=>x"6300", 352=>x"2d00",
---- 353=>x"e300", 354=>x"a300", 355=>x"2600", 356=>x"d700",
---- 357=>x"cb00", 358=>x"4300", 359=>x"2100", 360=>x"e300",
---- 361=>x"7f00", 362=>x"2a00", 363=>x"2a00", 364=>x"a100",
---- 365=>x"3000", 366=>x"3300", 367=>x"2b00", 368=>x"3300",
---- 369=>x"2300", 370=>x"2800", 371=>x"2a00", 372=>x"2900",
---- 373=>x"d500", 374=>x"2d00", 375=>x"3000", 376=>x"2e00",
---- 377=>x"2e00", 378=>x"2d00", 379=>x"3300", 380=>x"3000",
---- 381=>x"2f00", 382=>x"3400", 383=>x"3600", 384=>x"2f00",
---- 385=>x"3400", 386=>x"3800", 387=>x"3500", 388=>x"3700",
---- 389=>x"3b00", 390=>x"3800", 391=>x"3400", 392=>x"3500",
---- 393=>x"3700", 394=>x"3600", 395=>x"3300", 396=>x"3500",
---- 397=>x"3400", 398=>x"3600", 399=>x"3400", 400=>x"3500",
---- 401=>x"3700", 402=>x"3500", 403=>x"3700", 404=>x"3800",
---- 405=>x"3900", 406=>x"3f00", 407=>x"3600", 408=>x"3800",
---- 409=>x"3b00", 410=>x"3700", 411=>x"2f00", 412=>x"3700",
---- 413=>x"3800", 414=>x"3700", 415=>x"3100", 416=>x"3600",
---- 417=>x"3700", 418=>x"3500", 419=>x"d000", 420=>x"3700",
---- 421=>x"3a00", 422=>x"3300", 423=>x"2a00", 424=>x"3800",
---- 425=>x"3500", 426=>x"3000", 427=>x"2900", 428=>x"3900",
---- 429=>x"3000", 430=>x"3000", 431=>x"2c00", 432=>x"3600",
---- 433=>x"2f00", 434=>x"3500", 435=>x"2d00", 436=>x"3700",
---- 437=>x"2f00", 438=>x"2d00", 439=>x"2e00", 440=>x"3200",
---- 441=>x"3000", 442=>x"2e00", 443=>x"2a00", 444=>x"2e00",
---- 445=>x"2c00", 446=>x"2d00", 447=>x"2d00", 448=>x"2f00",
---- 449=>x"2d00", 450=>x"2d00", 451=>x"2f00", 452=>x"2e00",
---- 453=>x"2c00", 454=>x"3000", 455=>x"3300", 456=>x"2e00",
---- 457=>x"d300", 458=>x"3000", 459=>x"3300", 460=>x"2f00",
---- 461=>x"2e00", 462=>x"2e00", 463=>x"3300", 464=>x"2e00",
---- 465=>x"3300", 466=>x"3200", 467=>x"3600", 468=>x"2d00",
---- 469=>x"2e00", 470=>x"3700", 471=>x"3700", 472=>x"3300",
---- 473=>x"3300", 474=>x"3800", 475=>x"3300", 476=>x"3300",
---- 477=>x"3600", 478=>x"3600", 479=>x"3200", 480=>x"3000",
---- 481=>x"3400", 482=>x"3500", 483=>x"2e00", 484=>x"3300",
---- 485=>x"3900", 486=>x"3400", 487=>x"2c00", 488=>x"3400",
---- 489=>x"3800", 490=>x"3100", 491=>x"2d00", 492=>x"3400",
---- 493=>x"3600", 494=>x"2f00", 495=>x"2d00", 496=>x"3900",
---- 497=>x"3400", 498=>x"3000", 499=>x"2c00", 500=>x"3900",
---- 501=>x"3800", 502=>x"3300", 503=>x"3000", 504=>x"3800",
---- 505=>x"3a00", 506=>x"3700", 507=>x"3600", 508=>x"3600",
---- 509=>x"3100", 510=>x"3700", 511=>x"4400", 512=>x"3400",
---- 513=>x"2b00", 514=>x"3200", 515=>x"5000", 516=>x"3400",
---- 517=>x"2800", 518=>x"2c00", 519=>x"5a00", 520=>x"3400",
---- 521=>x"2700", 522=>x"2e00", 523=>x"6500", 524=>x"3100",
---- 525=>x"2c00", 526=>x"4200", 527=>x"7700", 528=>x"2d00",
---- 529=>x"3100", 530=>x"5900", 531=>x"8300", 532=>x"cd00",
---- 533=>x"4000", 534=>x"6900", 535=>x"8c00", 536=>x"3300",
---- 537=>x"4800", 538=>x"7800", 539=>x"8e00", 540=>x"2e00",
---- 541=>x"5400", 542=>x"8400", 543=>x"9100", 544=>x"3200",
---- 545=>x"6400", 546=>x"8800", 547=>x"8d00", 548=>x"4100",
---- 549=>x"7100", 550=>x"8c00", 551=>x"8b00", 552=>x"5f00",
---- 553=>x"7900", 554=>x"8d00", 555=>x"8800", 556=>x"6a00",
---- 557=>x"8500", 558=>x"8a00", 559=>x"8500", 560=>x"7900",
---- 561=>x"8b00", 562=>x"8800", 563=>x"8300", 564=>x"8100",
---- 565=>x"8900", 566=>x"8500", 567=>x"8100", 568=>x"8700",
---- 569=>x"8b00", 570=>x"8500", 571=>x"8500", 572=>x"8700",
---- 573=>x"8700", 574=>x"7b00", 575=>x"8800", 576=>x"8b00",
---- 577=>x"8800", 578=>x"8400", 579=>x"8b00", 580=>x"8d00",
---- 581=>x"8600", 582=>x"8400", 583=>x"9300", 584=>x"8b00",
---- 585=>x"8500", 586=>x"8600", 587=>x"9900", 588=>x"8b00",
---- 589=>x"8600", 590=>x"8a00", 591=>x"9b00", 592=>x"8c00",
---- 593=>x"8800", 594=>x"9200", 595=>x"9f00", 596=>x"8900",
---- 597=>x"8900", 598=>x"9800", 599=>x"a200", 600=>x"8900",
---- 601=>x"9000", 602=>x"a300", 603=>x"a700", 604=>x"8500",
---- 605=>x"9200", 606=>x"ae00", 607=>x"ac00", 608=>x"8800",
---- 609=>x"9a00", 610=>x"a000", 611=>x"a200", 612=>x"8c00",
---- 613=>x"9e00", 614=>x"a200", 615=>x"a000", 616=>x"9100",
---- 617=>x"a000", 618=>x"a000", 619=>x"9e00", 620=>x"9700",
---- 621=>x"a000", 622=>x"9f00", 623=>x"9f00", 624=>x"9b00",
---- 625=>x"a000", 626=>x"9d00", 627=>x"9d00", 628=>x"9e00",
---- 629=>x"a100", 630=>x"9c00", 631=>x"9d00", 632=>x"a000",
---- 633=>x"9f00", 634=>x"9c00", 635=>x"9a00", 636=>x"a100",
---- 637=>x"9d00", 638=>x"9c00", 639=>x"9c00", 640=>x"a000",
---- 641=>x"9e00", 642=>x"9c00", 643=>x"9a00", 644=>x"a000",
---- 645=>x"9d00", 646=>x"9c00", 647=>x"9a00", 648=>x"9d00",
---- 649=>x"9d00", 650=>x"9900", 651=>x"9900", 652=>x"9d00",
---- 653=>x"9d00", 654=>x"9b00", 655=>x"9900", 656=>x"9e00",
---- 657=>x"9b00", 658=>x"9900", 659=>x"9b00", 660=>x"9b00",
---- 661=>x"9b00", 662=>x"9b00", 663=>x"9a00", 664=>x"9a00",
---- 665=>x"9900", 666=>x"9a00", 667=>x"9a00", 668=>x"9c00",
---- 669=>x"9b00", 670=>x"6500", 671=>x"6600", 672=>x"9900",
---- 673=>x"9900", 674=>x"9900", 675=>x"9800", 676=>x"9a00",
---- 677=>x"9b00", 678=>x"9700", 679=>x"9800", 680=>x"9a00",
---- 681=>x"9a00", 682=>x"9800", 683=>x"9800", 684=>x"9b00",
---- 685=>x"9a00", 686=>x"9800", 687=>x"9800", 688=>x"9b00",
---- 689=>x"9900", 690=>x"9800", 691=>x"9700", 692=>x"9a00",
---- 693=>x"9900", 694=>x"9500", 695=>x"9700", 696=>x"9900",
---- 697=>x"9600", 698=>x"9800", 699=>x"9500", 700=>x"9600",
---- 701=>x"9800", 702=>x"9900", 703=>x"9800", 704=>x"9900",
---- 705=>x"9800", 706=>x"9700", 707=>x"9700", 708=>x"9700",
---- 709=>x"9800", 710=>x"9a00", 711=>x"9700", 712=>x"9600",
---- 713=>x"9800", 714=>x"9a00", 715=>x"9700", 716=>x"9b00",
---- 717=>x"9c00", 718=>x"9900", 719=>x"9800", 720=>x"9900",
---- 721=>x"9a00", 722=>x"9a00", 723=>x"9900", 724=>x"9900",
---- 725=>x"9700", 726=>x"9a00", 727=>x"9a00", 728=>x"9900",
---- 729=>x"9900", 730=>x"9b00", 731=>x"9900", 732=>x"9a00",
---- 733=>x"9b00", 734=>x"9b00", 735=>x"9800", 736=>x"9a00",
---- 737=>x"6600", 738=>x"9b00", 739=>x"9a00", 740=>x"9900",
---- 741=>x"9700", 742=>x"9c00", 743=>x"9800", 744=>x"9a00",
---- 745=>x"9800", 746=>x"9c00", 747=>x"9700", 748=>x"9a00",
---- 749=>x"9a00", 750=>x"9a00", 751=>x"9700", 752=>x"9500",
---- 753=>x"9800", 754=>x"9700", 755=>x"9600", 756=>x"9500",
---- 757=>x"9600", 758=>x"9800", 759=>x"9700", 760=>x"9200",
---- 761=>x"9500", 762=>x"9800", 763=>x"9800", 764=>x"9500",
---- 765=>x"9800", 766=>x"9400", 767=>x"9600", 768=>x"9200",
---- 769=>x"9300", 770=>x"9200", 771=>x"9600", 772=>x"8900",
---- 773=>x"8b00", 774=>x"8b00", 775=>x"8c00", 776=>x"7b00",
---- 777=>x"8400", 778=>x"8100", 779=>x"8100", 780=>x"7500",
---- 781=>x"7a00", 782=>x"7500", 783=>x"7a00", 784=>x"7200",
---- 785=>x"7100", 786=>x"7200", 787=>x"7400", 788=>x"7100",
---- 789=>x"6e00", 790=>x"7000", 791=>x"6f00", 792=>x"7500",
---- 793=>x"7100", 794=>x"6f00", 795=>x"6c00", 796=>x"7a00",
---- 797=>x"7b00", 798=>x"7700", 799=>x"7100", 800=>x"7c00",
---- 801=>x"8000", 802=>x"7f00", 803=>x"8500", 804=>x"8600",
---- 805=>x"8600", 806=>x"8200", 807=>x"8300", 808=>x"8800",
---- 809=>x"8900", 810=>x"8900", 811=>x"8900", 812=>x"8b00",
---- 813=>x"8a00", 814=>x"8a00", 815=>x"8700", 816=>x"8e00",
---- 817=>x"8e00", 818=>x"8c00", 819=>x"8800", 820=>x"9000",
---- 821=>x"8f00", 822=>x"8c00", 823=>x"8b00", 824=>x"8e00",
---- 825=>x"8d00", 826=>x"8e00", 827=>x"8d00", 828=>x"8f00",
---- 829=>x"8f00", 830=>x"8e00", 831=>x"8d00", 832=>x"8c00",
---- 833=>x"8e00", 834=>x"8d00", 835=>x"8d00", 836=>x"8f00",
---- 837=>x"9000", 838=>x"8f00", 839=>x"8f00", 840=>x"8d00",
---- 841=>x"8f00", 842=>x"8d00", 843=>x"8c00", 844=>x"8a00",
---- 845=>x"8c00", 846=>x"8d00", 847=>x"8a00", 848=>x"8b00",
---- 849=>x"8b00", 850=>x"8d00", 851=>x"8d00", 852=>x"8e00",
---- 853=>x"8d00", 854=>x"8d00", 855=>x"8b00", 856=>x"8f00",
---- 857=>x"8f00", 858=>x"8a00", 859=>x"8b00", 860=>x"8e00",
---- 861=>x"8d00", 862=>x"8b00", 863=>x"8a00", 864=>x"8b00",
---- 865=>x"8c00", 866=>x"8c00", 867=>x"8800", 868=>x"8a00",
---- 869=>x"8b00", 870=>x"8c00", 871=>x"8a00", 872=>x"8c00",
---- 873=>x"8d00", 874=>x"8900", 875=>x"8b00", 876=>x"8a00",
---- 877=>x"8d00", 878=>x"8d00", 879=>x"8900", 880=>x"8a00",
---- 881=>x"8c00", 882=>x"8d00", 883=>x"8a00", 884=>x"8b00",
---- 885=>x"8c00", 886=>x"8a00", 887=>x"8a00", 888=>x"8b00",
---- 889=>x"8e00", 890=>x"8b00", 891=>x"8c00", 892=>x"8a00",
---- 893=>x"8b00", 894=>x"8c00", 895=>x"8b00", 896=>x"8a00",
---- 897=>x"8b00", 898=>x"8d00", 899=>x"8a00", 900=>x"8c00",
---- 901=>x"8c00", 902=>x"8f00", 903=>x"8b00", 904=>x"8d00",
---- 905=>x"8f00", 906=>x"8d00", 907=>x"8b00", 908=>x"8e00",
---- 909=>x"8e00", 910=>x"8f00", 911=>x"8d00", 912=>x"8f00",
---- 913=>x"9000", 914=>x"8f00", 915=>x"9000", 916=>x"9100",
---- 917=>x"9200", 918=>x"9000", 919=>x"8f00", 920=>x"8b00",
---- 921=>x"8e00", 922=>x"8e00", 923=>x"8b00", 924=>x"7b00",
---- 925=>x"8000", 926=>x"8600", 927=>x"8500", 928=>x"6800",
---- 929=>x"6b00", 930=>x"7400", 931=>x"7600", 932=>x"5500",
---- 933=>x"5900", 934=>x"5d00", 935=>x"6200", 936=>x"4700",
---- 937=>x"4800", 938=>x"4a00", 939=>x"4900", 940=>x"3e00",
---- 941=>x"3900", 942=>x"3800", 943=>x"3700", 944=>x"3f00",
---- 945=>x"3900", 946=>x"3500", 947=>x"3100", 948=>x"b500",
---- 949=>x"3e00", 950=>x"3700", 951=>x"3300", 952=>x"5000",
---- 953=>x"4700", 954=>x"3f00", 955=>x"3600", 956=>x"5400",
---- 957=>x"4d00", 958=>x"4900", 959=>x"4100", 960=>x"5500",
---- 961=>x"5100", 962=>x"5200", 963=>x"4600", 964=>x"5b00",
---- 965=>x"5800", 966=>x"5200", 967=>x"4b00", 968=>x"5f00",
---- 969=>x"5e00", 970=>x"5500", 971=>x"4f00", 972=>x"9e00",
---- 973=>x"6200", 974=>x"5c00", 975=>x"5500", 976=>x"6200",
---- 977=>x"6600", 978=>x"5f00", 979=>x"5900", 980=>x"6700",
---- 981=>x"6500", 982=>x"6100", 983=>x"6000", 984=>x"6800",
---- 985=>x"6400", 986=>x"6400", 987=>x"6400", 988=>x"6d00",
---- 989=>x"6700", 990=>x"6700", 991=>x"6900", 992=>x"6e00",
---- 993=>x"6b00", 994=>x"6a00", 995=>x"7000", 996=>x"6d00",
---- 997=>x"7100", 998=>x"7300", 999=>x"7500", 1000=>x"6f00",
---- 1001=>x"7300", 1002=>x"7900", 1003=>x"7800", 1004=>x"6e00",
---- 1005=>x"7500", 1006=>x"7800", 1007=>x"7800", 1008=>x"7000",
---- 1009=>x"7500", 1010=>x"7600", 1011=>x"7800", 1012=>x"6e00",
---- 1013=>x"7300", 1014=>x"7600", 1015=>x"7500", 1016=>x"6d00",
---- 1017=>x"7200", 1018=>x"7100", 1019=>x"7300", 1020=>x"6900",
---- 1021=>x"6700", 1022=>x"7400", 1023=>x"7d00"),
----
---- 51 => (0=>x"d400", 1=>x"d500", 2=>x"da00", 3=>x"da00", 4=>x"d300",
---- 5=>x"d500", 6=>x"2500", 7=>x"da00", 8=>x"d200",
---- 9=>x"d600", 10=>x"d900", 11=>x"da00", 12=>x"d000",
---- 13=>x"d600", 14=>x"d800", 15=>x"da00", 16=>x"cc00",
---- 17=>x"d300", 18=>x"d500", 19=>x"d900", 20=>x"c300",
---- 21=>x"cf00", 22=>x"d600", 23=>x"d700", 24=>x"b400",
---- 25=>x"c800", 26=>x"d200", 27=>x"d600", 28=>x"a100",
---- 29=>x"c100", 30=>x"cc00", 31=>x"d400", 32=>x"9600",
---- 33=>x"b200", 34=>x"c900", 35=>x"d200", 36=>x"9200",
---- 37=>x"9c00", 38=>x"bb00", 39=>x"ce00", 40=>x"9600",
---- 41=>x"9200", 42=>x"a800", 43=>x"c500", 44=>x"9200",
---- 45=>x"7100", 46=>x"9800", 47=>x"b700", 48=>x"9500",
---- 49=>x"9100", 50=>x"9100", 51=>x"a500", 52=>x"9400",
---- 53=>x"9300", 54=>x"9100", 55=>x"9600", 56=>x"9400",
---- 57=>x"9300", 58=>x"9200", 59=>x"9000", 60=>x"9500",
---- 61=>x"9200", 62=>x"9100", 63=>x"9000", 64=>x"9600",
---- 65=>x"9500", 66=>x"9400", 67=>x"8d00", 68=>x"9800",
---- 69=>x"9400", 70=>x"9400", 71=>x"8f00", 72=>x"9700",
---- 73=>x"9500", 74=>x"9500", 75=>x"9100", 76=>x"9700",
---- 77=>x"9400", 78=>x"9400", 79=>x"9100", 80=>x"9500",
---- 81=>x"9400", 82=>x"9100", 83=>x"6d00", 84=>x"9200",
---- 85=>x"9200", 86=>x"9100", 87=>x"8f00", 88=>x"9000",
---- 89=>x"9000", 90=>x"8f00", 91=>x"9000", 92=>x"9100",
---- 93=>x"9000", 94=>x"8f00", 95=>x"8f00", 96=>x"9200",
---- 97=>x"9000", 98=>x"8e00", 99=>x"8e00", 100=>x"8f00",
---- 101=>x"8f00", 102=>x"8b00", 103=>x"8e00", 104=>x"8d00",
---- 105=>x"8d00", 106=>x"8c00", 107=>x"8e00", 108=>x"8e00",
---- 109=>x"8b00", 110=>x"7200", 111=>x"8c00", 112=>x"8c00",
---- 113=>x"8c00", 114=>x"8a00", 115=>x"8d00", 116=>x"8b00",
---- 117=>x"8d00", 118=>x"8a00", 119=>x"8a00", 120=>x"8d00",
---- 121=>x"8b00", 122=>x"8d00", 123=>x"8d00", 124=>x"8d00",
---- 125=>x"8d00", 126=>x"8d00", 127=>x"8e00", 128=>x"8d00",
---- 129=>x"8b00", 130=>x"8d00", 131=>x"8e00", 132=>x"8e00",
---- 133=>x"8c00", 134=>x"8e00", 135=>x"8e00", 136=>x"8d00",
---- 137=>x"8d00", 138=>x"8c00", 139=>x"8f00", 140=>x"8e00",
---- 141=>x"8d00", 142=>x"8f00", 143=>x"8f00", 144=>x"8e00",
---- 145=>x"8f00", 146=>x"9000", 147=>x"9000", 148=>x"9000",
---- 149=>x"8e00", 150=>x"9000", 151=>x"9100", 152=>x"8f00",
---- 153=>x"9000", 154=>x"9100", 155=>x"9100", 156=>x"8f00",
---- 157=>x"8f00", 158=>x"9000", 159=>x"9000", 160=>x"9000",
---- 161=>x"9200", 162=>x"9000", 163=>x"9100", 164=>x"9000",
---- 165=>x"9100", 166=>x"9100", 167=>x"9200", 168=>x"8e00",
---- 169=>x"8f00", 170=>x"9200", 171=>x"9300", 172=>x"8e00",
---- 173=>x"8f00", 174=>x"9100", 175=>x"9000", 176=>x"9000",
---- 177=>x"8f00", 178=>x"8f00", 179=>x"9100", 180=>x"9100",
---- 181=>x"9100", 182=>x"9100", 183=>x"6c00", 184=>x"8f00",
---- 185=>x"8f00", 186=>x"9200", 187=>x"9000", 188=>x"9100",
---- 189=>x"9000", 190=>x"8f00", 191=>x"9000", 192=>x"8f00",
---- 193=>x"9100", 194=>x"9000", 195=>x"9200", 196=>x"8d00",
---- 197=>x"9000", 198=>x"6e00", 199=>x"9100", 200=>x"8f00",
---- 201=>x"8f00", 202=>x"9100", 203=>x"9200", 204=>x"8f00",
---- 205=>x"8e00", 206=>x"9400", 207=>x"9400", 208=>x"8b00",
---- 209=>x"6f00", 210=>x"9200", 211=>x"9300", 212=>x"8c00",
---- 213=>x"9000", 214=>x"9300", 215=>x"6900", 216=>x"8e00",
---- 217=>x"8f00", 218=>x"9300", 219=>x"9500", 220=>x"8900",
---- 221=>x"9300", 222=>x"9700", 223=>x"9500", 224=>x"a500",
---- 225=>x"c200", 226=>x"ae00", 227=>x"8e00", 228=>x"d500",
---- 229=>x"d900", 230=>x"d700", 231=>x"ac00", 232=>x"da00",
---- 233=>x"da00", 234=>x"dc00", 235=>x"d400", 236=>x"e500",
---- 237=>x"e900", 238=>x"df00", 239=>x"e300", 240=>x"e000",
---- 241=>x"e400", 242=>x"e800", 243=>x"ed00", 244=>x"de00",
---- 245=>x"de00", 246=>x"e200", 247=>x"eb00", 248=>x"d300",
---- 249=>x"d600", 250=>x"df00", 251=>x"e800", 252=>x"c900",
---- 253=>x"d200", 254=>x"dc00", 255=>x"e600", 256=>x"d100",
---- 257=>x"d700", 258=>x"dc00", 259=>x"e200", 260=>x"d400",
---- 261=>x"db00", 262=>x"de00", 263=>x"e300", 264=>x"d700",
---- 265=>x"d900", 266=>x"dd00", 267=>x"e100", 268=>x"d900",
---- 269=>x"dc00", 270=>x"de00", 271=>x"e000", 272=>x"2700",
---- 273=>x"da00", 274=>x"de00", 275=>x"e100", 276=>x"d800",
---- 277=>x"db00", 278=>x"dd00", 279=>x"e200", 280=>x"da00",
---- 281=>x"de00", 282=>x"dc00", 283=>x"e500", 284=>x"db00",
---- 285=>x"dd00", 286=>x"dc00", 287=>x"e600", 288=>x"da00",
---- 289=>x"de00", 290=>x"dd00", 291=>x"e600", 292=>x"db00",
---- 293=>x"de00", 294=>x"e000", 295=>x"e000", 296=>x"db00",
---- 297=>x"de00", 298=>x"e100", 299=>x"ca00", 300=>x"d800",
---- 301=>x"d800", 302=>x"df00", 303=>x"a400", 304=>x"d700",
---- 305=>x"d800", 306=>x"dc00", 307=>x"7500", 308=>x"d300",
---- 309=>x"d700", 310=>x"c900", 311=>x"4100", 312=>x"cb00",
---- 313=>x"db00", 314=>x"9700", 315=>x"2400", 316=>x"c600",
---- 317=>x"d500", 318=>x"5900", 319=>x"2500", 320=>x"d300",
---- 321=>x"b600", 322=>x"2d00", 323=>x"2600", 324=>x"de00",
---- 325=>x"8f00", 326=>x"1d00", 327=>x"2900", 328=>x"dc00",
---- 329=>x"5600", 330=>x"2000", 331=>x"2d00", 332=>x"b900",
---- 333=>x"3000", 334=>x"2600", 335=>x"2c00", 336=>x"7d00",
---- 337=>x"1d00", 338=>x"2900", 339=>x"2a00", 340=>x"4b00",
---- 341=>x"1f00", 342=>x"d900", 343=>x"2c00", 344=>x"2500",
---- 345=>x"2200", 346=>x"2300", 347=>x"2a00", 348=>x"1c00",
---- 349=>x"2700", 350=>x"2600", 351=>x"2b00", 352=>x"2300",
---- 353=>x"2c00", 354=>x"2e00", 355=>x"2e00", 356=>x"2700",
---- 357=>x"d500", 358=>x"3200", 359=>x"3100", 360=>x"2a00",
---- 361=>x"2f00", 362=>x"3000", 363=>x"3300", 364=>x"2b00",
---- 365=>x"3100", 366=>x"3400", 367=>x"3200", 368=>x"3100",
---- 369=>x"3400", 370=>x"3300", 371=>x"3000", 372=>x"3400",
---- 373=>x"3200", 374=>x"3000", 375=>x"2c00", 376=>x"3300",
---- 377=>x"3500", 378=>x"2f00", 379=>x"2e00", 380=>x"3700",
---- 381=>x"3500", 382=>x"2e00", 383=>x"2c00", 384=>x"3600",
---- 385=>x"3800", 386=>x"2f00", 387=>x"2f00", 388=>x"3200",
---- 389=>x"3000", 390=>x"3100", 391=>x"3200", 392=>x"c700",
---- 393=>x"3100", 394=>x"2d00", 395=>x"2d00", 396=>x"3700",
---- 397=>x"3100", 398=>x"2c00", 399=>x"2f00", 400=>x"3500",
---- 401=>x"3100", 402=>x"2e00", 403=>x"2e00", 404=>x"3300",
---- 405=>x"3200", 406=>x"2e00", 407=>x"2c00", 408=>x"2c00",
---- 409=>x"3000", 410=>x"2c00", 411=>x"2c00", 412=>x"2e00",
---- 413=>x"2e00", 414=>x"2f00", 415=>x"2e00", 416=>x"2b00",
---- 417=>x"2f00", 418=>x"2d00", 419=>x"3100", 420=>x"2900",
---- 421=>x"2f00", 422=>x"3000", 423=>x"3400", 424=>x"2900",
---- 425=>x"3000", 426=>x"3600", 427=>x"3700", 428=>x"2900",
---- 429=>x"2c00", 430=>x"3200", 431=>x"3500", 432=>x"2900",
---- 433=>x"2c00", 434=>x"3300", 435=>x"3300", 436=>x"2d00",
---- 437=>x"3300", 438=>x"3400", 439=>x"d300", 440=>x"2e00",
---- 441=>x"3400", 442=>x"3100", 443=>x"2f00", 444=>x"2e00",
---- 445=>x"3600", 446=>x"2e00", 447=>x"3000", 448=>x"3400",
---- 449=>x"3600", 450=>x"2b00", 451=>x"2c00", 452=>x"3800",
---- 453=>x"3700", 454=>x"2d00", 455=>x"2a00", 456=>x"3700",
---- 457=>x"3300", 458=>x"2a00", 459=>x"2d00", 460=>x"3500",
---- 461=>x"2e00", 462=>x"2b00", 463=>x"3a00", 464=>x"3900",
---- 465=>x"2e00", 466=>x"2a00", 467=>x"4700", 468=>x"3000",
---- 469=>x"2b00", 470=>x"2d00", 471=>x"5600", 472=>x"2a00",
---- 473=>x"2c00", 474=>x"4300", 475=>x"6e00", 476=>x"2a00",
---- 477=>x"3100", 478=>x"5700", 479=>x"7e00", 480=>x"2b00",
---- 481=>x"3600", 482=>x"6300", 483=>x"8600", 484=>x"3100",
---- 485=>x"4b00", 486=>x"7000", 487=>x"8900", 488=>x"3400",
---- 489=>x"5800", 490=>x"7f00", 491=>x"8b00", 492=>x"c200",
---- 493=>x"6400", 494=>x"8500", 495=>x"8d00", 496=>x"4500",
---- 497=>x"7000", 498=>x"8900", 499=>x"8a00", 500=>x"4e00",
---- 501=>x"7f00", 502=>x"8e00", 503=>x"8600", 504=>x"5b00",
---- 505=>x"8400", 506=>x"8d00", 507=>x"8400", 508=>x"6c00",
---- 509=>x"8900", 510=>x"8b00", 511=>x"8200", 512=>x"7d00",
---- 513=>x"8d00", 514=>x"8900", 515=>x"7f00", 516=>x"8700",
---- 517=>x"8d00", 518=>x"8600", 519=>x"8100", 520=>x"8e00",
---- 521=>x"8c00", 522=>x"8500", 523=>x"8600", 524=>x"8e00",
---- 525=>x"8d00", 526=>x"8700", 527=>x"8b00", 528=>x"9100",
---- 529=>x"8e00", 530=>x"8700", 531=>x"9100", 532=>x"8e00",
---- 533=>x"8b00", 534=>x"8900", 535=>x"9500", 536=>x"8e00",
---- 537=>x"8800", 538=>x"8a00", 539=>x"9600", 540=>x"8c00",
---- 541=>x"8900", 542=>x"8f00", 543=>x"9a00", 544=>x"8a00",
---- 545=>x"8a00", 546=>x"9400", 547=>x"a100", 548=>x"8700",
---- 549=>x"8b00", 550=>x"9800", 551=>x"9f00", 552=>x"8600",
---- 553=>x"8d00", 554=>x"9c00", 555=>x"9f00", 556=>x"8700",
---- 557=>x"9200", 558=>x"a000", 559=>x"a000", 560=>x"8900",
---- 561=>x"9b00", 562=>x"a000", 563=>x"9d00", 564=>x"8d00",
---- 565=>x"9d00", 566=>x"9e00", 567=>x"9d00", 568=>x"9100",
---- 569=>x"9c00", 570=>x"9d00", 571=>x"9b00", 572=>x"9800",
---- 573=>x"9d00", 574=>x"9c00", 575=>x"9c00", 576=>x"9c00",
---- 577=>x"9f00", 578=>x"9e00", 579=>x"9b00", 580=>x"a000",
---- 581=>x"9e00", 582=>x"9c00", 583=>x"9b00", 584=>x"9f00",
---- 585=>x"9e00", 586=>x"9b00", 587=>x"9b00", 588=>x"a100",
---- 589=>x"a000", 590=>x"9d00", 591=>x"9c00", 592=>x"a100",
---- 593=>x"9d00", 594=>x"9a00", 595=>x"9900", 596=>x"a100",
---- 597=>x"9d00", 598=>x"9b00", 599=>x"9800", 600=>x"a000",
---- 601=>x"9c00", 602=>x"9c00", 603=>x"9a00", 604=>x"9c00",
---- 605=>x"9d00", 606=>x"9c00", 607=>x"9a00", 608=>x"9e00",
---- 609=>x"9c00", 610=>x"9c00", 611=>x"9a00", 612=>x"5e00",
---- 613=>x"9d00", 614=>x"9c00", 615=>x"9a00", 616=>x"9d00",
---- 617=>x"9c00", 618=>x"9a00", 619=>x"9900", 620=>x"9e00",
---- 621=>x"9c00", 622=>x"9500", 623=>x"9800", 624=>x"9d00",
---- 625=>x"9b00", 626=>x"9600", 627=>x"9800", 628=>x"9b00",
---- 629=>x"9800", 630=>x"9b00", 631=>x"9800", 632=>x"9a00",
---- 633=>x"9a00", 634=>x"9800", 635=>x"9500", 636=>x"9b00",
---- 637=>x"9b00", 638=>x"9700", 639=>x"9600", 640=>x"9800",
---- 641=>x"9900", 642=>x"9900", 643=>x"9600", 644=>x"9a00",
---- 645=>x"9900", 646=>x"9600", 647=>x"9500", 648=>x"9900",
---- 649=>x"9500", 650=>x"9600", 651=>x"9700", 652=>x"9600",
---- 653=>x"9500", 654=>x"9700", 655=>x"9600", 656=>x"9900",
---- 657=>x"9600", 658=>x"9800", 659=>x"9700", 660=>x"9700",
---- 661=>x"9900", 662=>x"9800", 663=>x"9700", 664=>x"9700",
---- 665=>x"9700", 666=>x"9900", 667=>x"9500", 668=>x"6900",
---- 669=>x"9600", 670=>x"9700", 671=>x"9800", 672=>x"9600",
---- 673=>x"9900", 674=>x"9600", 675=>x"9600", 676=>x"9600",
---- 677=>x"9600", 678=>x"9600", 679=>x"9300", 680=>x"9800",
---- 681=>x"9500", 682=>x"9400", 683=>x"9800", 684=>x"9800",
---- 685=>x"9400", 686=>x"9400", 687=>x"9600", 688=>x"9700",
---- 689=>x"9600", 690=>x"9200", 691=>x"6b00", 692=>x"9600",
---- 693=>x"9400", 694=>x"9300", 695=>x"9200", 696=>x"9500",
---- 697=>x"9400", 698=>x"9400", 699=>x"9200", 700=>x"9700",
---- 701=>x"9600", 702=>x"9500", 703=>x"9300", 704=>x"9800",
---- 705=>x"9600", 706=>x"9700", 707=>x"9400", 708=>x"9800",
---- 709=>x"9600", 710=>x"9a00", 711=>x"6b00", 712=>x"9a00",
---- 713=>x"9800", 714=>x"9800", 715=>x"9500", 716=>x"9800",
---- 717=>x"9900", 718=>x"9500", 719=>x"9900", 720=>x"9a00",
---- 721=>x"9800", 722=>x"9900", 723=>x"9800", 724=>x"9b00",
---- 725=>x"9800", 726=>x"9600", 727=>x"9700", 728=>x"9b00",
---- 729=>x"9900", 730=>x"9700", 731=>x"9a00", 732=>x"9c00",
---- 733=>x"9900", 734=>x"9c00", 735=>x"9d00", 736=>x"9a00",
---- 737=>x"9a00", 738=>x"9b00", 739=>x"9a00", 740=>x"9900",
---- 741=>x"9800", 742=>x"9700", 743=>x"9800", 744=>x"9600",
---- 745=>x"9800", 746=>x"9500", 747=>x"9800", 748=>x"9800",
---- 749=>x"9900", 750=>x"9600", 751=>x"9800", 752=>x"9600",
---- 753=>x"9500", 754=>x"9500", 755=>x"9700", 756=>x"9700",
---- 757=>x"9600", 758=>x"9800", 759=>x"6b00", 760=>x"9700",
---- 761=>x"9700", 762=>x"9500", 763=>x"9400", 764=>x"9600",
---- 765=>x"9600", 766=>x"9500", 767=>x"9400", 768=>x"9700",
---- 769=>x"9400", 770=>x"9800", 771=>x"9500", 772=>x"6e00",
---- 773=>x"9300", 774=>x"9200", 775=>x"9300", 776=>x"8800",
---- 777=>x"8c00", 778=>x"8c00", 779=>x"8b00", 780=>x"7c00",
---- 781=>x"7d00", 782=>x"8100", 783=>x"8500", 784=>x"7200",
---- 785=>x"7500", 786=>x"7600", 787=>x"7600", 788=>x"6d00",
---- 789=>x"6d00", 790=>x"6d00", 791=>x"6d00", 792=>x"6a00",
---- 793=>x"6900", 794=>x"6b00", 795=>x"6800", 796=>x"6f00",
---- 797=>x"6b00", 798=>x"6900", 799=>x"6500", 800=>x"7a00",
---- 801=>x"7400", 802=>x"9300", 803=>x"6b00", 804=>x"8000",
---- 805=>x"7b00", 806=>x"7a00", 807=>x"7500", 808=>x"8600",
---- 809=>x"8000", 810=>x"7e00", 811=>x"7900", 812=>x"8800",
---- 813=>x"8500", 814=>x"8200", 815=>x"7f00", 816=>x"8800",
---- 817=>x"8700", 818=>x"8700", 819=>x"8200", 820=>x"8900",
---- 821=>x"8700", 822=>x"8a00", 823=>x"8800", 824=>x"8b00",
---- 825=>x"8a00", 826=>x"8900", 827=>x"8900", 828=>x"8d00",
---- 829=>x"8a00", 830=>x"8a00", 831=>x"8600", 832=>x"8d00",
---- 833=>x"8c00", 834=>x"8d00", 835=>x"8700", 836=>x"8d00",
---- 837=>x"8d00", 838=>x"8b00", 839=>x"8b00", 840=>x"8d00",
---- 841=>x"8b00", 842=>x"8a00", 843=>x"8a00", 844=>x"8d00",
---- 845=>x"8a00", 846=>x"7300", 847=>x"8a00", 848=>x"8a00",
---- 849=>x"8600", 850=>x"8900", 851=>x"8b00", 852=>x"8900",
---- 853=>x"8800", 854=>x"8600", 855=>x"8900", 856=>x"8a00",
---- 857=>x"8800", 858=>x"8700", 859=>x"8600", 860=>x"8400",
---- 861=>x"8400", 862=>x"8500", 863=>x"8600", 864=>x"8500",
---- 865=>x"8500", 866=>x"8700", 867=>x"8400", 868=>x"8900",
---- 869=>x"8600", 870=>x"8500", 871=>x"8500", 872=>x"8700",
---- 873=>x"8400", 874=>x"8700", 875=>x"8600", 876=>x"8900",
---- 877=>x"8500", 878=>x"8300", 879=>x"8400", 880=>x"8900",
---- 881=>x"8700", 882=>x"8500", 883=>x"8400", 884=>x"8900",
---- 885=>x"8700", 886=>x"8800", 887=>x"8200", 888=>x"8d00",
---- 889=>x"8700", 890=>x"8800", 891=>x"8100", 892=>x"8a00",
---- 893=>x"8600", 894=>x"8800", 895=>x"8700", 896=>x"8a00",
---- 897=>x"8a00", 898=>x"8600", 899=>x"8300", 900=>x"8900",
---- 901=>x"8800", 902=>x"8500", 903=>x"8200", 904=>x"8c00",
---- 905=>x"8b00", 906=>x"8800", 907=>x"8500", 908=>x"8a00",
---- 909=>x"8800", 910=>x"8800", 911=>x"8400", 912=>x"8e00",
---- 913=>x"8b00", 914=>x"8b00", 915=>x"8800", 916=>x"8d00",
---- 917=>x"8c00", 918=>x"8b00", 919=>x"8c00", 920=>x"8c00",
---- 921=>x"8e00", 922=>x"8e00", 923=>x"8b00", 924=>x"8800",
---- 925=>x"8a00", 926=>x"8c00", 927=>x"8e00", 928=>x"7900",
---- 929=>x"7c00", 930=>x"8600", 931=>x"8900", 932=>x"6500",
---- 933=>x"6900", 934=>x"7300", 935=>x"7c00", 936=>x"4f00",
---- 937=>x"4d00", 938=>x"5a00", 939=>x"6700", 940=>x"3300",
---- 941=>x"3500", 942=>x"3d00", 943=>x"4800", 944=>x"2b00",
---- 945=>x"2f00", 946=>x"2900", 947=>x"3000", 948=>x"2e00",
---- 949=>x"2900", 950=>x"2300", 951=>x"2700", 952=>x"2d00",
---- 953=>x"2d00", 954=>x"2800", 955=>x"2600", 956=>x"3900",
---- 957=>x"2f00", 958=>x"2a00", 959=>x"2900", 960=>x"4200",
---- 961=>x"3600", 962=>x"2e00", 963=>x"2e00", 964=>x"4800",
---- 965=>x"4200", 966=>x"3c00", 967=>x"3800", 968=>x"5100",
---- 969=>x"4b00", 970=>x"4a00", 971=>x"4d00", 972=>x"5400",
---- 973=>x"5400", 974=>x"5700", 975=>x"5900", 976=>x"5800",
---- 977=>x"5e00", 978=>x"5f00", 979=>x"5e00", 980=>x"6500",
---- 981=>x"6600", 982=>x"6a00", 983=>x"6600", 984=>x"6800",
---- 985=>x"6d00", 986=>x"6f00", 987=>x"6f00", 988=>x"7000",
---- 989=>x"7400", 990=>x"7400", 991=>x"7100", 992=>x"7500",
---- 993=>x"7400", 994=>x"7400", 995=>x"7200", 996=>x"7600",
---- 997=>x"7900", 998=>x"7600", 999=>x"7200", 1000=>x"7600",
---- 1001=>x"7700", 1002=>x"7200", 1003=>x"7300", 1004=>x"7c00",
---- 1005=>x"7300", 1006=>x"7600", 1007=>x"7400", 1008=>x"7600",
---- 1009=>x"7900", 1010=>x"8700", 1011=>x"7500", 1012=>x"7700",
---- 1013=>x"7c00", 1014=>x"7c00", 1015=>x"7a00", 1016=>x"7d00",
---- 1017=>x"8200", 1018=>x"7f00", 1019=>x"7b00", 1020=>x"8200",
---- 1021=>x"8700", 1022=>x"8300", 1023=>x"7d00"),
----
---- 52 => (0=>x"da00", 1=>x"d300", 2=>x"c000", 3=>x"9600", 4=>x"da00",
---- 5=>x"d300", 6=>x"c000", 7=>x"9500", 8=>x"db00",
---- 9=>x"d400", 10=>x"c100", 11=>x"9800", 12=>x"db00",
---- 13=>x"d900", 14=>x"ce00", 15=>x"b100", 16=>x"d900",
---- 17=>x"d900", 18=>x"2a00", 19=>x"c200", 20=>x"d900",
---- 21=>x"db00", 22=>x"d900", 23=>x"d000", 24=>x"db00",
---- 25=>x"db00", 26=>x"da00", 27=>x"d800", 28=>x"d800",
---- 29=>x"d900", 30=>x"db00", 31=>x"db00", 32=>x"d800",
---- 33=>x"d900", 34=>x"dc00", 35=>x"dc00", 36=>x"d500",
---- 37=>x"d900", 38=>x"da00", 39=>x"db00", 40=>x"d000",
---- 41=>x"d600", 42=>x"d900", 43=>x"dc00", 44=>x"cc00",
---- 45=>x"d300", 46=>x"d700", 47=>x"d900", 48=>x"c300",
---- 49=>x"cf00", 50=>x"d600", 51=>x"d800", 52=>x"b500",
---- 53=>x"cc00", 54=>x"d300", 55=>x"d700", 56=>x"a100",
---- 57=>x"c200", 58=>x"d000", 59=>x"d700", 60=>x"9000",
---- 61=>x"b000", 62=>x"ca00", 63=>x"d200", 64=>x"8a00",
---- 65=>x"9800", 66=>x"b800", 67=>x"3700", 68=>x"8c00",
---- 69=>x"8f00", 70=>x"aa00", 71=>x"c800", 72=>x"9000",
---- 73=>x"8e00", 74=>x"9700", 75=>x"b900", 76=>x"8e00",
---- 77=>x"8d00", 78=>x"8c00", 79=>x"a300", 80=>x"8f00",
---- 81=>x"8e00", 82=>x"8c00", 83=>x"9200", 84=>x"8e00",
---- 85=>x"8c00", 86=>x"8c00", 87=>x"8b00", 88=>x"8d00",
---- 89=>x"8e00", 90=>x"8c00", 91=>x"8e00", 92=>x"8e00",
---- 93=>x"9000", 94=>x"9000", 95=>x"8e00", 96=>x"8f00",
---- 97=>x"8e00", 98=>x"8f00", 99=>x"8c00", 100=>x"8e00",
---- 101=>x"8b00", 102=>x"8d00", 103=>x"8c00", 104=>x"8c00",
---- 105=>x"8e00", 106=>x"8e00", 107=>x"8c00", 108=>x"8d00",
---- 109=>x"8c00", 110=>x"8e00", 111=>x"8d00", 112=>x"8d00",
---- 113=>x"8e00", 114=>x"8e00", 115=>x"8c00", 116=>x"8b00",
---- 117=>x"8a00", 118=>x"8e00", 119=>x"8c00", 120=>x"8d00",
---- 121=>x"8c00", 122=>x"8d00", 123=>x"8e00", 124=>x"8e00",
---- 125=>x"8e00", 126=>x"8f00", 127=>x"8e00", 128=>x"8a00",
---- 129=>x"8b00", 130=>x"9200", 131=>x"9000", 132=>x"8c00",
---- 133=>x"8d00", 134=>x"9000", 135=>x"9100", 136=>x"8e00",
---- 137=>x"8f00", 138=>x"8f00", 139=>x"9200", 140=>x"9000",
---- 141=>x"9000", 142=>x"8e00", 143=>x"9000", 144=>x"9100",
---- 145=>x"9000", 146=>x"6f00", 147=>x"9000", 148=>x"9000",
---- 149=>x"9000", 150=>x"9100", 151=>x"9400", 152=>x"9000",
---- 153=>x"9200", 154=>x"9200", 155=>x"9300", 156=>x"9000",
---- 157=>x"8c00", 158=>x"9300", 159=>x"9100", 160=>x"8f00",
---- 161=>x"9000", 162=>x"6c00", 163=>x"9000", 164=>x"9200",
---- 165=>x"9100", 166=>x"9100", 167=>x"9400", 168=>x"9000",
---- 169=>x"9100", 170=>x"9100", 171=>x"9200", 172=>x"8e00",
---- 173=>x"8f00", 174=>x"9000", 175=>x"9100", 176=>x"8d00",
---- 177=>x"8f00", 178=>x"9000", 179=>x"9100", 180=>x"9000",
---- 181=>x"9200", 182=>x"9400", 183=>x"9300", 184=>x"9100",
---- 185=>x"9100", 186=>x"9300", 187=>x"9600", 188=>x"9100",
---- 189=>x"9100", 190=>x"9300", 191=>x"9500", 192=>x"9200",
---- 193=>x"9300", 194=>x"9700", 195=>x"9900", 196=>x"9200",
---- 197=>x"9600", 198=>x"9a00", 199=>x"9a00", 200=>x"9300",
---- 201=>x"6800", 202=>x"9b00", 203=>x"9700", 204=>x"9500",
---- 205=>x"9b00", 206=>x"9900", 207=>x"8700", 208=>x"9800",
---- 209=>x"9a00", 210=>x"9200", 211=>x"6200", 212=>x"9900",
---- 213=>x"9700", 214=>x"7500", 215=>x"3c00", 216=>x"9b00",
---- 217=>x"8b00", 218=>x"4d00", 219=>x"2900", 220=>x"9200",
---- 221=>x"6200", 222=>x"3000", 223=>x"2a00", 224=>x"7400",
---- 225=>x"3a00", 226=>x"2900", 227=>x"2a00", 228=>x"b600",
---- 229=>x"2900", 230=>x"2b00", 231=>x"2d00", 232=>x"5b00",
---- 233=>x"1d00", 234=>x"2c00", 235=>x"2d00", 236=>x"9100",
---- 237=>x"2000", 238=>x"2b00", 239=>x"2c00", 240=>x"c600",
---- 241=>x"3800", 242=>x"2700", 243=>x"2c00", 244=>x"de00",
---- 245=>x"5700", 246=>x"2200", 247=>x"2c00", 248=>x"e400",
---- 249=>x"7700", 250=>x"2300", 251=>x"2c00", 252=>x"eb00",
---- 253=>x"7500", 254=>x"2200", 255=>x"2c00", 256=>x"ec00",
---- 257=>x"8800", 258=>x"1f00", 259=>x"2a00", 260=>x"e900",
---- 261=>x"8600", 262=>x"1c00", 263=>x"2900", 264=>x"e400",
---- 265=>x"7b00", 266=>x"2000", 267=>x"2d00", 268=>x"e200",
---- 269=>x"6800", 270=>x"2500", 271=>x"2a00", 272=>x"d800",
---- 273=>x"4c00", 274=>x"2700", 275=>x"3000", 276=>x"c700",
---- 277=>x"3a00", 278=>x"2600", 279=>x"2c00", 280=>x"b100",
---- 281=>x"2c00", 282=>x"d400", 283=>x"3300", 284=>x"9400",
---- 285=>x"2700", 286=>x"3100", 287=>x"3100", 288=>x"7d00",
---- 289=>x"2000", 290=>x"3100", 291=>x"3300", 292=>x"5d00",
---- 293=>x"1e00", 294=>x"2f00", 295=>x"2c00", 296=>x"3c00",
---- 297=>x"2100", 298=>x"2c00", 299=>x"2b00", 300=>x"2800",
---- 301=>x"2400", 302=>x"2c00", 303=>x"2e00", 304=>x"2300",
---- 305=>x"2800", 306=>x"2b00", 307=>x"2a00", 308=>x"2500",
---- 309=>x"2b00", 310=>x"2b00", 311=>x"2d00", 312=>x"2a00",
---- 313=>x"3400", 314=>x"3500", 315=>x"3100", 316=>x"2800",
---- 317=>x"3300", 318=>x"3b00", 319=>x"3200", 320=>x"2800",
---- 321=>x"2800", 322=>x"3100", 323=>x"3a00", 324=>x"2800",
---- 325=>x"2a00", 326=>x"3200", 327=>x"3400", 328=>x"2b00",
---- 329=>x"2c00", 330=>x"3000", 331=>x"3100", 332=>x"3100",
---- 333=>x"2f00", 334=>x"3000", 335=>x"3200", 336=>x"2f00",
---- 337=>x"3500", 338=>x"3500", 339=>x"3100", 340=>x"3100",
---- 341=>x"3600", 342=>x"3700", 343=>x"3100", 344=>x"2f00",
---- 345=>x"2e00", 346=>x"3000", 347=>x"2d00", 348=>x"3100",
---- 349=>x"3100", 350=>x"3200", 351=>x"2c00", 352=>x"3000",
---- 353=>x"2f00", 354=>x"3200", 355=>x"2b00", 356=>x"2f00",
---- 357=>x"3000", 358=>x"2e00", 359=>x"2a00", 360=>x"3000",
---- 361=>x"3000", 362=>x"2d00", 363=>x"3100", 364=>x"3400",
---- 365=>x"3300", 366=>x"3100", 367=>x"2a00", 368=>x"3000",
---- 369=>x"3200", 370=>x"3400", 371=>x"3200", 372=>x"3000",
---- 373=>x"2b00", 374=>x"3100", 375=>x"3300", 376=>x"2e00",
---- 377=>x"2d00", 378=>x"3200", 379=>x"3500", 380=>x"2c00",
---- 381=>x"2b00", 382=>x"3300", 383=>x"3b00", 384=>x"2a00",
---- 385=>x"2a00", 386=>x"3400", 387=>x"4000", 388=>x"3200",
---- 389=>x"2e00", 390=>x"3600", 391=>x"3500", 392=>x"3000",
---- 393=>x"3300", 394=>x"3600", 395=>x"3500", 396=>x"2f00",
---- 397=>x"3400", 398=>x"3600", 399=>x"3400", 400=>x"3100",
---- 401=>x"3400", 402=>x"3300", 403=>x"3100", 404=>x"3000",
---- 405=>x"3300", 406=>x"3500", 407=>x"2f00", 408=>x"ce00",
---- 409=>x"3500", 410=>x"3400", 411=>x"3600", 412=>x"3700",
---- 413=>x"3900", 414=>x"3200", 415=>x"3b00", 416=>x"3800",
---- 417=>x"3300", 418=>x"3400", 419=>x"3d00", 420=>x"3600",
---- 421=>x"2f00", 422=>x"3600", 423=>x"4400", 424=>x"3000",
---- 425=>x"3300", 426=>x"3e00", 427=>x"4a00", 428=>x"3000",
---- 429=>x"3400", 430=>x"3e00", 431=>x"5800", 432=>x"2e00",
---- 433=>x"3100", 434=>x"b800", 435=>x"6c00", 436=>x"2e00",
---- 437=>x"3500", 438=>x"5300", 439=>x"7b00", 440=>x"3200",
---- 441=>x"3f00", 442=>x"6300", 443=>x"8400", 444=>x"3700",
---- 445=>x"4c00", 446=>x"7700", 447=>x"8b00", 448=>x"3900",
---- 449=>x"5f00", 450=>x"8400", 451=>x"9200", 452=>x"3b00",
---- 453=>x"6e00", 454=>x"8c00", 455=>x"8f00", 456=>x"4a00",
---- 457=>x"7900", 458=>x"8e00", 459=>x"8c00", 460=>x"6100",
---- 461=>x"8600", 462=>x"9000", 463=>x"8c00", 464=>x"7a00",
---- 465=>x"9100", 466=>x"8f00", 467=>x"8700", 468=>x"8500",
---- 469=>x"9200", 470=>x"8e00", 471=>x"8400", 472=>x"8900",
---- 473=>x"9000", 474=>x"8800", 475=>x"8500", 476=>x"8b00",
---- 477=>x"8b00", 478=>x"8600", 479=>x"7600", 480=>x"8d00",
---- 481=>x"8700", 482=>x"8000", 483=>x"8a00", 484=>x"8d00",
---- 485=>x"8500", 486=>x"8100", 487=>x"9000", 488=>x"8900",
---- 489=>x"8200", 490=>x"8400", 491=>x"9500", 492=>x"8700",
---- 493=>x"8100", 494=>x"8900", 495=>x"9a00", 496=>x"8500",
---- 497=>x"7e00", 498=>x"9000", 499=>x"9f00", 500=>x"7f00",
---- 501=>x"8400", 502=>x"9600", 503=>x"a200", 504=>x"8000",
---- 505=>x"8d00", 506=>x"9c00", 507=>x"a100", 508=>x"8000",
---- 509=>x"8f00", 510=>x"9e00", 511=>x"a000", 512=>x"8300",
---- 513=>x"9600", 514=>x"a000", 515=>x"a000", 516=>x"8a00",
---- 517=>x"9900", 518=>x"a000", 519=>x"a000", 520=>x"9500",
---- 521=>x"a100", 522=>x"a100", 523=>x"a000", 524=>x"9900",
---- 525=>x"a300", 526=>x"9e00", 527=>x"9e00", 528=>x"9d00",
---- 529=>x"a000", 530=>x"9f00", 531=>x"9e00", 532=>x"9f00",
---- 533=>x"9e00", 534=>x"9f00", 535=>x"9c00", 536=>x"9e00",
---- 537=>x"9e00", 538=>x"9f00", 539=>x"9d00", 540=>x"9e00",
---- 541=>x"9d00", 542=>x"9c00", 543=>x"9c00", 544=>x"9f00",
---- 545=>x"9d00", 546=>x"9b00", 547=>x"9b00", 548=>x"9d00",
---- 549=>x"9a00", 550=>x"9d00", 551=>x"9a00", 552=>x"9b00",
---- 553=>x"9b00", 554=>x"9c00", 555=>x"9d00", 556=>x"9e00",
---- 557=>x"9b00", 558=>x"9b00", 559=>x"9a00", 560=>x"9e00",
---- 561=>x"9900", 562=>x"9a00", 563=>x"9900", 564=>x"9b00",
---- 565=>x"9700", 566=>x"9a00", 567=>x"9b00", 568=>x"9a00",
---- 569=>x"9b00", 570=>x"9800", 571=>x"9900", 572=>x"9d00",
---- 573=>x"9b00", 574=>x"9800", 575=>x"9700", 576=>x"6400",
---- 577=>x"9900", 578=>x"9a00", 579=>x"9600", 580=>x"9c00",
---- 581=>x"9800", 582=>x"9900", 583=>x"9900", 584=>x"9900",
---- 585=>x"9800", 586=>x"9a00", 587=>x"9700", 588=>x"9b00",
---- 589=>x"9b00", 590=>x"9b00", 591=>x"9a00", 592=>x"9a00",
---- 593=>x"9c00", 594=>x"9a00", 595=>x"9800", 596=>x"9900",
---- 597=>x"9a00", 598=>x"9900", 599=>x"9900", 600=>x"9b00",
---- 601=>x"9b00", 602=>x"9a00", 603=>x"9700", 604=>x"9d00",
---- 605=>x"9900", 606=>x"9900", 607=>x"9800", 608=>x"9800",
---- 609=>x"9900", 610=>x"9900", 611=>x"9700", 612=>x"9b00",
---- 613=>x"9a00", 614=>x"9a00", 615=>x"9800", 616=>x"9900",
---- 617=>x"9a00", 618=>x"9b00", 619=>x"9700", 620=>x"9b00",
---- 621=>x"9b00", 622=>x"9b00", 623=>x"9900", 624=>x"9700",
---- 625=>x"9900", 626=>x"9700", 627=>x"9a00", 628=>x"9700",
---- 629=>x"9700", 630=>x"9400", 631=>x"9700", 632=>x"9700",
---- 633=>x"9700", 634=>x"9600", 635=>x"9300", 636=>x"9600",
---- 637=>x"9500", 638=>x"9700", 639=>x"6a00", 640=>x"9600",
---- 641=>x"9700", 642=>x"9700", 643=>x"6900", 644=>x"9700",
---- 645=>x"9700", 646=>x"9600", 647=>x"9600", 648=>x"9500",
---- 649=>x"9400", 650=>x"9400", 651=>x"9600", 652=>x"9600",
---- 653=>x"9500", 654=>x"9700", 655=>x"9800", 656=>x"9500",
---- 657=>x"9500", 658=>x"9800", 659=>x"9500", 660=>x"9400",
---- 661=>x"9600", 662=>x"6b00", 663=>x"9400", 664=>x"9400",
---- 665=>x"9500", 666=>x"9500", 667=>x"9200", 668=>x"9200",
---- 669=>x"9400", 670=>x"9600", 671=>x"9600", 672=>x"9400",
---- 673=>x"9500", 674=>x"9400", 675=>x"9300", 676=>x"9300",
---- 677=>x"9500", 678=>x"9400", 679=>x"9500", 680=>x"9300",
---- 681=>x"9400", 682=>x"9600", 683=>x"9400", 684=>x"9200",
---- 685=>x"9300", 686=>x"9500", 687=>x"9400", 688=>x"9400",
---- 689=>x"9600", 690=>x"9500", 691=>x"9300", 692=>x"9300",
---- 693=>x"9800", 694=>x"9300", 695=>x"9200", 696=>x"9300",
---- 697=>x"9400", 698=>x"9400", 699=>x"9400", 700=>x"9400",
---- 701=>x"9500", 702=>x"9400", 703=>x"9100", 704=>x"9200",
---- 705=>x"9500", 706=>x"9300", 707=>x"9200", 708=>x"9100",
---- 709=>x"9300", 710=>x"9200", 711=>x"9000", 712=>x"9500",
---- 713=>x"9700", 714=>x"6b00", 715=>x"9300", 716=>x"9800",
---- 717=>x"9600", 718=>x"9500", 719=>x"9700", 720=>x"9700",
---- 721=>x"9500", 722=>x"9500", 723=>x"9800", 724=>x"9500",
---- 725=>x"9500", 726=>x"9500", 727=>x"9400", 728=>x"9900",
---- 729=>x"9700", 730=>x"9500", 731=>x"9500", 732=>x"9d00",
---- 733=>x"9a00", 734=>x"9800", 735=>x"9700", 736=>x"9a00",
---- 737=>x"9600", 738=>x"9700", 739=>x"9600", 740=>x"9700",
---- 741=>x"9900", 742=>x"9500", 743=>x"9500", 744=>x"9900",
---- 745=>x"9b00", 746=>x"9600", 747=>x"9400", 748=>x"9900",
---- 749=>x"9700", 750=>x"9600", 751=>x"9800", 752=>x"9800",
---- 753=>x"9800", 754=>x"9800", 755=>x"9700", 756=>x"9500",
---- 757=>x"9700", 758=>x"9500", 759=>x"9400", 760=>x"9700",
---- 761=>x"9500", 762=>x"9500", 763=>x"9400", 764=>x"9400",
---- 765=>x"9600", 766=>x"9500", 767=>x"9200", 768=>x"9700",
---- 769=>x"9300", 770=>x"9400", 771=>x"9300", 772=>x"9400",
---- 773=>x"9500", 774=>x"9200", 775=>x"9100", 776=>x"8f00",
---- 777=>x"9600", 778=>x"9500", 779=>x"9300", 780=>x"8700",
---- 781=>x"8b00", 782=>x"7200", 783=>x"8f00", 784=>x"7c00",
---- 785=>x"8000", 786=>x"8100", 787=>x"8400", 788=>x"6f00",
---- 789=>x"7200", 790=>x"7500", 791=>x"7900", 792=>x"6600",
---- 793=>x"6600", 794=>x"6900", 795=>x"7000", 796=>x"6500",
---- 797=>x"6400", 798=>x"6400", 799=>x"6200", 800=>x"6a00",
---- 801=>x"6400", 802=>x"6400", 803=>x"6100", 804=>x"7100",
---- 805=>x"6e00", 806=>x"6900", 807=>x"6500", 808=>x"7a00",
---- 809=>x"7600", 810=>x"7200", 811=>x"6b00", 812=>x"7e00",
---- 813=>x"7a00", 814=>x"7500", 815=>x"7500", 816=>x"8100",
---- 817=>x"7d00", 818=>x"7b00", 819=>x"7900", 820=>x"8200",
---- 821=>x"7f00", 822=>x"8300", 823=>x"8100", 824=>x"8700",
---- 825=>x"8200", 826=>x"8200", 827=>x"8000", 828=>x"8600",
---- 829=>x"8600", 830=>x"8200", 831=>x"8400", 832=>x"8500",
---- 833=>x"8600", 834=>x"8500", 835=>x"8400", 836=>x"8600",
---- 837=>x"8700", 838=>x"8600", 839=>x"8200", 840=>x"8700",
---- 841=>x"8a00", 842=>x"8400", 843=>x"8500", 844=>x"8900",
---- 845=>x"8900", 846=>x"8600", 847=>x"8300", 848=>x"8900",
---- 849=>x"8300", 850=>x"8700", 851=>x"8300", 852=>x"8600",
---- 853=>x"8500", 854=>x"8500", 855=>x"8100", 856=>x"8700",
---- 857=>x"8400", 858=>x"8200", 859=>x"8000", 860=>x"8600",
---- 861=>x"8200", 862=>x"8000", 863=>x"7d00", 864=>x"8100",
---- 865=>x"8100", 866=>x"8200", 867=>x"7e00", 868=>x"7f00",
---- 869=>x"7f00", 870=>x"8000", 871=>x"7e00", 872=>x"8200",
---- 873=>x"7f00", 874=>x"8200", 875=>x"7c00", 876=>x"8200",
---- 877=>x"7e00", 878=>x"7c00", 879=>x"7900", 880=>x"8300",
---- 881=>x"7d00", 882=>x"7f00", 883=>x"7d00", 884=>x"8000",
---- 885=>x"8100", 886=>x"7b00", 887=>x"7a00", 888=>x"7e00",
---- 889=>x"7c00", 890=>x"7b00", 891=>x"7d00", 892=>x"7f00",
---- 893=>x"7f00", 894=>x"7f00", 895=>x"7f00", 896=>x"8200",
---- 897=>x"7e00", 898=>x"8000", 899=>x"8200", 900=>x"7e00",
---- 901=>x"8200", 902=>x"8500", 903=>x"8400", 904=>x"8000",
---- 905=>x"8300", 906=>x"8400", 907=>x"8500", 908=>x"8300",
---- 909=>x"8600", 910=>x"8800", 911=>x"8700", 912=>x"8800",
---- 913=>x"8800", 914=>x"8d00", 915=>x"8d00", 916=>x"8800",
---- 917=>x"6f00", 918=>x"9100", 919=>x"9300", 920=>x"8a00",
---- 921=>x"8d00", 922=>x"9600", 923=>x"9800", 924=>x"9200",
---- 925=>x"9500", 926=>x"9900", 927=>x"9b00", 928=>x"9000",
---- 929=>x"9900", 930=>x"a000", 931=>x"9e00", 932=>x"8900",
---- 933=>x"9100", 934=>x"9d00", 935=>x"a100", 936=>x"7700",
---- 937=>x"8600", 938=>x"8e00", 939=>x"9200", 940=>x"5b00",
---- 941=>x"6c00", 942=>x"7100", 943=>x"8900", 944=>x"3c00",
---- 945=>x"5000", 946=>x"6d00", 947=>x"a200", 948=>x"2b00",
---- 949=>x"4300", 950=>x"8a00", 951=>x"bd00", 952=>x"2000",
---- 953=>x"4500", 954=>x"9b00", 955=>x"c800", 956=>x"2700",
---- 957=>x"4500", 958=>x"9800", 959=>x"c400", 960=>x"3100",
---- 961=>x"4a00", 962=>x"8d00", 963=>x"b900", 964=>x"3d00",
---- 965=>x"4800", 966=>x"7e00", 967=>x"b500", 968=>x"4d00",
---- 969=>x"5700", 970=>x"8300", 971=>x"b700", 972=>x"5200",
---- 973=>x"5f00", 974=>x"8c00", 975=>x"b500", 976=>x"5900",
---- 977=>x"5e00", 978=>x"8800", 979=>x"b200", 980=>x"6100",
---- 981=>x"6100", 982=>x"7b00", 983=>x"a200", 984=>x"6900",
---- 985=>x"6800", 986=>x"7000", 987=>x"8900", 988=>x"7000",
---- 989=>x"7000", 990=>x"6d00", 991=>x"7100", 992=>x"7300",
---- 993=>x"7200", 994=>x"6e00", 995=>x"6b00", 996=>x"7200",
---- 997=>x"7100", 998=>x"8f00", 999=>x"6800", 1000=>x"7400",
---- 1001=>x"7200", 1002=>x"7000", 1003=>x"6d00", 1004=>x"7200",
---- 1005=>x"7400", 1006=>x"7100", 1007=>x"7000", 1008=>x"7300",
---- 1009=>x"7400", 1010=>x"7100", 1011=>x"6e00", 1012=>x"7500",
---- 1013=>x"7500", 1014=>x"7100", 1015=>x"7500", 1016=>x"7a00",
---- 1017=>x"7700", 1018=>x"7600", 1019=>x"7900", 1020=>x"7b00",
---- 1021=>x"7d00", 1022=>x"7d00", 1023=>x"8400"),
----
---- 53 => (0=>x"6c00", 1=>x"6500", 2=>x"6900", 3=>x"6c00", 4=>x"6a00",
---- 5=>x"6600", 6=>x"6900", 7=>x"6c00", 8=>x"6c00",
---- 9=>x"6500", 10=>x"9600", 11=>x"6d00", 12=>x"7f00",
---- 13=>x"6400", 14=>x"6600", 15=>x"6c00", 16=>x"9d00",
---- 17=>x"6f00", 18=>x"6700", 19=>x"6b00", 20=>x"b600",
---- 21=>x"8900", 22=>x"6800", 23=>x"6700", 24=>x"c800",
---- 25=>x"a600", 26=>x"8a00", 27=>x"6700", 28=>x"d300",
---- 29=>x"c000", 30=>x"9400", 31=>x"6a00", 32=>x"d900",
---- 33=>x"ce00", 34=>x"b300", 35=>x"8000", 36=>x"db00",
---- 37=>x"d600", 38=>x"c400", 39=>x"9c00", 40=>x"dc00",
---- 41=>x"da00", 42=>x"d100", 43=>x"b900", 44=>x"db00",
---- 45=>x"de00", 46=>x"da00", 47=>x"c900", 48=>x"db00",
---- 49=>x"dc00", 50=>x"db00", 51=>x"d300", 52=>x"da00",
---- 53=>x"dc00", 54=>x"de00", 55=>x"d900", 56=>x"2600",
---- 57=>x"db00", 58=>x"dd00", 59=>x"de00", 60=>x"d800",
---- 61=>x"da00", 62=>x"dd00", 63=>x"de00", 64=>x"cf00",
---- 65=>x"d600", 66=>x"2400", 67=>x"2200", 68=>x"d200",
---- 69=>x"d700", 70=>x"db00", 71=>x"df00", 72=>x"ce00",
---- 73=>x"d700", 74=>x"db00", 75=>x"dd00", 76=>x"c600",
---- 77=>x"d200", 78=>x"d800", 79=>x"dd00", 80=>x"b700",
---- 81=>x"ce00", 82=>x"d600", 83=>x"db00", 84=>x"a200",
---- 85=>x"c500", 86=>x"d200", 87=>x"d900", 88=>x"9100",
---- 89=>x"b400", 90=>x"ce00", 91=>x"d500", 92=>x"8c00",
---- 93=>x"9e00", 94=>x"c200", 95=>x"d000", 96=>x"8e00",
---- 97=>x"9200", 98=>x"ae00", 99=>x"cb00", 100=>x"8e00",
---- 101=>x"8f00", 102=>x"9a00", 103=>x"bc00", 104=>x"8c00",
---- 105=>x"8d00", 106=>x"8f00", 107=>x"a700", 108=>x"8b00",
---- 109=>x"8d00", 110=>x"8a00", 111=>x"8d00", 112=>x"8b00",
---- 113=>x"8d00", 114=>x"8a00", 115=>x"8700", 116=>x"8d00",
---- 117=>x"8d00", 118=>x"8b00", 119=>x"8800", 120=>x"8e00",
---- 121=>x"8f00", 122=>x"8d00", 123=>x"8a00", 124=>x"9000",
---- 125=>x"8f00", 126=>x"8c00", 127=>x"8c00", 128=>x"9000",
---- 129=>x"9100", 130=>x"8e00", 131=>x"8d00", 132=>x"8f00",
---- 133=>x"8f00", 134=>x"9100", 135=>x"8e00", 136=>x"7200",
---- 137=>x"8f00", 138=>x"9100", 139=>x"9100", 140=>x"9100",
---- 141=>x"9000", 142=>x"6e00", 143=>x"9200", 144=>x"9200",
---- 145=>x"9200", 146=>x"9400", 147=>x"9500", 148=>x"9200",
---- 149=>x"9100", 150=>x"9600", 151=>x"9400", 152=>x"9000",
---- 153=>x"9200", 154=>x"9400", 155=>x"9700", 156=>x"9100",
---- 157=>x"9600", 158=>x"9500", 159=>x"9800", 160=>x"9400",
---- 161=>x"9400", 162=>x"9600", 163=>x"9400", 164=>x"9300",
---- 165=>x"9400", 166=>x"9400", 167=>x"9a00", 168=>x"9400",
---- 169=>x"9500", 170=>x"9600", 171=>x"9c00", 172=>x"9300",
---- 173=>x"9600", 174=>x"9a00", 175=>x"9d00", 176=>x"9400",
---- 177=>x"9600", 178=>x"9c00", 179=>x"9900", 180=>x"9700",
---- 181=>x"9b00", 182=>x"9900", 183=>x"7e00", 184=>x"9900",
---- 185=>x"a000", 186=>x"8f00", 187=>x"5600", 188=>x"9b00",
---- 189=>x"9a00", 190=>x"7400", 191=>x"3500", 192=>x"6400",
---- 193=>x"8400", 194=>x"4a00", 195=>x"2e00", 196=>x"8f00",
---- 197=>x"6200", 198=>x"2c00", 199=>x"2900", 200=>x"7300",
---- 201=>x"3800", 202=>x"2600", 203=>x"2900", 204=>x"4900",
---- 205=>x"2900", 206=>x"2500", 207=>x"2800", 208=>x"2d00",
---- 209=>x"2a00", 210=>x"2900", 211=>x"2e00", 212=>x"2800",
---- 213=>x"2c00", 214=>x"2800", 215=>x"2a00", 216=>x"2b00",
---- 217=>x"2b00", 218=>x"2b00", 219=>x"2c00", 220=>x"2b00",
---- 221=>x"2d00", 222=>x"2c00", 223=>x"2f00", 224=>x"2d00",
---- 225=>x"3000", 226=>x"3200", 227=>x"2f00", 228=>x"2a00",
---- 229=>x"3500", 230=>x"2d00", 231=>x"3100", 232=>x"2d00",
---- 233=>x"2f00", 234=>x"2e00", 235=>x"3100", 236=>x"2f00",
---- 237=>x"2e00", 238=>x"3100", 239=>x"3a00", 240=>x"2e00",
---- 241=>x"2d00", 242=>x"2f00", 243=>x"3400", 244=>x"2c00",
---- 245=>x"2e00", 246=>x"3200", 247=>x"3200", 248=>x"2c00",
---- 249=>x"d000", 250=>x"3200", 251=>x"3400", 252=>x"2b00",
---- 253=>x"2c00", 254=>x"2e00", 255=>x"3200", 256=>x"2c00",
---- 257=>x"2e00", 258=>x"3400", 259=>x"3700", 260=>x"2e00",
---- 261=>x"3100", 262=>x"3500", 263=>x"3c00", 264=>x"2f00",
---- 265=>x"3200", 266=>x"3300", 267=>x"3600", 268=>x"2d00",
---- 269=>x"3000", 270=>x"2f00", 271=>x"3100", 272=>x"3100",
---- 273=>x"3400", 274=>x"2f00", 275=>x"3100", 276=>x"3300",
---- 277=>x"3200", 278=>x"3200", 279=>x"2e00", 280=>x"3600",
---- 281=>x"3300", 282=>x"3400", 283=>x"3200", 284=>x"3300",
---- 285=>x"3500", 286=>x"3500", 287=>x"3300", 288=>x"3300",
---- 289=>x"3800", 290=>x"3300", 291=>x"3300", 292=>x"2e00",
---- 293=>x"2e00", 294=>x"3100", 295=>x"3900", 296=>x"3200",
---- 297=>x"2d00", 298=>x"2e00", 299=>x"3400", 300=>x"2e00",
---- 301=>x"3000", 302=>x"3100", 303=>x"3400", 304=>x"2c00",
---- 305=>x"3300", 306=>x"3100", 307=>x"3800", 308=>x"3000",
---- 309=>x"3200", 310=>x"2e00", 311=>x"3400", 312=>x"2f00",
---- 313=>x"3500", 314=>x"3500", 315=>x"3300", 316=>x"3500",
---- 317=>x"3500", 318=>x"3200", 319=>x"2d00", 320=>x"4200",
---- 321=>x"3100", 322=>x"2d00", 323=>x"2800", 324=>x"3400",
---- 325=>x"d100", 326=>x"2b00", 327=>x"2a00", 328=>x"3100",
---- 329=>x"3800", 330=>x"2900", 331=>x"2900", 332=>x"3000",
---- 333=>x"2e00", 334=>x"3400", 335=>x"3300", 336=>x"3a00",
---- 337=>x"3000", 338=>x"3700", 339=>x"4200", 340=>x"3400",
---- 341=>x"3000", 342=>x"3100", 343=>x"4200", 344=>x"2e00",
---- 345=>x"2d00", 346=>x"3300", 347=>x"3a00", 348=>x"2c00",
---- 349=>x"3200", 350=>x"3500", 351=>x"3800", 352=>x"2a00",
---- 353=>x"3100", 354=>x"3600", 355=>x"3800", 356=>x"2b00",
---- 357=>x"3100", 358=>x"3800", 359=>x"3300", 360=>x"3300",
---- 361=>x"3600", 362=>x"3600", 363=>x"2e00", 364=>x"3300",
---- 365=>x"3900", 366=>x"2f00", 367=>x"2d00", 368=>x"3700",
---- 369=>x"3900", 370=>x"2f00", 371=>x"2800", 372=>x"3800",
---- 373=>x"3700", 374=>x"3100", 375=>x"2c00", 376=>x"3c00",
---- 377=>x"3c00", 378=>x"3300", 379=>x"3000", 380=>x"3700",
---- 381=>x"3d00", 382=>x"3c00", 383=>x"3400", 384=>x"3e00",
---- 385=>x"3500", 386=>x"3200", 387=>x"3f00", 388=>x"2a00",
---- 389=>x"2e00", 390=>x"2f00", 391=>x"5200", 392=>x"2b00",
---- 393=>x"3100", 394=>x"3500", 395=>x"6800", 396=>x"3300",
---- 397=>x"3200", 398=>x"4900", 399=>x"7900", 400=>x"3300",
---- 401=>x"3800", 402=>x"6000", 403=>x"8400", 404=>x"3400",
---- 405=>x"4500", 406=>x"6b00", 407=>x"8700", 408=>x"4200",
---- 409=>x"5000", 410=>x"7800", 411=>x"8a00", 412=>x"4700",
---- 413=>x"6200", 414=>x"8200", 415=>x"8900", 416=>x"4c00",
---- 417=>x"7400", 418=>x"8600", 419=>x"8500", 420=>x"5900",
---- 421=>x"7c00", 422=>x"8500", 423=>x"8000", 424=>x"7000",
---- 425=>x"8700", 426=>x"8500", 427=>x"7a00", 428=>x"7b00",
---- 429=>x"8800", 430=>x"8100", 431=>x"7a00", 432=>x"8400",
---- 433=>x"8900", 434=>x"8100", 435=>x"7a00", 436=>x"8d00",
---- 437=>x"8800", 438=>x"7e00", 439=>x"7e00", 440=>x"8e00",
---- 441=>x"8600", 442=>x"7f00", 443=>x"8800", 444=>x"8b00",
---- 445=>x"8200", 446=>x"8100", 447=>x"9300", 448=>x"8900",
---- 449=>x"7e00", 450=>x"8800", 451=>x"9900", 452=>x"8600",
---- 453=>x"8100", 454=>x"9000", 455=>x"a000", 456=>x"8300",
---- 457=>x"8900", 458=>x"9900", 459=>x"a300", 460=>x"8200",
---- 461=>x"8e00", 462=>x"9e00", 463=>x"a700", 464=>x"8400",
---- 465=>x"6c00", 466=>x"a200", 467=>x"a500", 468=>x"8900",
---- 469=>x"9a00", 470=>x"a500", 471=>x"a700", 472=>x"8f00",
---- 473=>x"9f00", 474=>x"a600", 475=>x"a300", 476=>x"9400",
---- 477=>x"a000", 478=>x"a500", 479=>x"a400", 480=>x"9a00",
---- 481=>x"a300", 482=>x"a200", 483=>x"a400", 484=>x"9d00",
---- 485=>x"a200", 486=>x"a300", 487=>x"a400", 488=>x"a000",
---- 489=>x"a000", 490=>x"a000", 491=>x"a000", 492=>x"a200",
---- 493=>x"a100", 494=>x"a000", 495=>x"9f00", 496=>x"a500",
---- 497=>x"a400", 498=>x"9f00", 499=>x"9f00", 500=>x"a100",
---- 501=>x"a200", 502=>x"9f00", 503=>x"9f00", 504=>x"a300",
---- 505=>x"a100", 506=>x"9f00", 507=>x"a000", 508=>x"a100",
---- 509=>x"9f00", 510=>x"9e00", 511=>x"9e00", 512=>x"9f00",
---- 513=>x"9f00", 514=>x"9e00", 515=>x"9b00", 516=>x"9f00",
---- 517=>x"9f00", 518=>x"9d00", 519=>x"9c00", 520=>x"9d00",
---- 521=>x"9c00", 522=>x"9d00", 523=>x"9a00", 524=>x"9d00",
---- 525=>x"9c00", 526=>x"9b00", 527=>x"6500", 528=>x"9d00",
---- 529=>x"9c00", 530=>x"9c00", 531=>x"6600", 532=>x"9d00",
---- 533=>x"9e00", 534=>x"9c00", 535=>x"9800", 536=>x"9c00",
---- 537=>x"9f00", 538=>x"9b00", 539=>x"9900", 540=>x"9b00",
---- 541=>x"9c00", 542=>x"9800", 543=>x"9900", 544=>x"9b00",
---- 545=>x"9a00", 546=>x"9a00", 547=>x"9900", 548=>x"9800",
---- 549=>x"9800", 550=>x"9900", 551=>x"9800", 552=>x"9800",
---- 553=>x"9700", 554=>x"9900", 555=>x"9400", 556=>x"9900",
---- 557=>x"9900", 558=>x"9900", 559=>x"9800", 560=>x"9a00",
---- 561=>x"9700", 562=>x"9800", 563=>x"9800", 564=>x"9800",
---- 565=>x"9500", 566=>x"9600", 567=>x"9600", 568=>x"9800",
---- 569=>x"9700", 570=>x"9500", 571=>x"6600", 572=>x"9800",
---- 573=>x"9700", 574=>x"9600", 575=>x"9600", 576=>x"9500",
---- 577=>x"9700", 578=>x"9700", 579=>x"9700", 580=>x"9900",
---- 581=>x"9a00", 582=>x"9800", 583=>x"9500", 584=>x"9700",
---- 585=>x"9700", 586=>x"9600", 587=>x"9600", 588=>x"9500",
---- 589=>x"9800", 590=>x"9900", 591=>x"9700", 592=>x"9600",
---- 593=>x"9700", 594=>x"9700", 595=>x"9600", 596=>x"9800",
---- 597=>x"6a00", 598=>x"9300", 599=>x"9700", 600=>x"9700",
---- 601=>x"9700", 602=>x"9700", 603=>x"9400", 604=>x"9800",
---- 605=>x"9500", 606=>x"9400", 607=>x"9500", 608=>x"9600",
---- 609=>x"9500", 610=>x"9400", 611=>x"9500", 612=>x"9800",
---- 613=>x"9700", 614=>x"9500", 615=>x"9600", 616=>x"9700",
---- 617=>x"9900", 618=>x"9600", 619=>x"9600", 620=>x"9600",
---- 621=>x"9700", 622=>x"9800", 623=>x"9600", 624=>x"9900",
---- 625=>x"9700", 626=>x"9700", 627=>x"9500", 628=>x"9800",
---- 629=>x"9800", 630=>x"9600", 631=>x"9400", 632=>x"9600",
---- 633=>x"9500", 634=>x"9600", 635=>x"9900", 636=>x"9700",
---- 637=>x"9600", 638=>x"9300", 639=>x"9400", 640=>x"9700",
---- 641=>x"9500", 642=>x"9500", 643=>x"9500", 644=>x"9700",
---- 645=>x"9600", 646=>x"9400", 647=>x"9000", 648=>x"9500",
---- 649=>x"9500", 650=>x"9300", 651=>x"9400", 652=>x"9600",
---- 653=>x"9400", 654=>x"9400", 655=>x"9500", 656=>x"9500",
---- 657=>x"9700", 658=>x"9500", 659=>x"9400", 660=>x"9300",
---- 661=>x"9400", 662=>x"9600", 663=>x"9300", 664=>x"9500",
---- 665=>x"9600", 666=>x"9300", 667=>x"9200", 668=>x"9500",
---- 669=>x"9300", 670=>x"9000", 671=>x"9400", 672=>x"9200",
---- 673=>x"9100", 674=>x"9100", 675=>x"9100", 676=>x"9300",
---- 677=>x"8e00", 678=>x"9000", 679=>x"9200", 680=>x"9100",
---- 681=>x"9100", 682=>x"9000", 683=>x"9200", 684=>x"9000",
---- 685=>x"9300", 686=>x"9400", 687=>x"9000", 688=>x"9300",
---- 689=>x"9400", 690=>x"9000", 691=>x"9200", 692=>x"9500",
---- 693=>x"9400", 694=>x"9000", 695=>x"9100", 696=>x"9400",
---- 697=>x"9300", 698=>x"9300", 699=>x"9100", 700=>x"9200",
---- 701=>x"9400", 702=>x"9500", 703=>x"6e00", 704=>x"9400",
---- 705=>x"9500", 706=>x"9200", 707=>x"9100", 708=>x"9400",
---- 709=>x"9300", 710=>x"9200", 711=>x"9200", 712=>x"9400",
---- 713=>x"9300", 714=>x"9100", 715=>x"9000", 716=>x"9300",
---- 717=>x"9200", 718=>x"9100", 719=>x"9000", 720=>x"9500",
---- 721=>x"9300", 722=>x"9100", 723=>x"9200", 724=>x"9600",
---- 725=>x"9200", 726=>x"9100", 727=>x"9100", 728=>x"9500",
---- 729=>x"9500", 730=>x"9200", 731=>x"9200", 732=>x"9500",
---- 733=>x"9400", 734=>x"9200", 735=>x"9100", 736=>x"9500",
---- 737=>x"9400", 738=>x"9200", 739=>x"9200", 740=>x"9400",
---- 741=>x"9400", 742=>x"9400", 743=>x"9100", 744=>x"9600",
---- 745=>x"9500", 746=>x"9000", 747=>x"9000", 748=>x"9600",
---- 749=>x"9500", 750=>x"6e00", 751=>x"8f00", 752=>x"9400",
---- 753=>x"9300", 754=>x"9000", 755=>x"8e00", 756=>x"9500",
---- 757=>x"9300", 758=>x"9000", 759=>x"8e00", 760=>x"9100",
---- 761=>x"8f00", 762=>x"8e00", 763=>x"8d00", 764=>x"9100",
---- 765=>x"8f00", 766=>x"8f00", 767=>x"8c00", 768=>x"9200",
---- 769=>x"9000", 770=>x"8f00", 771=>x"8d00", 772=>x"9000",
---- 773=>x"9100", 774=>x"8d00", 775=>x"7300", 776=>x"6f00",
---- 777=>x"8f00", 778=>x"8f00", 779=>x"8c00", 780=>x"8e00",
---- 781=>x"8c00", 782=>x"8c00", 783=>x"8c00", 784=>x"8500",
---- 785=>x"8600", 786=>x"8800", 787=>x"8900", 788=>x"7800",
---- 789=>x"7a00", 790=>x"7b00", 791=>x"7d00", 792=>x"7000",
---- 793=>x"7300", 794=>x"7000", 795=>x"7000", 796=>x"6400",
---- 797=>x"6900", 798=>x"6600", 799=>x"9b00", 800=>x"5f00",
---- 801=>x"6100", 802=>x"6000", 803=>x"5c00", 804=>x"6100",
---- 805=>x"5f00", 806=>x"5e00", 807=>x"5700", 808=>x"6800",
---- 809=>x"6b00", 810=>x"5f00", 811=>x"5800", 812=>x"7200",
---- 813=>x"6d00", 814=>x"6800", 815=>x"6100", 816=>x"7600",
---- 817=>x"7500", 818=>x"7400", 819=>x"9600", 820=>x"7b00",
---- 821=>x"7c00", 822=>x"7700", 823=>x"7100", 824=>x"7f00",
---- 825=>x"7f00", 826=>x"7800", 827=>x"7700", 828=>x"7f00",
---- 829=>x"7e00", 830=>x"7a00", 831=>x"7b00", 832=>x"7f00",
---- 833=>x"8000", 834=>x"7c00", 835=>x"7e00", 836=>x"8100",
---- 837=>x"7e00", 838=>x"8100", 839=>x"7f00", 840=>x"8100",
---- 841=>x"7e00", 842=>x"8200", 843=>x"7f00", 844=>x"8200",
---- 845=>x"8200", 846=>x"7e00", 847=>x"7b00", 848=>x"7f00",
---- 849=>x"7e00", 850=>x"7d00", 851=>x"7a00", 852=>x"7d00",
---- 853=>x"7b00", 854=>x"7b00", 855=>x"7900", 856=>x"7c00",
---- 857=>x"7e00", 858=>x"7a00", 859=>x"7f00", 860=>x"7a00",
---- 861=>x"7b00", 862=>x"7900", 863=>x"8b00", 864=>x"8000",
---- 865=>x"7800", 866=>x"7b00", 867=>x"9d00", 868=>x"7f00",
---- 869=>x"7700", 870=>x"8000", 871=>x"ae00", 872=>x"7900",
---- 873=>x"7700", 874=>x"8500", 875=>x"ba00", 876=>x"7800",
---- 877=>x"7800", 878=>x"6f00", 879=>x"c100", 880=>x"7a00",
---- 881=>x"7c00", 882=>x"9600", 883=>x"c400", 884=>x"7b00",
---- 885=>x"8200", 886=>x"9c00", 887=>x"c700", 888=>x"7f00",
---- 889=>x"8300", 890=>x"a300", 891=>x"ca00", 892=>x"7f00",
---- 893=>x"8200", 894=>x"a800", 895=>x"cb00", 896=>x"7e00",
---- 897=>x"8400", 898=>x"a200", 899=>x"c200", 900=>x"8100",
---- 901=>x"8400", 902=>x"9600", 903=>x"b800", 904=>x"8800",
---- 905=>x"8600", 906=>x"8a00", 907=>x"9d00", 908=>x"8c00",
---- 909=>x"8a00", 910=>x"8a00", 911=>x"8b00", 912=>x"8e00",
---- 913=>x"8d00", 914=>x"8c00", 915=>x"8a00", 916=>x"9400",
---- 917=>x"9200", 918=>x"8f00", 919=>x"8c00", 920=>x"9600",
---- 921=>x"9100", 922=>x"9000", 923=>x"8c00", 924=>x"9400",
---- 925=>x"8d00", 926=>x"8700", 927=>x"8300", 928=>x"9700",
---- 929=>x"8e00", 930=>x"7c00", 931=>x"7d00", 932=>x"9600",
---- 933=>x"8f00", 934=>x"9100", 935=>x"9200", 936=>x"9400",
---- 937=>x"a200", 938=>x"a700", 939=>x"9b00", 940=>x"ad00",
---- 941=>x"bc00", 942=>x"b400", 943=>x"a000", 944=>x"c300",
---- 945=>x"c300", 946=>x"bd00", 947=>x"a800", 948=>x"ca00",
---- 949=>x"ca00", 950=>x"bb00", 951=>x"9f00", 952=>x"ce00",
---- 953=>x"d000", 954=>x"b100", 955=>x"9400", 956=>x"cc00",
---- 957=>x"cb00", 958=>x"ae00", 959=>x"9f00", 960=>x"ca00",
---- 961=>x"c900", 962=>x"bd00", 963=>x"b800", 964=>x"c900",
---- 965=>x"ca00", 966=>x"ca00", 967=>x"c500", 968=>x"cd00",
---- 969=>x"d200", 970=>x"d100", 971=>x"c800", 972=>x"cd00",
---- 973=>x"d500", 974=>x"d000", 975=>x"bf00", 976=>x"ca00",
---- 977=>x"ce00", 978=>x"c300", 979=>x"ab00", 980=>x"b700",
---- 981=>x"b600", 982=>x"a700", 983=>x"7b00", 984=>x"9400",
---- 985=>x"8c00", 986=>x"7300", 987=>x"5800", 988=>x"7500",
---- 989=>x"6e00", 990=>x"6000", 991=>x"5700", 992=>x"6900",
---- 993=>x"6500", 994=>x"5f00", 995=>x"5b00", 996=>x"6700",
---- 997=>x"6600", 998=>x"6200", 999=>x"6000", 1000=>x"6a00",
---- 1001=>x"6800", 1002=>x"6500", 1003=>x"6200", 1004=>x"6b00",
---- 1005=>x"6b00", 1006=>x"6a00", 1007=>x"6e00", 1008=>x"6e00",
---- 1009=>x"7100", 1010=>x"7300", 1011=>x"7800", 1012=>x"7600",
---- 1013=>x"7500", 1014=>x"7b00", 1015=>x"7f00", 1016=>x"7d00",
---- 1017=>x"8200", 1018=>x"8700", 1019=>x"8500", 1020=>x"8400",
---- 1021=>x"8a00", 1022=>x"8b00", 1023=>x"8600"),
----
---- 54 => (0=>x"7300", 1=>x"7600", 2=>x"7600", 3=>x"7900", 4=>x"7300",
---- 5=>x"7600", 6=>x"7600", 7=>x"7900", 8=>x"7300",
---- 9=>x"7600", 10=>x"7600", 11=>x"7800", 12=>x"7100",
---- 13=>x"7400", 14=>x"7700", 15=>x"7600", 16=>x"6f00",
---- 17=>x"8f00", 18=>x"7500", 19=>x"7700", 20=>x"6a00",
---- 21=>x"6e00", 22=>x"7100", 23=>x"7300", 24=>x"6800",
---- 25=>x"6e00", 26=>x"7000", 27=>x"7300", 28=>x"6a00",
---- 29=>x"6d00", 30=>x"6e00", 31=>x"7000", 32=>x"6800",
---- 33=>x"6800", 34=>x"6c00", 35=>x"6e00", 36=>x"6d00",
---- 37=>x"6700", 38=>x"6900", 39=>x"9300", 40=>x"8600",
---- 41=>x"6600", 42=>x"6d00", 43=>x"6a00", 44=>x"a300",
---- 45=>x"7100", 46=>x"6900", 47=>x"6a00", 48=>x"c000",
---- 49=>x"9100", 50=>x"6700", 51=>x"6900", 52=>x"ce00",
---- 53=>x"b100", 54=>x"7800", 55=>x"6400", 56=>x"d500",
---- 57=>x"c700", 58=>x"9a00", 59=>x"6900", 60=>x"dc00",
---- 61=>x"d500", 62=>x"ba00", 63=>x"7f00", 64=>x"de00",
---- 65=>x"dc00", 66=>x"d100", 67=>x"b100", 68=>x"df00",
---- 69=>x"de00", 70=>x"d800", 71=>x"c300", 72=>x"de00",
---- 73=>x"e100", 74=>x"db00", 75=>x"cf00", 76=>x"de00",
---- 77=>x"df00", 78=>x"e100", 79=>x"d900", 80=>x"df00",
---- 81=>x"de00", 82=>x"e100", 83=>x"de00", 84=>x"dc00",
---- 85=>x"de00", 86=>x"2000", 87=>x"df00", 88=>x"da00",
---- 89=>x"dd00", 90=>x"df00", 91=>x"e100", 92=>x"d900",
---- 93=>x"dc00", 94=>x"e000", 95=>x"e000", 96=>x"d300",
---- 97=>x"da00", 98=>x"dc00", 99=>x"dc00", 100=>x"d000",
---- 101=>x"d700", 102=>x"d900", 103=>x"de00", 104=>x"c500",
---- 105=>x"d300", 106=>x"2700", 107=>x"db00", 108=>x"b400",
---- 109=>x"cd00", 110=>x"d600", 111=>x"dc00", 112=>x"9b00",
---- 113=>x"c200", 114=>x"d200", 115=>x"db00", 116=>x"8a00",
---- 117=>x"ac00", 118=>x"cd00", 119=>x"d700", 120=>x"7700",
---- 121=>x"9300", 122=>x"bd00", 123=>x"d000", 124=>x"8c00",
---- 125=>x"8b00", 126=>x"a500", 127=>x"c600", 128=>x"8d00",
---- 129=>x"8c00", 130=>x"9200", 131=>x"b300", 132=>x"8f00",
---- 133=>x"8f00", 134=>x"8e00", 135=>x"9900", 136=>x"9100",
---- 137=>x"9300", 138=>x"9300", 139=>x"9100", 140=>x"9200",
---- 141=>x"9400", 142=>x"9800", 143=>x"9600", 144=>x"9400",
---- 145=>x"6b00", 146=>x"9900", 147=>x"9a00", 148=>x"9600",
---- 149=>x"9600", 150=>x"9900", 151=>x"9e00", 152=>x"9600",
---- 153=>x"9900", 154=>x"9c00", 155=>x"9d00", 156=>x"9900",
---- 157=>x"9b00", 158=>x"9e00", 159=>x"8b00", 160=>x"9a00",
---- 161=>x"9d00", 162=>x"9100", 163=>x"6700", 164=>x"9d00",
---- 165=>x"9800", 166=>x"7500", 167=>x"3d00", 168=>x"9b00",
---- 169=>x"8400", 170=>x"4e00", 171=>x"2c00", 172=>x"9200",
---- 173=>x"5d00", 174=>x"2d00", 175=>x"2500", 176=>x"7100",
---- 177=>x"3700", 178=>x"2800", 179=>x"2700", 180=>x"4500",
---- 181=>x"2900", 182=>x"3c00", 183=>x"4100", 184=>x"2e00",
---- 185=>x"2e00", 186=>x"3500", 187=>x"3500", 188=>x"2700",
---- 189=>x"2600", 190=>x"2900", 191=>x"2b00", 192=>x"2700",
---- 193=>x"2400", 194=>x"2c00", 195=>x"2b00", 196=>x"2700",
---- 197=>x"2700", 198=>x"2800", 199=>x"2e00", 200=>x"2600",
---- 201=>x"2800", 202=>x"2b00", 203=>x"2d00", 204=>x"2900",
---- 205=>x"2900", 206=>x"2f00", 207=>x"2f00", 208=>x"2d00",
---- 209=>x"2f00", 210=>x"3000", 211=>x"3200", 212=>x"2c00",
---- 213=>x"2e00", 214=>x"3300", 215=>x"3700", 216=>x"ce00",
---- 217=>x"2f00", 218=>x"3500", 219=>x"3400", 220=>x"3300",
---- 221=>x"3500", 222=>x"3c00", 223=>x"3600", 224=>x"3400",
---- 225=>x"3500", 226=>x"3900", 227=>x"3600", 228=>x"3a00",
---- 229=>x"3500", 230=>x"3500", 231=>x"3400", 232=>x"3a00",
---- 233=>x"3900", 234=>x"3400", 235=>x"c500", 236=>x"3700",
---- 237=>x"3400", 238=>x"3200", 239=>x"3b00", 240=>x"3800",
---- 241=>x"3600", 242=>x"3700", 243=>x"3600", 244=>x"3600",
---- 245=>x"3800", 246=>x"3a00", 247=>x"3100", 248=>x"3500",
---- 249=>x"3500", 250=>x"3500", 251=>x"3300", 252=>x"3400",
---- 253=>x"3400", 254=>x"3800", 255=>x"3100", 256=>x"3400",
---- 257=>x"3100", 258=>x"2f00", 259=>x"2b00", 260=>x"3a00",
---- 261=>x"2f00", 262=>x"2f00", 263=>x"2d00", 264=>x"3a00",
---- 265=>x"2f00", 266=>x"3200", 267=>x"3000", 268=>x"3900",
---- 269=>x"3700", 270=>x"3900", 271=>x"3200", 272=>x"3300",
---- 273=>x"3400", 274=>x"3500", 275=>x"3000", 276=>x"3200",
---- 277=>x"3200", 278=>x"3500", 279=>x"3000", 280=>x"3300",
---- 281=>x"3200", 282=>x"2e00", 283=>x"2f00", 284=>x"3400",
---- 285=>x"3100", 286=>x"2e00", 287=>x"2800", 288=>x"3800",
---- 289=>x"3100", 290=>x"2f00", 291=>x"2c00", 292=>x"3800",
---- 293=>x"3200", 294=>x"2e00", 295=>x"2800", 296=>x"2f00",
---- 297=>x"2d00", 298=>x"2b00", 299=>x"2d00", 300=>x"3300",
---- 301=>x"2e00", 302=>x"2a00", 303=>x"3000", 304=>x"3f00",
---- 305=>x"2d00", 306=>x"2e00", 307=>x"2f00", 308=>x"3200",
---- 309=>x"2d00", 310=>x"2e00", 311=>x"3000", 312=>x"2d00",
---- 313=>x"2a00", 314=>x"d100", 315=>x"d000", 316=>x"2c00",
---- 317=>x"2b00", 318=>x"3200", 319=>x"2f00", 320=>x"2d00",
---- 321=>x"3200", 322=>x"3300", 323=>x"2d00", 324=>x"3100",
---- 325=>x"3500", 326=>x"3200", 327=>x"2e00", 328=>x"3000",
---- 329=>x"3500", 330=>x"2f00", 331=>x"2e00", 332=>x"3400",
---- 333=>x"3600", 334=>x"3000", 335=>x"3400", 336=>x"3a00",
---- 337=>x"3500", 338=>x"3200", 339=>x"3300", 340=>x"3a00",
---- 341=>x"3400", 342=>x"3500", 343=>x"3800", 344=>x"3200",
---- 345=>x"3500", 346=>x"3800", 347=>x"3b00", 348=>x"3400",
---- 349=>x"3200", 350=>x"3600", 351=>x"4100", 352=>x"3500",
---- 353=>x"3000", 354=>x"3900", 355=>x"5600", 356=>x"2d00",
---- 357=>x"2e00", 358=>x"4300", 359=>x"6b00", 360=>x"2900",
---- 361=>x"2c00", 362=>x"5100", 363=>x"8000", 364=>x"2900",
---- 365=>x"3400", 366=>x"6200", 367=>x"8c00", 368=>x"2500",
---- 369=>x"4400", 370=>x"7900", 371=>x"6b00", 372=>x"3200",
---- 373=>x"5d00", 374=>x"8700", 375=>x"9500", 376=>x"4300",
---- 377=>x"7300", 378=>x"9000", 379=>x"9600", 380=>x"5800",
---- 381=>x"8600", 382=>x"9500", 383=>x"9600", 384=>x"7100",
---- 385=>x"8f00", 386=>x"9600", 387=>x"9400", 388=>x"8000",
---- 389=>x"9400", 390=>x"9300", 391=>x"9300", 392=>x"8f00",
---- 393=>x"9700", 394=>x"9200", 395=>x"9100", 396=>x"9200",
---- 397=>x"9300", 398=>x"8f00", 399=>x"8e00", 400=>x"9000",
---- 401=>x"9100", 402=>x"8c00", 403=>x"8d00", 404=>x"8a00",
---- 405=>x"8a00", 406=>x"8700", 407=>x"8f00", 408=>x"8400",
---- 409=>x"8400", 410=>x"8200", 411=>x"9600", 412=>x"7f00",
---- 413=>x"7b00", 414=>x"8600", 415=>x"9d00", 416=>x"7c00",
---- 417=>x"7c00", 418=>x"8e00", 419=>x"a300", 420=>x"7b00",
---- 421=>x"8000", 422=>x"9400", 423=>x"a500", 424=>x"7a00",
---- 425=>x"8600", 426=>x"9900", 427=>x"a500", 428=>x"7c00",
---- 429=>x"8e00", 430=>x"9b00", 431=>x"a200", 432=>x"8100",
---- 433=>x"9600", 434=>x"a000", 435=>x"a100", 436=>x"8c00",
---- 437=>x"9a00", 438=>x"9b00", 439=>x"9e00", 440=>x"6c00",
---- 441=>x"6600", 442=>x"9600", 443=>x"9600", 444=>x"9a00",
---- 445=>x"9800", 446=>x"9700", 447=>x"9600", 448=>x"a100",
---- 449=>x"9b00", 450=>x"9800", 451=>x"9700", 452=>x"a200",
---- 453=>x"9d00", 454=>x"9900", 455=>x"9800", 456=>x"a300",
---- 457=>x"9e00", 458=>x"9a00", 459=>x"9a00", 460=>x"a500",
---- 461=>x"a100", 462=>x"9f00", 463=>x"9c00", 464=>x"a400",
---- 465=>x"a300", 466=>x"a400", 467=>x"a200", 468=>x"a500",
---- 469=>x"a200", 470=>x"a300", 471=>x"a200", 472=>x"a000",
---- 473=>x"a200", 474=>x"a200", 475=>x"a400", 476=>x"a100",
---- 477=>x"a200", 478=>x"a100", 479=>x"a000", 480=>x"a200",
---- 481=>x"a300", 482=>x"a200", 483=>x"a100", 484=>x"a300",
---- 485=>x"a200", 486=>x"a100", 487=>x"9f00", 488=>x"a000",
---- 489=>x"a100", 490=>x"a000", 491=>x"a000", 492=>x"6000",
---- 493=>x"9d00", 494=>x"9e00", 495=>x"9f00", 496=>x"9e00",
---- 497=>x"9d00", 498=>x"9e00", 499=>x"9f00", 500=>x"9d00",
---- 501=>x"9d00", 502=>x"9e00", 503=>x"9e00", 504=>x"9e00",
---- 505=>x"9c00", 506=>x"9c00", 507=>x"9d00", 508=>x"9d00",
---- 509=>x"9b00", 510=>x"9c00", 511=>x"9d00", 512=>x"9c00",
---- 513=>x"9c00", 514=>x"9d00", 515=>x"9c00", 516=>x"9b00",
---- 517=>x"9b00", 518=>x"9b00", 519=>x"9b00", 520=>x"9b00",
---- 521=>x"6500", 522=>x"9900", 523=>x"9800", 524=>x"9900",
---- 525=>x"9800", 526=>x"9800", 527=>x"9a00", 528=>x"9a00",
---- 529=>x"9d00", 530=>x"9800", 531=>x"9900", 532=>x"9800",
---- 533=>x"9900", 534=>x"9900", 535=>x"9800", 536=>x"6600",
---- 537=>x"6800", 538=>x"9800", 539=>x"9700", 540=>x"9800",
---- 541=>x"9700", 542=>x"9900", 543=>x"9700", 544=>x"9700",
---- 545=>x"9900", 546=>x"9800", 547=>x"9800", 548=>x"6a00",
---- 549=>x"9700", 550=>x"9800", 551=>x"9900", 552=>x"9300",
---- 553=>x"9700", 554=>x"9800", 555=>x"9800", 556=>x"9600",
---- 557=>x"9500", 558=>x"9600", 559=>x"9700", 560=>x"9800",
---- 561=>x"9700", 562=>x"9700", 563=>x"9800", 564=>x"9800",
---- 565=>x"9600", 566=>x"9700", 567=>x"9700", 568=>x"9800",
---- 569=>x"9700", 570=>x"9800", 571=>x"9700", 572=>x"9600",
---- 573=>x"9800", 574=>x"9800", 575=>x"9600", 576=>x"9500",
---- 577=>x"9800", 578=>x"9900", 579=>x"9700", 580=>x"9900",
---- 581=>x"9900", 582=>x"9700", 583=>x"9800", 584=>x"9600",
---- 585=>x"9600", 586=>x"9900", 587=>x"9900", 588=>x"9600",
---- 589=>x"9600", 590=>x"9700", 591=>x"9500", 592=>x"9500",
---- 593=>x"9500", 594=>x"9600", 595=>x"9500", 596=>x"9600",
---- 597=>x"6900", 598=>x"9300", 599=>x"9200", 600=>x"9300",
---- 601=>x"9600", 602=>x"9300", 603=>x"9100", 604=>x"9400",
---- 605=>x"9300", 606=>x"9200", 607=>x"9300", 608=>x"9400",
---- 609=>x"9000", 610=>x"9200", 611=>x"9200", 612=>x"9300",
---- 613=>x"9200", 614=>x"9300", 615=>x"9100", 616=>x"9400",
---- 617=>x"9400", 618=>x"9300", 619=>x"9400", 620=>x"9300",
---- 621=>x"9300", 622=>x"9400", 623=>x"9300", 624=>x"9600",
---- 625=>x"9400", 626=>x"9600", 627=>x"9300", 628=>x"9400",
---- 629=>x"9200", 630=>x"9400", 631=>x"9400", 632=>x"9700",
---- 633=>x"9500", 634=>x"9400", 635=>x"9400", 636=>x"9600",
---- 637=>x"9500", 638=>x"9200", 639=>x"9400", 640=>x"9300",
---- 641=>x"9500", 642=>x"9500", 643=>x"6a00", 644=>x"9300",
---- 645=>x"9300", 646=>x"9400", 647=>x"9000", 648=>x"9400",
---- 649=>x"9100", 650=>x"9100", 651=>x"9000", 652=>x"9300",
---- 653=>x"9100", 654=>x"6d00", 655=>x"8f00", 656=>x"9200",
---- 657=>x"9100", 658=>x"9300", 659=>x"9000", 660=>x"9200",
---- 661=>x"9400", 662=>x"9100", 663=>x"9100", 664=>x"9200",
---- 665=>x"9300", 666=>x"9200", 667=>x"9100", 668=>x"9300",
---- 669=>x"9300", 670=>x"9400", 671=>x"9100", 672=>x"9300",
---- 673=>x"9100", 674=>x"9000", 675=>x"9300", 676=>x"8f00",
---- 677=>x"9100", 678=>x"9200", 679=>x"9000", 680=>x"9100",
---- 681=>x"6e00", 682=>x"9200", 683=>x"9000", 684=>x"9100",
---- 685=>x"9200", 686=>x"9000", 687=>x"9100", 688=>x"8f00",
---- 689=>x"9200", 690=>x"9100", 691=>x"9000", 692=>x"9200",
---- 693=>x"9000", 694=>x"9000", 695=>x"8f00", 696=>x"9100",
---- 697=>x"9000", 698=>x"9000", 699=>x"8f00", 700=>x"8f00",
---- 701=>x"8f00", 702=>x"9000", 703=>x"9000", 704=>x"8f00",
---- 705=>x"9100", 706=>x"9100", 707=>x"9000", 708=>x"9000",
---- 709=>x"9200", 710=>x"9000", 711=>x"6d00", 712=>x"9200",
---- 713=>x"9400", 714=>x"8f00", 715=>x"9100", 716=>x"9300",
---- 717=>x"9200", 718=>x"8d00", 719=>x"9000", 720=>x"9300",
---- 721=>x"9000", 722=>x"9100", 723=>x"9100", 724=>x"6e00",
---- 725=>x"8f00", 726=>x"8e00", 727=>x"8c00", 728=>x"9000",
---- 729=>x"8f00", 730=>x"8d00", 731=>x"8d00", 732=>x"8f00",
---- 733=>x"9000", 734=>x"8f00", 735=>x"8e00", 736=>x"9000",
---- 737=>x"8d00", 738=>x"8e00", 739=>x"8d00", 740=>x"9300",
---- 741=>x"8f00", 742=>x"8e00", 743=>x"8c00", 744=>x"8f00",
---- 745=>x"8e00", 746=>x"8c00", 747=>x"8b00", 748=>x"8e00",
---- 749=>x"8d00", 750=>x"8c00", 751=>x"8d00", 752=>x"8e00",
---- 753=>x"8c00", 754=>x"8c00", 755=>x"8800", 756=>x"8d00",
---- 757=>x"8b00", 758=>x"8c00", 759=>x"8b00", 760=>x"8c00",
---- 761=>x"8800", 762=>x"8a00", 763=>x"8900", 764=>x"8a00",
---- 765=>x"8b00", 766=>x"8900", 767=>x"8900", 768=>x"8d00",
---- 769=>x"8b00", 770=>x"8700", 771=>x"8700", 772=>x"8d00",
---- 773=>x"8800", 774=>x"8500", 775=>x"8500", 776=>x"8900",
---- 777=>x"8700", 778=>x"8700", 779=>x"8300", 780=>x"8900",
---- 781=>x"8a00", 782=>x"8700", 783=>x"8100", 784=>x"8700",
---- 785=>x"8700", 786=>x"8600", 787=>x"8200", 788=>x"8100",
---- 789=>x"8000", 790=>x"8100", 791=>x"7f00", 792=>x"7300",
---- 793=>x"7300", 794=>x"7400", 795=>x"7300", 796=>x"9900",
---- 797=>x"6800", 798=>x"6a00", 799=>x"6d00", 800=>x"5f00",
---- 801=>x"6000", 802=>x"6c00", 803=>x"6f00", 804=>x"5b00",
---- 805=>x"6400", 806=>x"7600", 807=>x"7700", 808=>x"6200",
---- 809=>x"6d00", 810=>x"7f00", 811=>x"8000", 812=>x"6400",
---- 813=>x"7400", 814=>x"8100", 815=>x"8600", 816=>x"6b00",
---- 817=>x"7600", 818=>x"8300", 819=>x"8700", 820=>x"7100",
---- 821=>x"7c00", 822=>x"8100", 823=>x"8300", 824=>x"7500",
---- 825=>x"7c00", 826=>x"7e00", 827=>x"8500", 828=>x"7900",
---- 829=>x"7c00", 830=>x"8500", 831=>x"8400", 832=>x"7d00",
---- 833=>x"8300", 834=>x"8900", 835=>x"8900", 836=>x"7e00",
---- 837=>x"8700", 838=>x"8a00", 839=>x"8b00", 840=>x"7d00",
---- 841=>x"8400", 842=>x"8700", 843=>x"8900", 844=>x"7900",
---- 845=>x"7d00", 846=>x"8b00", 847=>x"9700", 848=>x"7a00",
---- 849=>x"8600", 850=>x"9800", 851=>x"a500", 852=>x"8200",
---- 853=>x"9900", 854=>x"aa00", 855=>x"b800", 856=>x"9600",
---- 857=>x"ad00", 858=>x"bc00", 859=>x"c600", 860=>x"ae00",
---- 861=>x"c300", 862=>x"ca00", 863=>x"cb00", 864=>x"c100",
---- 865=>x"2f00", 866=>x"d400", 867=>x"d200", 868=>x"ce00",
---- 869=>x"d600", 870=>x"d900", 871=>x"d800", 872=>x"d300",
---- 873=>x"d900", 874=>x"db00", 875=>x"d700", 876=>x"d300",
---- 877=>x"da00", 878=>x"d900", 879=>x"d500", 880=>x"d500",
---- 881=>x"d800", 882=>x"d600", 883=>x"d000", 884=>x"d400",
---- 885=>x"d700", 886=>x"d300", 887=>x"cd00", 888=>x"d400",
---- 889=>x"d700", 890=>x"d300", 891=>x"cd00", 892=>x"d300",
---- 893=>x"d900", 894=>x"d200", 895=>x"ca00", 896=>x"d000",
---- 897=>x"d500", 898=>x"d100", 899=>x"cb00", 900=>x"c900",
---- 901=>x"cd00", 902=>x"cc00", 903=>x"ca00", 904=>x"b600",
---- 905=>x"bf00", 906=>x"bf00", 907=>x"c100", 908=>x"9700",
---- 909=>x"a600", 910=>x"a900", 911=>x"b300", 912=>x"8500",
---- 913=>x"8c00", 914=>x"9500", 915=>x"b100", 916=>x"8400",
---- 917=>x"8700", 918=>x"9400", 919=>x"b600", 920=>x"8700",
---- 921=>x"8b00", 922=>x"9900", 923=>x"be00", 924=>x"8500",
---- 925=>x"8d00", 926=>x"a600", 927=>x"3700", 928=>x"8100",
---- 929=>x"9200", 930=>x"b600", 931=>x"cf00", 932=>x"8c00",
---- 933=>x"9600", 934=>x"bc00", 935=>x"d300", 936=>x"9500",
---- 937=>x"a400", 938=>x"c400", 939=>x"d500", 940=>x"9700",
---- 941=>x"b300", 942=>x"cb00", 943=>x"d700", 944=>x"a000",
---- 945=>x"4700", 946=>x"ce00", 947=>x"d600", 948=>x"a000",
---- 949=>x"c100", 950=>x"d100", 951=>x"d800", 952=>x"ab00",
---- 953=>x"c800", 954=>x"d300", 955=>x"d600", 956=>x"b600",
---- 957=>x"c800", 958=>x"cf00", 959=>x"cf00", 960=>x"be00",
---- 961=>x"c800", 962=>x"c800", 963=>x"bf00", 964=>x"bf00",
---- 965=>x"ba00", 966=>x"b200", 967=>x"9f00", 968=>x"b800",
---- 969=>x"a200", 970=>x"8f00", 971=>x"7200", 972=>x"a100",
---- 973=>x"8000", 974=>x"5d00", 975=>x"4b00", 976=>x"7a00",
---- 977=>x"a800", 978=>x"4c00", 979=>x"4700", 980=>x"5700",
---- 981=>x"5000", 982=>x"5500", 983=>x"5000", 984=>x"5200",
---- 985=>x"4c00", 986=>x"4c00", 987=>x"4c00", 988=>x"5500",
---- 989=>x"5500", 990=>x"5400", 991=>x"5900", 992=>x"5b00",
---- 993=>x"9f00", 994=>x"6000", 995=>x"6400", 996=>x"6000",
---- 997=>x"6900", 998=>x"9300", 999=>x"6800", 1000=>x"6b00",
---- 1001=>x"7100", 1002=>x"7100", 1003=>x"6a00", 1004=>x"7400",
---- 1005=>x"7600", 1006=>x"7200", 1007=>x"6b00", 1008=>x"7d00",
---- 1009=>x"7a00", 1010=>x"7200", 1011=>x"9600", 1012=>x"8100",
---- 1013=>x"7b00", 1014=>x"7000", 1015=>x"6600", 1016=>x"7d00",
---- 1017=>x"7700", 1018=>x"6f00", 1019=>x"6100", 1020=>x"7d00",
---- 1021=>x"7400", 1022=>x"6500", 1023=>x"5900"),
----
---- 55 => (0=>x"8100", 1=>x"7600", 2=>x"7900", 3=>x"7900", 4=>x"7d00",
---- 5=>x"7600", 6=>x"7900", 7=>x"7900", 8=>x"7d00",
---- 9=>x"7600", 10=>x"7800", 11=>x"7b00", 12=>x"7700",
---- 13=>x"7900", 14=>x"8800", 15=>x"7b00", 16=>x"7700",
---- 17=>x"7800", 18=>x"7700", 19=>x"7a00", 20=>x"7a00",
---- 21=>x"8800", 22=>x"7700", 23=>x"7900", 24=>x"7500",
---- 25=>x"7a00", 26=>x"7700", 27=>x"7800", 28=>x"7500",
---- 29=>x"7500", 30=>x"7400", 31=>x"7600", 32=>x"7600",
---- 33=>x"7400", 34=>x"7400", 35=>x"7800", 36=>x"7100",
---- 37=>x"7400", 38=>x"7500", 39=>x"7700", 40=>x"7000",
---- 41=>x"7000", 42=>x"7200", 43=>x"7600", 44=>x"6f00",
---- 45=>x"7100", 46=>x"7300", 47=>x"7500", 48=>x"6d00",
---- 49=>x"6f00", 50=>x"7400", 51=>x"7800", 52=>x"6b00",
---- 53=>x"6f00", 54=>x"7300", 55=>x"7200", 56=>x"6900",
---- 57=>x"6d00", 58=>x"7200", 59=>x"7200", 60=>x"6500",
---- 61=>x"6d00", 62=>x"6f00", 63=>x"7400", 64=>x"7c00",
---- 65=>x"6d00", 66=>x"6e00", 67=>x"7000", 68=>x"9000",
---- 69=>x"6800", 70=>x"6900", 71=>x"6b00", 72=>x"b300",
---- 73=>x"7a00", 74=>x"6400", 75=>x"6800", 76=>x"ca00",
---- 77=>x"9c00", 78=>x"6700", 79=>x"6000", 80=>x"d400",
---- 81=>x"bc00", 82=>x"8400", 83=>x"6200", 84=>x"db00",
---- 85=>x"ca00", 86=>x"a300", 87=>x"6c00", 88=>x"df00",
---- 89=>x"d400", 90=>x"bf00", 91=>x"8600", 92=>x"e000",
---- 93=>x"db00", 94=>x"cf00", 95=>x"ab00", 96=>x"df00",
---- 97=>x"2000", 98=>x"d800", 99=>x"c600", 100=>x"e000",
---- 101=>x"e200", 102=>x"df00", 103=>x"d300", 104=>x"df00",
---- 105=>x"e200", 106=>x"e300", 107=>x"dd00", 108=>x"df00",
---- 109=>x"e000", 110=>x"1c00", 111=>x"e200", 112=>x"df00",
---- 113=>x"e000", 114=>x"e200", 115=>x"e400", 116=>x"dd00",
---- 117=>x"df00", 118=>x"e200", 119=>x"e300", 120=>x"d900",
---- 121=>x"dd00", 122=>x"e200", 123=>x"e400", 124=>x"d500",
---- 125=>x"dc00", 126=>x"e100", 127=>x"e500", 128=>x"d300",
---- 129=>x"dc00", 130=>x"e400", 131=>x"e600", 132=>x"c500",
---- 133=>x"da00", 134=>x"e100", 135=>x"e000", 136=>x"ae00",
---- 137=>x"d200", 138=>x"db00", 139=>x"d100", 140=>x"a300",
---- 141=>x"c900", 142=>x"c400", 143=>x"8500", 144=>x"a000",
---- 145=>x"a300", 146=>x"7500", 147=>x"3600", 148=>x"9900",
---- 149=>x"6f00", 150=>x"3900", 151=>x"2d00", 152=>x"8300",
---- 153=>x"4700", 154=>x"2900", 155=>x"2d00", 156=>x"5800",
---- 157=>x"3200", 158=>x"2a00", 159=>x"2b00", 160=>x"3000",
---- 161=>x"2e00", 162=>x"2c00", 163=>x"2e00", 164=>x"2900",
---- 165=>x"2c00", 166=>x"2800", 167=>x"2b00", 168=>x"2b00",
---- 169=>x"2600", 170=>x"2500", 171=>x"2a00", 172=>x"2700",
---- 173=>x"2900", 174=>x"2800", 175=>x"d600", 176=>x"2b00",
---- 177=>x"2a00", 178=>x"2b00", 179=>x"2d00", 180=>x"3700",
---- 181=>x"2c00", 182=>x"2a00", 183=>x"3300", 184=>x"2f00",
---- 185=>x"d200", 186=>x"2c00", 187=>x"3300", 188=>x"2a00",
---- 189=>x"2f00", 190=>x"3200", 191=>x"3600", 192=>x"3000",
---- 193=>x"3400", 194=>x"3900", 195=>x"3800", 196=>x"3200",
---- 197=>x"3b00", 198=>x"3a00", 199=>x"3800", 200=>x"3500",
---- 201=>x"3600", 202=>x"3900", 203=>x"3a00", 204=>x"3600",
---- 205=>x"3a00", 206=>x"3500", 207=>x"3400", 208=>x"3600",
---- 209=>x"3700", 210=>x"3300", 211=>x"3300", 212=>x"3600",
---- 213=>x"3500", 214=>x"3b00", 215=>x"3500", 216=>x"3400",
---- 217=>x"3700", 218=>x"3700", 219=>x"3300", 220=>x"2e00",
---- 221=>x"3600", 222=>x"3600", 223=>x"3600", 224=>x"3200",
---- 225=>x"3700", 226=>x"3a00", 227=>x"3b00", 228=>x"3400",
---- 229=>x"3800", 230=>x"3f00", 231=>x"c700", 232=>x"3900",
---- 233=>x"3200", 234=>x"3200", 235=>x"3300", 236=>x"3e00",
---- 237=>x"3600", 238=>x"3400", 239=>x"3200", 240=>x"3300",
---- 241=>x"3100", 242=>x"2e00", 243=>x"3000", 244=>x"3300",
---- 245=>x"2f00", 246=>x"3000", 247=>x"3600", 248=>x"3200",
---- 249=>x"3100", 250=>x"3200", 251=>x"3100", 252=>x"2c00",
---- 253=>x"3000", 254=>x"3100", 255=>x"2e00", 256=>x"2c00",
---- 257=>x"3200", 258=>x"2f00", 259=>x"2c00", 260=>x"2b00",
---- 261=>x"2d00", 262=>x"2c00", 263=>x"2e00", 264=>x"2f00",
---- 265=>x"2f00", 266=>x"2b00", 267=>x"2e00", 268=>x"2f00",
---- 269=>x"2f00", 270=>x"3100", 271=>x"3500", 272=>x"2b00",
---- 273=>x"2b00", 274=>x"2b00", 275=>x"3300", 276=>x"2c00",
---- 277=>x"2e00", 278=>x"2900", 279=>x"3000", 280=>x"2900",
---- 281=>x"2a00", 282=>x"2c00", 283=>x"3200", 284=>x"2900",
---- 285=>x"3100", 286=>x"3100", 287=>x"3400", 288=>x"2e00",
---- 289=>x"3200", 290=>x"2f00", 291=>x"3200", 292=>x"2e00",
---- 293=>x"3100", 294=>x"2e00", 295=>x"3400", 296=>x"2e00",
---- 297=>x"3500", 298=>x"3700", 299=>x"3600", 300=>x"2d00",
---- 301=>x"3700", 302=>x"3900", 303=>x"3100", 304=>x"3300",
---- 305=>x"3800", 306=>x"3900", 307=>x"2d00", 308=>x"3100",
---- 309=>x"3100", 310=>x"3500", 311=>x"3100", 312=>x"2a00",
---- 313=>x"2d00", 314=>x"3900", 315=>x"4300", 316=>x"2c00",
---- 317=>x"3200", 318=>x"4400", 319=>x"5100", 320=>x"2f00",
---- 321=>x"3900", 322=>x"4700", 323=>x"5b00", 324=>x"3100",
---- 325=>x"4200", 326=>x"4b00", 327=>x"6a00", 328=>x"3800",
---- 329=>x"4400", 330=>x"5b00", 331=>x"7f00", 332=>x"4000",
---- 333=>x"4700", 334=>x"6c00", 335=>x"9000", 336=>x"3d00",
---- 337=>x"5800", 338=>x"8100", 339=>x"9800", 340=>x"4200",
---- 341=>x"6b00", 342=>x"9000", 343=>x"9b00", 344=>x"5600",
---- 345=>x"7f00", 346=>x"9800", 347=>x"9a00", 348=>x"6900",
---- 349=>x"8d00", 350=>x"9700", 351=>x"9800", 352=>x"7c00",
---- 353=>x"9600", 354=>x"9700", 355=>x"9300", 356=>x"8e00",
---- 357=>x"9900", 358=>x"9600", 359=>x"9100", 360=>x"9500",
---- 361=>x"9500", 362=>x"9100", 363=>x"8e00", 364=>x"9500",
---- 365=>x"9300", 366=>x"8f00", 367=>x"8f00", 368=>x"6800",
---- 369=>x"9100", 370=>x"9000", 371=>x"9300", 372=>x"9700",
---- 373=>x"8f00", 374=>x"8e00", 375=>x"9700", 376=>x"9500",
---- 377=>x"8e00", 378=>x"9300", 379=>x"9e00", 380=>x"9300",
---- 381=>x"8e00", 382=>x"9700", 383=>x"a100", 384=>x"9000",
---- 385=>x"9000", 386=>x"9d00", 387=>x"a400", 388=>x"8b00",
---- 389=>x"9200", 390=>x"a200", 391=>x"a500", 392=>x"8f00",
---- 393=>x"9b00", 394=>x"a400", 395=>x"a700", 396=>x"9400",
---- 397=>x"a000", 398=>x"a500", 399=>x"a400", 400=>x"9a00",
---- 401=>x"a400", 402=>x"a600", 403=>x"a800", 404=>x"a000",
---- 405=>x"a600", 406=>x"a600", 407=>x"a700", 408=>x"a500",
---- 409=>x"a600", 410=>x"a500", 411=>x"a700", 412=>x"a700",
---- 413=>x"a700", 414=>x"a700", 415=>x"a700", 416=>x"a800",
---- 417=>x"a900", 418=>x"a800", 419=>x"a700", 420=>x"a900",
---- 421=>x"a700", 422=>x"a700", 423=>x"a700", 424=>x"a700",
---- 425=>x"a500", 426=>x"a700", 427=>x"a500", 428=>x"a600",
---- 429=>x"a700", 430=>x"a600", 431=>x"a500", 432=>x"a300",
---- 433=>x"a600", 434=>x"a400", 435=>x"a500", 436=>x"a100",
---- 437=>x"a500", 438=>x"a700", 439=>x"a500", 440=>x"9b00",
---- 441=>x"a000", 442=>x"a400", 443=>x"a400", 444=>x"9800",
---- 445=>x"9800", 446=>x"9b00", 447=>x"a000", 448=>x"9800",
---- 449=>x"9600", 450=>x"9500", 451=>x"9900", 452=>x"9800",
---- 453=>x"9600", 454=>x"9600", 455=>x"9500", 456=>x"9b00",
---- 457=>x"9700", 458=>x"9900", 459=>x"6700", 460=>x"9b00",
---- 461=>x"9900", 462=>x"9800", 463=>x"9800", 464=>x"a000",
---- 465=>x"9d00", 466=>x"9900", 467=>x"9800", 468=>x"a100",
---- 469=>x"9f00", 470=>x"9d00", 471=>x"a000", 472=>x"a000",
---- 473=>x"9e00", 474=>x"a300", 475=>x"a500", 476=>x"9f00",
---- 477=>x"a000", 478=>x"a200", 479=>x"a400", 480=>x"a100",
---- 481=>x"a000", 482=>x"a100", 483=>x"a500", 484=>x"9f00",
---- 485=>x"a000", 486=>x"a100", 487=>x"a200", 488=>x"9f00",
---- 489=>x"a000", 490=>x"a000", 491=>x"a000", 492=>x"9f00",
---- 493=>x"9d00", 494=>x"9d00", 495=>x"9f00", 496=>x"9c00",
---- 497=>x"9d00", 498=>x"9c00", 499=>x"a000", 500=>x"9e00",
---- 501=>x"9e00", 502=>x"6400", 503=>x"9b00", 504=>x"9d00",
---- 505=>x"6400", 506=>x"9b00", 507=>x"9c00", 508=>x"9c00",
---- 509=>x"9c00", 510=>x"9b00", 511=>x"9a00", 512=>x"9d00",
---- 513=>x"9b00", 514=>x"9a00", 515=>x"9a00", 516=>x"9d00",
---- 517=>x"9c00", 518=>x"9a00", 519=>x"9b00", 520=>x"9b00",
---- 521=>x"9b00", 522=>x"9b00", 523=>x"9e00", 524=>x"9b00",
---- 525=>x"9700", 526=>x"9800", 527=>x"9d00", 528=>x"9800",
---- 529=>x"9900", 530=>x"9900", 531=>x"9b00", 532=>x"9a00",
---- 533=>x"9b00", 534=>x"9800", 535=>x"9a00", 536=>x"9600",
---- 537=>x"9700", 538=>x"9700", 539=>x"9900", 540=>x"9900",
---- 541=>x"9600", 542=>x"9700", 543=>x"9a00", 544=>x"9f00",
---- 545=>x"9a00", 546=>x"9600", 547=>x"9900", 548=>x"9e00",
---- 549=>x"a400", 550=>x"9800", 551=>x"9a00", 552=>x"9f00",
---- 553=>x"a900", 554=>x"9900", 555=>x"9800", 556=>x"9a00",
---- 557=>x"9700", 558=>x"9500", 559=>x"9900", 560=>x"9600",
---- 561=>x"9600", 562=>x"9700", 563=>x"9800", 564=>x"9700",
---- 565=>x"9400", 566=>x"9600", 567=>x"9500", 568=>x"9800",
---- 569=>x"9700", 570=>x"9600", 571=>x"9700", 572=>x"9700",
---- 573=>x"9500", 574=>x"9400", 575=>x"9700", 576=>x"9600",
---- 577=>x"6c00", 578=>x"9500", 579=>x"9700", 580=>x"9800",
---- 581=>x"9400", 582=>x"9300", 583=>x"9300", 584=>x"9600",
---- 585=>x"9200", 586=>x"9300", 587=>x"9300", 588=>x"9500",
---- 589=>x"9400", 590=>x"9200", 591=>x"9200", 592=>x"9500",
---- 593=>x"9300", 594=>x"9300", 595=>x"9300", 596=>x"9400",
---- 597=>x"9300", 598=>x"9400", 599=>x"9400", 600=>x"9500",
---- 601=>x"9200", 602=>x"9200", 603=>x"9400", 604=>x"9200",
---- 605=>x"6f00", 606=>x"9000", 607=>x"8e00", 608=>x"9200",
---- 609=>x"9000", 610=>x"9000", 611=>x"9300", 612=>x"9200",
---- 613=>x"9000", 614=>x"8e00", 615=>x"8f00", 616=>x"9300",
---- 617=>x"9100", 618=>x"8f00", 619=>x"9000", 620=>x"9200",
---- 621=>x"9200", 622=>x"9000", 623=>x"9000", 624=>x"9100",
---- 625=>x"9100", 626=>x"8f00", 627=>x"9100", 628=>x"9400",
---- 629=>x"9300", 630=>x"9100", 631=>x"8e00", 632=>x"9400",
---- 633=>x"9200", 634=>x"9500", 635=>x"9000", 636=>x"9300",
---- 637=>x"9100", 638=>x"9300", 639=>x"9100", 640=>x"6c00",
---- 641=>x"9000", 642=>x"9000", 643=>x"8e00", 644=>x"9000",
---- 645=>x"9100", 646=>x"9000", 647=>x"8e00", 648=>x"9000",
---- 649=>x"9200", 650=>x"9000", 651=>x"8d00", 652=>x"9200",
---- 653=>x"9000", 654=>x"8c00", 655=>x"8e00", 656=>x"8f00",
---- 657=>x"8e00", 658=>x"8f00", 659=>x"9100", 660=>x"9200",
---- 661=>x"8e00", 662=>x"8d00", 663=>x"8d00", 664=>x"9000",
---- 665=>x"9000", 666=>x"8e00", 667=>x"8d00", 668=>x"8e00",
---- 669=>x"8d00", 670=>x"8c00", 671=>x"8e00", 672=>x"9000",
---- 673=>x"8e00", 674=>x"8c00", 675=>x"8d00", 676=>x"9000",
---- 677=>x"8d00", 678=>x"8d00", 679=>x"8d00", 680=>x"8f00",
---- 681=>x"8f00", 682=>x"8a00", 683=>x"8500", 684=>x"9000",
---- 685=>x"8e00", 686=>x"8900", 687=>x"8500", 688=>x"8e00",
---- 689=>x"8c00", 690=>x"8b00", 691=>x"8a00", 692=>x"8d00",
---- 693=>x"8b00", 694=>x"8b00", 695=>x"8800", 696=>x"9000",
---- 697=>x"8d00", 698=>x"8b00", 699=>x"7700", 700=>x"9100",
---- 701=>x"8f00", 702=>x"8a00", 703=>x"8500", 704=>x"8f00",
---- 705=>x"8d00", 706=>x"8900", 707=>x"8600", 708=>x"9100",
---- 709=>x"8b00", 710=>x"8a00", 711=>x"8500", 712=>x"8e00",
---- 713=>x"8d00", 714=>x"8700", 715=>x"8400", 716=>x"8f00",
---- 717=>x"8c00", 718=>x"8700", 719=>x"8300", 720=>x"9200",
---- 721=>x"8c00", 722=>x"8600", 723=>x"8400", 724=>x"8e00",
---- 725=>x"8a00", 726=>x"8300", 727=>x"8400", 728=>x"8b00",
---- 729=>x"8900", 730=>x"8300", 731=>x"7f00", 732=>x"8e00",
---- 733=>x"8700", 734=>x"8300", 735=>x"7e00", 736=>x"8c00",
---- 737=>x"8700", 738=>x"8000", 739=>x"7e00", 740=>x"8900",
---- 741=>x"7a00", 742=>x"7f00", 743=>x"7a00", 744=>x"8a00",
---- 745=>x"8700", 746=>x"7f00", 747=>x"7800", 748=>x"8900",
---- 749=>x"8800", 750=>x"8000", 751=>x"7b00", 752=>x"8600",
---- 753=>x"8500", 754=>x"8100", 755=>x"7d00", 756=>x"8800",
---- 757=>x"8400", 758=>x"8000", 759=>x"7900", 760=>x"8600",
---- 761=>x"8200", 762=>x"7e00", 763=>x"7700", 764=>x"8700",
---- 765=>x"8100", 766=>x"7e00", 767=>x"7800", 768=>x"8800",
---- 769=>x"8000", 770=>x"7a00", 771=>x"7400", 772=>x"8200",
---- 773=>x"7c00", 774=>x"8700", 775=>x"7200", 776=>x"8000",
---- 777=>x"7d00", 778=>x"7500", 779=>x"7000", 780=>x"7d00",
---- 781=>x"7900", 782=>x"7500", 783=>x"7100", 784=>x"7e00",
---- 785=>x"7a00", 786=>x"7500", 787=>x"8c00", 788=>x"7d00",
---- 789=>x"7a00", 790=>x"7400", 791=>x"7300", 792=>x"7500",
---- 793=>x"8e00", 794=>x"6d00", 795=>x"7100", 796=>x"6c00",
---- 797=>x"6300", 798=>x"6000", 799=>x"6600", 800=>x"6b00",
---- 801=>x"5d00", 802=>x"4e00", 803=>x"5600", 804=>x"7200",
---- 805=>x"6100", 806=>x"4c00", 807=>x"4e00", 808=>x"7400",
---- 809=>x"6500", 810=>x"4b00", 811=>x"5000", 812=>x"7600",
---- 813=>x"6300", 814=>x"4d00", 815=>x"5f00", 816=>x"8700",
---- 817=>x"6500", 818=>x"5500", 819=>x"7900", 820=>x"7800",
---- 821=>x"6c00", 822=>x"6200", 823=>x"8d00", 824=>x"8000",
---- 825=>x"7100", 826=>x"6f00", 827=>x"9d00", 828=>x"8000",
---- 829=>x"7600", 830=>x"7e00", 831=>x"af00", 832=>x"8300",
---- 833=>x"7900", 834=>x"8b00", 835=>x"bd00", 836=>x"8900",
---- 837=>x"7f00", 838=>x"9600", 839=>x"c200", 840=>x"8b00",
---- 841=>x"8700", 842=>x"a300", 843=>x"c600", 844=>x"9e00",
---- 845=>x"a400", 846=>x"b500", 847=>x"c700", 848=>x"b300",
---- 849=>x"bc00", 850=>x"c700", 851=>x"cd00", 852=>x"c000",
---- 853=>x"c400", 854=>x"ca00", 855=>x"d100", 856=>x"c700",
---- 857=>x"ca00", 858=>x"cf00", 859=>x"d600", 860=>x"c900",
---- 861=>x"cb00", 862=>x"cf00", 863=>x"d600", 864=>x"ce00",
---- 865=>x"cb00", 866=>x"cd00", 867=>x"d500", 868=>x"d100",
---- 869=>x"cf00", 870=>x"d100", 871=>x"d400", 872=>x"d200",
---- 873=>x"d200", 874=>x"d400", 875=>x"d700", 876=>x"d000",
---- 877=>x"d000", 878=>x"d500", 879=>x"d800", 880=>x"ce00",
---- 881=>x"d100", 882=>x"d500", 883=>x"da00", 884=>x"cc00",
---- 885=>x"d100", 886=>x"d500", 887=>x"2400", 888=>x"cc00",
---- 889=>x"d100", 890=>x"2900", 891=>x"da00", 892=>x"cc00",
---- 893=>x"d000", 894=>x"d800", 895=>x"dc00", 896=>x"ca00",
---- 897=>x"d100", 898=>x"d800", 899=>x"db00", 900=>x"ca00",
---- 901=>x"d200", 902=>x"da00", 903=>x"db00", 904=>x"c900",
---- 905=>x"d600", 906=>x"db00", 907=>x"d900", 908=>x"c900",
---- 909=>x"d400", 910=>x"db00", 911=>x"d700", 912=>x"cc00",
---- 913=>x"d800", 914=>x"dc00", 915=>x"d800", 916=>x"cf00",
---- 917=>x"dc00", 918=>x"dc00", 919=>x"d700", 920=>x"d300",
---- 921=>x"dd00", 922=>x"dc00", 923=>x"d500", 924=>x"d500",
---- 925=>x"dc00", 926=>x"da00", 927=>x"d100", 928=>x"d800",
---- 929=>x"de00", 930=>x"2700", 931=>x"ce00", 932=>x"da00",
---- 933=>x"dc00", 934=>x"d500", 935=>x"c500", 936=>x"dc00",
---- 937=>x"da00", 938=>x"3000", 939=>x"b800", 940=>x"2500",
---- 941=>x"d500", 942=>x"c900", 943=>x"ad00", 944=>x"d900",
---- 945=>x"d200", 946=>x"c100", 947=>x"a100", 948=>x"d600",
---- 949=>x"cd00", 950=>x"b500", 951=>x"8c00", 952=>x"d200",
---- 953=>x"c300", 954=>x"a000", 955=>x"6400", 956=>x"c500",
---- 957=>x"a800", 958=>x"7300", 959=>x"4200", 960=>x"a700",
---- 961=>x"7700", 962=>x"4400", 963=>x"3700", 964=>x"7900",
---- 965=>x"5000", 966=>x"3800", 967=>x"3400", 968=>x"5100",
---- 969=>x"4300", 970=>x"3500", 971=>x"3400", 972=>x"4300",
---- 973=>x"3b00", 974=>x"3600", 975=>x"3c00", 976=>x"4200",
---- 977=>x"3e00", 978=>x"4100", 979=>x"4800", 980=>x"4800",
---- 981=>x"4700", 982=>x"4d00", 983=>x"4b00", 984=>x"4f00",
---- 985=>x"5400", 986=>x"5100", 987=>x"4f00", 988=>x"5b00",
---- 989=>x"5600", 990=>x"aa00", 991=>x"4e00", 992=>x"5f00",
---- 993=>x"5600", 994=>x"5500", 995=>x"4c00", 996=>x"6100",
---- 997=>x"5a00", 998=>x"5300", 999=>x"4f00", 1000=>x"6100",
---- 1001=>x"5c00", 1002=>x"5300", 1003=>x"5400", 1004=>x"6200",
---- 1005=>x"5c00", 1006=>x"5700", 1007=>x"5e00", 1008=>x"6000",
---- 1009=>x"5e00", 1010=>x"5f00", 1011=>x"6600", 1012=>x"5d00",
---- 1013=>x"5d00", 1014=>x"a100", 1015=>x"6300", 1016=>x"6000",
---- 1017=>x"a200", 1018=>x"5900", 1019=>x"5900", 1020=>x"5c00",
---- 1021=>x"5700", 1022=>x"4f00", 1023=>x"4c00"),
----
---- 56 => (0=>x"7900", 1=>x"7e00", 2=>x"7a00", 3=>x"7800", 4=>x"7900",
---- 5=>x"7f00", 6=>x"7a00", 7=>x"7800", 8=>x"7b00",
---- 9=>x"7c00", 10=>x"7a00", 11=>x"7700", 12=>x"7a00",
---- 13=>x"7c00", 14=>x"7a00", 15=>x"7800", 16=>x"7700",
---- 17=>x"7900", 18=>x"7b00", 19=>x"7a00", 20=>x"7900",
---- 21=>x"7a00", 22=>x"7800", 23=>x"7900", 24=>x"7900",
---- 25=>x"7a00", 26=>x"7800", 27=>x"7900", 28=>x"7700",
---- 29=>x"7700", 30=>x"7c00", 31=>x"7a00", 32=>x"7800",
---- 33=>x"7700", 34=>x"7a00", 35=>x"7800", 36=>x"7700",
---- 37=>x"7a00", 38=>x"7c00", 39=>x"8500", 40=>x"7600",
---- 41=>x"7a00", 42=>x"7900", 43=>x"7b00", 44=>x"7500",
---- 45=>x"7400", 46=>x"7200", 47=>x"7a00", 48=>x"7700",
---- 49=>x"7900", 50=>x"7800", 51=>x"7800", 52=>x"7a00",
---- 53=>x"7b00", 54=>x"7c00", 55=>x"7b00", 56=>x"7700",
---- 57=>x"7900", 58=>x"7900", 59=>x"7a00", 60=>x"7300",
---- 61=>x"7400", 62=>x"7500", 63=>x"7a00", 64=>x"7300",
---- 65=>x"7700", 66=>x"7500", 67=>x"7800", 68=>x"7000",
---- 69=>x"7200", 70=>x"7400", 71=>x"7500", 72=>x"6c00",
---- 73=>x"7200", 74=>x"7300", 75=>x"7300", 76=>x"6b00",
---- 77=>x"6e00", 78=>x"7000", 79=>x"7200", 80=>x"6a00",
---- 81=>x"6e00", 82=>x"6b00", 83=>x"7200", 84=>x"6300",
---- 85=>x"6b00", 86=>x"6b00", 87=>x"6e00", 88=>x"6200",
---- 89=>x"6800", 90=>x"6a00", 91=>x"6c00", 92=>x"6e00",
---- 93=>x"6a00", 94=>x"6f00", 95=>x"6d00", 96=>x"9200",
---- 97=>x"6c00", 98=>x"6c00", 99=>x"6e00", 100=>x"b600",
---- 101=>x"7f00", 102=>x"6a00", 103=>x"7300", 104=>x"cd00",
---- 105=>x"a400", 106=>x"7600", 107=>x"7400", 108=>x"da00",
---- 109=>x"c600", 110=>x"9000", 111=>x"7800", 112=>x"e100",
---- 113=>x"d800", 114=>x"b500", 115=>x"7a00", 116=>x"e400",
---- 117=>x"df00", 118=>x"d100", 119=>x"8100", 120=>x"e400",
---- 121=>x"e400", 122=>x"db00", 123=>x"7700", 124=>x"e600",
---- 125=>x"e400", 126=>x"c100", 127=>x"4600", 128=>x"e100",
---- 129=>x"d300", 130=>x"7600", 131=>x"2000", 132=>x"d500",
---- 133=>x"9000", 134=>x"3100", 135=>x"2300", 136=>x"9400",
---- 137=>x"3700", 138=>x"2600", 139=>x"2900", 140=>x"3700",
---- 141=>x"2800", 142=>x"2f00", 143=>x"2c00", 144=>x"2a00",
---- 145=>x"2e00", 146=>x"3000", 147=>x"2a00", 148=>x"2e00",
---- 149=>x"2c00", 150=>x"2a00", 151=>x"2c00", 152=>x"2a00",
---- 153=>x"2b00", 154=>x"2e00", 155=>x"2900", 156=>x"3000",
---- 157=>x"2700", 158=>x"2d00", 159=>x"2d00", 160=>x"2b00",
---- 161=>x"2a00", 162=>x"3200", 163=>x"3000", 164=>x"2b00",
---- 165=>x"2c00", 166=>x"2e00", 167=>x"3000", 168=>x"2f00",
---- 169=>x"2d00", 170=>x"3300", 171=>x"3400", 172=>x"2b00",
---- 173=>x"3000", 174=>x"3700", 175=>x"3800", 176=>x"3300",
---- 177=>x"3b00", 178=>x"3900", 179=>x"3500", 180=>x"3a00",
---- 181=>x"3800", 182=>x"3400", 183=>x"3700", 184=>x"3400",
---- 185=>x"3400", 186=>x"3200", 187=>x"3400", 188=>x"ca00",
---- 189=>x"3400", 190=>x"3800", 191=>x"3700", 192=>x"3900",
---- 193=>x"3200", 194=>x"3600", 195=>x"3100", 196=>x"3600",
---- 197=>x"3400", 198=>x"3400", 199=>x"2f00", 200=>x"3800",
---- 201=>x"3500", 202=>x"3400", 203=>x"3200", 204=>x"3500",
---- 205=>x"3800", 206=>x"ce00", 207=>x"2e00", 208=>x"3b00",
---- 209=>x"3700", 210=>x"2f00", 211=>x"2c00", 212=>x"3700",
---- 213=>x"3300", 214=>x"2f00", 215=>x"2d00", 216=>x"3600",
---- 217=>x"2e00", 218=>x"2e00", 219=>x"3500", 220=>x"3300",
---- 221=>x"3000", 222=>x"3300", 223=>x"3600", 224=>x"3400",
---- 225=>x"3500", 226=>x"3200", 227=>x"3600", 228=>x"3200",
---- 229=>x"3800", 230=>x"3600", 231=>x"3200", 232=>x"3600",
---- 233=>x"3500", 234=>x"3800", 235=>x"3400", 236=>x"3400",
---- 237=>x"3500", 238=>x"3500", 239=>x"3200", 240=>x"3300",
---- 241=>x"3400", 242=>x"2e00", 243=>x"2e00", 244=>x"3700",
---- 245=>x"d000", 246=>x"2f00", 247=>x"3000", 248=>x"2a00",
---- 249=>x"2800", 250=>x"3300", 251=>x"3100", 252=>x"2800",
---- 253=>x"2e00", 254=>x"3300", 255=>x"3000", 256=>x"d200",
---- 257=>x"2e00", 258=>x"3100", 259=>x"3300", 260=>x"3200",
---- 261=>x"3300", 262=>x"3400", 263=>x"3300", 264=>x"3500",
---- 265=>x"3700", 266=>x"3600", 267=>x"3700", 268=>x"3300",
---- 269=>x"3400", 270=>x"3600", 271=>x"3400", 272=>x"3300",
---- 273=>x"3500", 274=>x"3500", 275=>x"3000", 276=>x"3400",
---- 277=>x"3200", 278=>x"3000", 279=>x"2d00", 280=>x"3400",
---- 281=>x"3500", 282=>x"3600", 283=>x"ca00", 284=>x"3300",
---- 285=>x"3700", 286=>x"3c00", 287=>x"4100", 288=>x"3200",
---- 289=>x"3600", 290=>x"3f00", 291=>x"4400", 292=>x"3b00",
---- 293=>x"4000", 294=>x"4600", 295=>x"5700", 296=>x"3500",
---- 297=>x"3900", 298=>x"4c00", 299=>x"6900", 300=>x"2c00",
---- 301=>x"3b00", 302=>x"5c00", 303=>x"7f00", 304=>x"2700",
---- 305=>x"4000", 306=>x"6d00", 307=>x"8e00", 308=>x"3000",
---- 309=>x"5400", 310=>x"8000", 311=>x"9700", 312=>x"4700",
---- 313=>x"6e00", 314=>x"8e00", 315=>x"9900", 316=>x"6300",
---- 317=>x"7b00", 318=>x"9500", 319=>x"9700", 320=>x"7b00",
---- 321=>x"9200", 322=>x"9700", 323=>x"9500", 324=>x"8c00",
---- 325=>x"9c00", 326=>x"9800", 327=>x"9200", 328=>x"9600",
---- 329=>x"9b00", 330=>x"9400", 331=>x"9100", 332=>x"9a00",
---- 333=>x"9800", 334=>x"9100", 335=>x"8e00", 336=>x"9900",
---- 337=>x"9400", 338=>x"9400", 339=>x"8e00", 340=>x"9500",
---- 341=>x"9300", 342=>x"9100", 343=>x"9400", 344=>x"9200",
---- 345=>x"9100", 346=>x"9300", 347=>x"9900", 348=>x"9300",
---- 349=>x"9100", 350=>x"9600", 351=>x"9e00", 352=>x"9000",
---- 353=>x"9300", 354=>x"9900", 355=>x"9f00", 356=>x"8e00",
---- 357=>x"9700", 358=>x"a000", 359=>x"a100", 360=>x"6f00",
---- 361=>x"9c00", 362=>x"a000", 363=>x"a100", 364=>x"9800",
---- 365=>x"a000", 366=>x"a300", 367=>x"a100", 368=>x"9b00",
---- 369=>x"a300", 370=>x"a300", 371=>x"a100", 372=>x"9f00",
---- 373=>x"a400", 374=>x"a400", 375=>x"a200", 376=>x"a500",
---- 377=>x"a600", 378=>x"a400", 379=>x"a300", 380=>x"a400",
---- 381=>x"a500", 382=>x"a400", 383=>x"a200", 384=>x"a500",
---- 385=>x"a400", 386=>x"a400", 387=>x"a300", 388=>x"a300",
---- 389=>x"a400", 390=>x"a600", 391=>x"a500", 392=>x"a400",
---- 393=>x"a400", 394=>x"a400", 395=>x"a500", 396=>x"a700",
---- 397=>x"a600", 398=>x"a400", 399=>x"a600", 400=>x"a400",
---- 401=>x"a600", 402=>x"a500", 403=>x"a500", 404=>x"a400",
---- 405=>x"a400", 406=>x"5900", 407=>x"a600", 408=>x"a600",
---- 409=>x"a500", 410=>x"a100", 411=>x"a500", 412=>x"a400",
---- 413=>x"a400", 414=>x"a200", 415=>x"a300", 416=>x"a300",
---- 417=>x"a200", 418=>x"a200", 419=>x"a300", 420=>x"a600",
---- 421=>x"a200", 422=>x"a400", 423=>x"a300", 424=>x"a600",
---- 425=>x"a400", 426=>x"a600", 427=>x"a300", 428=>x"a500",
---- 429=>x"a700", 430=>x"a500", 431=>x"a200", 432=>x"a200",
---- 433=>x"a500", 434=>x"a300", 435=>x"a300", 436=>x"a400",
---- 437=>x"a500", 438=>x"a600", 439=>x"a500", 440=>x"a600",
---- 441=>x"a700", 442=>x"a600", 443=>x"a500", 444=>x"9f00",
---- 445=>x"a300", 446=>x"a500", 447=>x"a200", 448=>x"9a00",
---- 449=>x"9a00", 450=>x"9e00", 451=>x"9e00", 452=>x"9500",
---- 453=>x"9700", 454=>x"9600", 455=>x"9800", 456=>x"9700",
---- 457=>x"9600", 458=>x"9400", 459=>x"9600", 460=>x"9700",
---- 461=>x"9500", 462=>x"9400", 463=>x"9300", 464=>x"9600",
---- 465=>x"9800", 466=>x"9700", 467=>x"9600", 468=>x"9e00",
---- 469=>x"9c00", 470=>x"9a00", 471=>x"9a00", 472=>x"a200",
---- 473=>x"9f00", 474=>x"a100", 475=>x"9e00", 476=>x"a300",
---- 477=>x"a300", 478=>x"a400", 479=>x"a400", 480=>x"a500",
---- 481=>x"a600", 482=>x"5a00", 483=>x"a500", 484=>x"a400",
---- 485=>x"a300", 486=>x"a800", 487=>x"a600", 488=>x"a300",
---- 489=>x"a300", 490=>x"a200", 491=>x"a400", 492=>x"9e00",
---- 493=>x"9f00", 494=>x"a200", 495=>x"a100", 496=>x"9d00",
---- 497=>x"9e00", 498=>x"9f00", 499=>x"9f00", 500=>x"9b00",
---- 501=>x"9e00", 502=>x"9c00", 503=>x"9e00", 504=>x"9c00",
---- 505=>x"9c00", 506=>x"9c00", 507=>x"9e00", 508=>x"9a00",
---- 509=>x"9a00", 510=>x"9d00", 511=>x"9e00", 512=>x"9c00",
---- 513=>x"9c00", 514=>x"9c00", 515=>x"9d00", 516=>x"9b00",
---- 517=>x"9c00", 518=>x"9c00", 519=>x"9c00", 520=>x"9a00",
---- 521=>x"9a00", 522=>x"9c00", 523=>x"9a00", 524=>x"9b00",
---- 525=>x"9900", 526=>x"9a00", 527=>x"9d00", 528=>x"9900",
---- 529=>x"9a00", 530=>x"9b00", 531=>x"9800", 532=>x"9800",
---- 533=>x"9900", 534=>x"9800", 535=>x"9600", 536=>x"9900",
---- 537=>x"9b00", 538=>x"9800", 539=>x"9800", 540=>x"9700",
---- 541=>x"9b00", 542=>x"9b00", 543=>x"9600", 544=>x"9900",
---- 545=>x"9800", 546=>x"9a00", 547=>x"9a00", 548=>x"9700",
---- 549=>x"9800", 550=>x"9b00", 551=>x"9900", 552=>x"9700",
---- 553=>x"9a00", 554=>x"9a00", 555=>x"9a00", 556=>x"9700",
---- 557=>x"9500", 558=>x"9600", 559=>x"9b00", 560=>x"9700",
---- 561=>x"9600", 562=>x"9600", 563=>x"9600", 564=>x"9600",
---- 565=>x"9800", 566=>x"9600", 567=>x"9700", 568=>x"9500",
---- 569=>x"9500", 570=>x"9600", 571=>x"9600", 572=>x"9500",
---- 573=>x"9400", 574=>x"9300", 575=>x"9300", 576=>x"9600",
---- 577=>x"9400", 578=>x"9300", 579=>x"9100", 580=>x"9300",
---- 581=>x"9100", 582=>x"9300", 583=>x"9200", 584=>x"9400",
---- 585=>x"9100", 586=>x"6c00", 587=>x"9100", 588=>x"9000",
---- 589=>x"9300", 590=>x"9000", 591=>x"8e00", 592=>x"9000",
---- 593=>x"9100", 594=>x"9300", 595=>x"8f00", 596=>x"9100",
---- 597=>x"9000", 598=>x"9300", 599=>x"9100", 600=>x"9000",
---- 601=>x"8f00", 602=>x"8f00", 603=>x"8f00", 604=>x"7000",
---- 605=>x"9100", 606=>x"6f00", 607=>x"8e00", 608=>x"9100",
---- 609=>x"8d00", 610=>x"9000", 611=>x"8d00", 612=>x"8f00",
---- 613=>x"8c00", 614=>x"8d00", 615=>x"8a00", 616=>x"8d00",
---- 617=>x"8b00", 618=>x"8900", 619=>x"8a00", 620=>x"8d00",
---- 621=>x"8900", 622=>x"8d00", 623=>x"8c00", 624=>x"8f00",
---- 625=>x"7500", 626=>x"8c00", 627=>x"8a00", 628=>x"8f00",
---- 629=>x"8d00", 630=>x"8900", 631=>x"8600", 632=>x"8d00",
---- 633=>x"8a00", 634=>x"8a00", 635=>x"8400", 636=>x"8f00",
---- 637=>x"8a00", 638=>x"8800", 639=>x"8200", 640=>x"8c00",
---- 641=>x"8b00", 642=>x"8700", 643=>x"8300", 644=>x"8d00",
---- 645=>x"8b00", 646=>x"8600", 647=>x"8100", 648=>x"7100",
---- 649=>x"8800", 650=>x"8600", 651=>x"8400", 652=>x"8d00",
---- 653=>x"7700", 654=>x"8700", 655=>x"8400", 656=>x"8c00",
---- 657=>x"8700", 658=>x"8400", 659=>x"8800", 660=>x"8900",
---- 661=>x"8600", 662=>x"8300", 663=>x"8900", 664=>x"8700",
---- 665=>x"8600", 666=>x"7a00", 667=>x"9100", 668=>x"8800",
---- 669=>x"8300", 670=>x"8300", 671=>x"9600", 672=>x"7500",
---- 673=>x"8300", 674=>x"8600", 675=>x"9a00", 676=>x"8900",
---- 677=>x"8400", 678=>x"8600", 679=>x"9e00", 680=>x"8300",
---- 681=>x"8200", 682=>x"8600", 683=>x"a200", 684=>x"8300",
---- 685=>x"8000", 686=>x"8800", 687=>x"a300", 688=>x"8500",
---- 689=>x"7f00", 690=>x"8900", 691=>x"a600", 692=>x"8400",
---- 693=>x"7e00", 694=>x"8b00", 695=>x"a600", 696=>x"8200",
---- 697=>x"7d00", 698=>x"8e00", 699=>x"5400", 700=>x"7f00",
---- 701=>x"7e00", 702=>x"9100", 703=>x"ad00", 704=>x"8100",
---- 705=>x"8000", 706=>x"9500", 707=>x"af00", 708=>x"7f00",
---- 709=>x"7f00", 710=>x"9800", 711=>x"b300", 712=>x"7e00",
---- 713=>x"7f00", 714=>x"9900", 715=>x"b500", 716=>x"7d00",
---- 717=>x"7e00", 718=>x"9d00", 719=>x"b800", 720=>x"7c00",
---- 721=>x"7e00", 722=>x"6300", 723=>x"ba00", 724=>x"7a00",
---- 725=>x"7d00", 726=>x"9e00", 727=>x"bf00", 728=>x"7700",
---- 729=>x"7b00", 730=>x"9e00", 731=>x"c000", 732=>x"7500",
---- 733=>x"7700", 734=>x"9b00", 735=>x"c300", 736=>x"7900",
---- 737=>x"7800", 738=>x"6300", 739=>x"c300", 740=>x"7700",
---- 741=>x"7400", 742=>x"9d00", 743=>x"c800", 744=>x"7600",
---- 745=>x"7600", 746=>x"a300", 747=>x"c800", 748=>x"7300",
---- 749=>x"7900", 750=>x"aa00", 751=>x"cd00", 752=>x"7300",
---- 753=>x"7e00", 754=>x"b300", 755=>x"2e00", 756=>x"7100",
---- 757=>x"8200", 758=>x"b800", 759=>x"d400", 760=>x"7500",
---- 761=>x"8c00", 762=>x"be00", 763=>x"d500", 764=>x"7400",
---- 765=>x"9600", 766=>x"c500", 767=>x"d600", 768=>x"7600",
---- 769=>x"a400", 770=>x"c900", 771=>x"d600", 772=>x"7e00",
---- 773=>x"b100", 774=>x"3000", 775=>x"d900", 776=>x"8700",
---- 777=>x"bc00", 778=>x"d100", 779=>x"d900", 780=>x"9600",
---- 781=>x"c400", 782=>x"d500", 783=>x"da00", 784=>x"9c00",
---- 785=>x"c800", 786=>x"d400", 787=>x"d700", 788=>x"9f00",
---- 789=>x"c900", 790=>x"d200", 791=>x"d600", 792=>x"9f00",
---- 793=>x"ca00", 794=>x"d000", 795=>x"d400", 796=>x"9c00",
---- 797=>x"3d00", 798=>x"ce00", 799=>x"d200", 800=>x"8e00",
---- 801=>x"c000", 802=>x"cf00", 803=>x"d100", 804=>x"8a00",
---- 805=>x"c200", 806=>x"cf00", 807=>x"cf00", 808=>x"9200",
---- 809=>x"c400", 810=>x"d100", 811=>x"d100", 812=>x"a200",
---- 813=>x"c800", 814=>x"d000", 815=>x"d200", 816=>x"b300",
---- 817=>x"cd00", 818=>x"d300", 819=>x"d400", 820=>x"be00",
---- 821=>x"cc00", 822=>x"d400", 823=>x"d400", 824=>x"c500",
---- 825=>x"d100", 826=>x"d400", 827=>x"d400", 828=>x"cb00",
---- 829=>x"d300", 830=>x"d500", 831=>x"d500", 832=>x"cd00",
---- 833=>x"d600", 834=>x"d600", 835=>x"d400", 836=>x"2d00",
---- 837=>x"d900", 838=>x"d600", 839=>x"d400", 840=>x"d300",
---- 841=>x"d900", 842=>x"d600", 843=>x"d400", 844=>x"d400",
---- 845=>x"d700", 846=>x"d600", 847=>x"d600", 848=>x"d400",
---- 849=>x"d700", 850=>x"d700", 851=>x"d700", 852=>x"d600",
---- 853=>x"d900", 854=>x"d700", 855=>x"d600", 856=>x"2700",
---- 857=>x"d900", 858=>x"d700", 859=>x"d700", 860=>x"da00",
---- 861=>x"d700", 862=>x"d800", 863=>x"d600", 864=>x"d800",
---- 865=>x"d800", 866=>x"d800", 867=>x"d600", 868=>x"da00",
---- 869=>x"d900", 870=>x"d900", 871=>x"d600", 872=>x"da00",
---- 873=>x"d900", 874=>x"d800", 875=>x"d500", 876=>x"d900",
---- 877=>x"d800", 878=>x"d500", 879=>x"d100", 880=>x"2600",
---- 881=>x"d800", 882=>x"d700", 883=>x"ce00", 884=>x"da00",
---- 885=>x"d700", 886=>x"d200", 887=>x"c800", 888=>x"d900",
---- 889=>x"d600", 890=>x"cf00", 891=>x"bd00", 892=>x"2700",
---- 893=>x"d400", 894=>x"c900", 895=>x"b300", 896=>x"d700",
---- 897=>x"d000", 898=>x"c500", 899=>x"a800", 900=>x"d600",
---- 901=>x"cd00", 902=>x"bf00", 903=>x"9f00", 904=>x"d200",
---- 905=>x"cc00", 906=>x"ba00", 907=>x"9600", 908=>x"d100",
---- 909=>x"c900", 910=>x"b400", 911=>x"8f00", 912=>x"d100",
---- 913=>x"c600", 914=>x"ab00", 915=>x"8700", 916=>x"d000",
---- 917=>x"be00", 918=>x"a000", 919=>x"8000", 920=>x"cc00",
---- 921=>x"b400", 922=>x"9300", 923=>x"7800", 924=>x"c500",
---- 925=>x"aa00", 926=>x"8700", 927=>x"7600", 928=>x"ba00",
---- 929=>x"9b00", 930=>x"8000", 931=>x"6e00", 932=>x"a700",
---- 933=>x"8a00", 934=>x"7500", 935=>x"6200", 936=>x"9800",
---- 937=>x"7d00", 938=>x"6300", 939=>x"5300", 940=>x"8a00",
---- 941=>x"6b00", 942=>x"5600", 943=>x"4700", 944=>x"7700",
---- 945=>x"5700", 946=>x"4b00", 947=>x"3e00", 948=>x"6100",
---- 949=>x"b800", 950=>x"3d00", 951=>x"3b00", 952=>x"4500",
---- 953=>x"3d00", 954=>x"ca00", 955=>x"3f00", 956=>x"3700",
---- 957=>x"3800", 958=>x"3d00", 959=>x"4200", 960=>x"3400",
---- 961=>x"3400", 962=>x"3e00", 963=>x"4600", 964=>x"3600",
---- 965=>x"3700", 966=>x"4300", 967=>x"4900", 968=>x"3d00",
---- 969=>x"4400", 970=>x"4900", 971=>x"4700", 972=>x"4400",
---- 973=>x"4c00", 974=>x"4800", 975=>x"4200", 976=>x"4c00",
---- 977=>x"4b00", 978=>x"b800", 979=>x"4700", 980=>x"4e00",
---- 981=>x"4900", 982=>x"4700", 983=>x"5000", 984=>x"4c00",
---- 985=>x"4600", 986=>x"4f00", 987=>x"5800", 988=>x"4800",
---- 989=>x"4800", 990=>x"5400", 991=>x"5f00", 992=>x"5000",
---- 993=>x"5100", 994=>x"5900", 995=>x"6700", 996=>x"5400",
---- 997=>x"5700", 998=>x"6000", 999=>x"6600", 1000=>x"5b00",
---- 1001=>x"6000", 1002=>x"6300", 1003=>x"5e00", 1004=>x"6100",
---- 1005=>x"6200", 1006=>x"6400", 1007=>x"5800", 1008=>x"6400",
---- 1009=>x"5d00", 1010=>x"5a00", 1011=>x"5700", 1012=>x"5b00",
---- 1013=>x"5600", 1014=>x"5000", 1015=>x"5100", 1016=>x"4f00",
---- 1017=>x"4e00", 1018=>x"4d00", 1019=>x"5500", 1020=>x"4a00",
---- 1021=>x"4a00", 1022=>x"5400", 1023=>x"5c00"),
----
---- 57 => (0=>x"7800", 1=>x"7a00", 2=>x"7900", 3=>x"7a00", 4=>x"7800",
---- 5=>x"7a00", 6=>x"7900", 7=>x"7a00", 8=>x"7800",
---- 9=>x"7a00", 10=>x"7800", 11=>x"7a00", 12=>x"7a00",
---- 13=>x"7900", 14=>x"7900", 15=>x"7c00", 16=>x"7800",
---- 17=>x"7800", 18=>x"7b00", 19=>x"7c00", 20=>x"7700",
---- 21=>x"7800", 22=>x"7800", 23=>x"7800", 24=>x"7a00",
---- 25=>x"7500", 26=>x"7800", 27=>x"7900", 28=>x"7800",
---- 29=>x"7800", 30=>x"7900", 31=>x"7a00", 32=>x"7700",
---- 33=>x"7c00", 34=>x"7900", 35=>x"7b00", 36=>x"7c00",
---- 37=>x"7f00", 38=>x"7a00", 39=>x"7b00", 40=>x"7a00",
---- 41=>x"7900", 42=>x"7900", 43=>x"7b00", 44=>x"7a00",
---- 45=>x"7900", 46=>x"7900", 47=>x"7800", 48=>x"7a00",
---- 49=>x"7a00", 50=>x"7a00", 51=>x"7800", 52=>x"8400",
---- 53=>x"7c00", 54=>x"7a00", 55=>x"7900", 56=>x"7b00",
---- 57=>x"7a00", 58=>x"7900", 59=>x"7a00", 60=>x"7b00",
---- 61=>x"7700", 62=>x"7a00", 63=>x"7800", 64=>x"7900",
---- 65=>x"7a00", 66=>x"7900", 67=>x"7900", 68=>x"7800",
---- 69=>x"7b00", 70=>x"7b00", 71=>x"7900", 72=>x"7700",
---- 73=>x"7b00", 74=>x"7b00", 75=>x"7d00", 76=>x"7400",
---- 77=>x"7900", 78=>x"7700", 79=>x"7d00", 80=>x"7300",
---- 81=>x"7300", 82=>x"7600", 83=>x"7b00", 84=>x"6f00",
---- 85=>x"7000", 86=>x"7400", 87=>x"7900", 88=>x"7200",
---- 89=>x"7100", 90=>x"7700", 91=>x"7c00", 92=>x"7500",
---- 93=>x"7300", 94=>x"7b00", 95=>x"7d00", 96=>x"7300",
---- 97=>x"7900", 98=>x"7a00", 99=>x"6d00", 100=>x"7800",
---- 101=>x"7b00", 102=>x"6a00", 103=>x"4800", 104=>x"7900",
---- 105=>x"7200", 106=>x"4b00", 107=>x"d000", 108=>x"7200",
---- 109=>x"5200", 110=>x"3200", 111=>x"2900", 112=>x"5300",
---- 113=>x"3000", 114=>x"2b00", 115=>x"2a00", 116=>x"3100",
---- 117=>x"2a00", 118=>x"2900", 119=>x"2900", 120=>x"2000",
---- 121=>x"2800", 122=>x"2800", 123=>x"2900", 124=>x"2100",
---- 125=>x"2900", 126=>x"2a00", 127=>x"2c00", 128=>x"2a00",
---- 129=>x"2700", 130=>x"2800", 131=>x"2b00", 132=>x"2800",
---- 133=>x"2b00", 134=>x"2a00", 135=>x"2900", 136=>x"2c00",
---- 137=>x"2c00", 138=>x"2d00", 139=>x"2c00", 140=>x"2c00",
---- 141=>x"2b00", 142=>x"2c00", 143=>x"2e00", 144=>x"2b00",
---- 145=>x"2e00", 146=>x"3100", 147=>x"3100", 148=>x"d600",
---- 149=>x"2c00", 150=>x"3100", 151=>x"3900", 152=>x"2900",
---- 153=>x"3100", 154=>x"3400", 155=>x"3500", 156=>x"2c00",
---- 157=>x"3300", 158=>x"3300", 159=>x"3400", 160=>x"2f00",
---- 161=>x"3700", 162=>x"3200", 163=>x"3400", 164=>x"3300",
---- 165=>x"3600", 166=>x"3500", 167=>x"3300", 168=>x"3700",
---- 169=>x"3400", 170=>x"3600", 171=>x"3400", 172=>x"3700",
---- 173=>x"3700", 174=>x"3500", 175=>x"3500", 176=>x"3500",
---- 177=>x"3600", 178=>x"3400", 179=>x"3200", 180=>x"3800",
---- 181=>x"3500", 182=>x"3100", 183=>x"2e00", 184=>x"3600",
---- 185=>x"3400", 186=>x"2e00", 187=>x"2d00", 188=>x"3100",
---- 189=>x"2c00", 190=>x"2800", 191=>x"2a00", 192=>x"2e00",
---- 193=>x"2900", 194=>x"2800", 195=>x"3200", 196=>x"2b00",
---- 197=>x"2d00", 198=>x"2e00", 199=>x"3a00", 200=>x"2700",
---- 201=>x"2b00", 202=>x"3600", 203=>x"3a00", 204=>x"d200",
---- 205=>x"3100", 206=>x"3900", 207=>x"3c00", 208=>x"3200",
---- 209=>x"3800", 210=>x"3500", 211=>x"2d00", 212=>x"3400",
---- 213=>x"3900", 214=>x"3200", 215=>x"2d00", 216=>x"c800",
---- 217=>x"3700", 218=>x"3100", 219=>x"2f00", 220=>x"3700",
---- 221=>x"3300", 222=>x"2f00", 223=>x"3100", 224=>x"3300",
---- 225=>x"2d00", 226=>x"3100", 227=>x"3800", 228=>x"2f00",
---- 229=>x"2f00", 230=>x"3200", 231=>x"3700", 232=>x"2f00",
---- 233=>x"3200", 234=>x"3900", 235=>x"4000", 236=>x"3100",
---- 237=>x"3400", 238=>x"3800", 239=>x"3800", 240=>x"3600",
---- 241=>x"3700", 242=>x"3500", 243=>x"3600", 244=>x"3200",
---- 245=>x"3500", 246=>x"3600", 247=>x"3400", 248=>x"3700",
---- 249=>x"3800", 250=>x"3700", 251=>x"3600", 252=>x"3700",
---- 253=>x"3800", 254=>x"3500", 255=>x"3000", 256=>x"3500",
---- 257=>x"3200", 258=>x"2e00", 259=>x"2c00", 260=>x"3200",
---- 261=>x"2700", 262=>x"2300", 263=>x"3000", 264=>x"2a00",
---- 265=>x"2100", 266=>x"2200", 267=>x"3b00", 268=>x"2600",
---- 269=>x"1f00", 270=>x"2a00", 271=>x"5b00", 272=>x"2300",
---- 273=>x"2400", 274=>x"4100", 275=>x"7400", 276=>x"2c00",
---- 277=>x"3b00", 278=>x"6300", 279=>x"8a00", 280=>x"c500",
---- 281=>x"5500", 282=>x"7d00", 283=>x"9400", 284=>x"4900",
---- 285=>x"6800", 286=>x"8e00", 287=>x"9600", 288=>x"5d00",
---- 289=>x"8100", 290=>x"9500", 291=>x"9800", 292=>x"7700",
---- 293=>x"9000", 294=>x"9900", 295=>x"9500", 296=>x"8700",
---- 297=>x"9800", 298=>x"9800", 299=>x"9400", 300=>x"9300",
---- 301=>x"9800", 302=>x"9600", 303=>x"9000", 304=>x"9a00",
---- 305=>x"6800", 306=>x"9100", 307=>x"9100", 308=>x"9b00",
---- 309=>x"9400", 310=>x"9000", 311=>x"9300", 312=>x"9700",
---- 313=>x"9300", 314=>x"9100", 315=>x"9800", 316=>x"9300",
---- 317=>x"8e00", 318=>x"9300", 319=>x"9b00", 320=>x"9100",
---- 321=>x"9200", 322=>x"9600", 323=>x"9f00", 324=>x"9100",
---- 325=>x"9400", 326=>x"9d00", 327=>x"a000", 328=>x"9100",
---- 329=>x"9600", 330=>x"9c00", 331=>x"9f00", 332=>x"9500",
---- 333=>x"6200", 334=>x"9e00", 335=>x"9f00", 336=>x"9800",
---- 337=>x"9d00", 338=>x"9e00", 339=>x"9f00", 340=>x"9c00",
---- 341=>x"9f00", 342=>x"a000", 343=>x"a100", 344=>x"9c00",
---- 345=>x"a000", 346=>x"9e00", 347=>x"a200", 348=>x"a100",
---- 349=>x"9f00", 350=>x"9f00", 351=>x"a100", 352=>x"a200",
---- 353=>x"a100", 354=>x"9f00", 355=>x"9e00", 356=>x"a100",
---- 357=>x"a000", 358=>x"a200", 359=>x"a000", 360=>x"a100",
---- 361=>x"a000", 362=>x"a000", 363=>x"9f00", 364=>x"9f00",
---- 365=>x"a100", 366=>x"a000", 367=>x"9f00", 368=>x"a400",
---- 369=>x"a100", 370=>x"9f00", 371=>x"a300", 372=>x"a200",
---- 373=>x"a100", 374=>x"9e00", 375=>x"9f00", 376=>x"a200",
---- 377=>x"a300", 378=>x"9f00", 379=>x"a000", 380=>x"a000",
---- 381=>x"a200", 382=>x"a100", 383=>x"a200", 384=>x"a200",
---- 385=>x"5b00", 386=>x"a300", 387=>x"a100", 388=>x"a700",
---- 389=>x"a500", 390=>x"a200", 391=>x"a100", 392=>x"a600",
---- 393=>x"a300", 394=>x"a200", 395=>x"a200", 396=>x"a800",
---- 397=>x"a300", 398=>x"a300", 399=>x"a300", 400=>x"a500",
---- 401=>x"a500", 402=>x"a400", 403=>x"a300", 404=>x"a400",
---- 405=>x"a100", 406=>x"a100", 407=>x"a400", 408=>x"a400",
---- 409=>x"a200", 410=>x"a000", 411=>x"a400", 412=>x"a400",
---- 413=>x"a200", 414=>x"a100", 415=>x"a400", 416=>x"a400",
---- 417=>x"a300", 418=>x"a300", 419=>x"a400", 420=>x"a200",
---- 421=>x"a400", 422=>x"a400", 423=>x"a400", 424=>x"a200",
---- 425=>x"a300", 426=>x"a300", 427=>x"a400", 428=>x"a400",
---- 429=>x"a300", 430=>x"a200", 431=>x"a400", 432=>x"a200",
---- 433=>x"a100", 434=>x"a300", 435=>x"a300", 436=>x"a200",
---- 437=>x"a100", 438=>x"9e00", 439=>x"a100", 440=>x"a400",
---- 441=>x"a300", 442=>x"a100", 443=>x"a200", 444=>x"a200",
---- 445=>x"a300", 446=>x"a300", 447=>x"a300", 448=>x"a100",
---- 449=>x"9f00", 450=>x"9f00", 451=>x"a100", 452=>x"9a00",
---- 453=>x"9b00", 454=>x"9e00", 455=>x"a000", 456=>x"9800",
---- 457=>x"9700", 458=>x"9600", 459=>x"9900", 460=>x"9400",
---- 461=>x"9700", 462=>x"9600", 463=>x"9600", 464=>x"9600",
---- 465=>x"9700", 466=>x"9400", 467=>x"9300", 468=>x"9900",
---- 469=>x"9900", 470=>x"9900", 471=>x"9500", 472=>x"9d00",
---- 473=>x"9c00", 474=>x"9900", 475=>x"9b00", 476=>x"a000",
---- 477=>x"9e00", 478=>x"9b00", 479=>x"9c00", 480=>x"a500",
---- 481=>x"a000", 482=>x"9e00", 483=>x"9d00", 484=>x"a400",
---- 485=>x"a300", 486=>x"a000", 487=>x"9e00", 488=>x"a400",
---- 489=>x"a300", 490=>x"9f00", 491=>x"9d00", 492=>x"a200",
---- 493=>x"a200", 494=>x"a200", 495=>x"9d00", 496=>x"9e00",
---- 497=>x"a100", 498=>x"a100", 499=>x"9c00", 500=>x"9f00",
---- 501=>x"9f00", 502=>x"9f00", 503=>x"9b00", 504=>x"9d00",
---- 505=>x"9e00", 506=>x"9e00", 507=>x"9c00", 508=>x"9f00",
---- 509=>x"a000", 510=>x"6200", 511=>x"9b00", 512=>x"9e00",
---- 513=>x"9d00", 514=>x"9b00", 515=>x"9b00", 516=>x"9d00",
---- 517=>x"9d00", 518=>x"9e00", 519=>x"9a00", 520=>x"9c00",
---- 521=>x"9b00", 522=>x"9a00", 523=>x"9a00", 524=>x"9d00",
---- 525=>x"9a00", 526=>x"9a00", 527=>x"9800", 528=>x"6600",
---- 529=>x"9900", 530=>x"9a00", 531=>x"9a00", 532=>x"9800",
---- 533=>x"9800", 534=>x"9800", 535=>x"9a00", 536=>x"9a00",
---- 537=>x"6500", 538=>x"9800", 539=>x"9700", 540=>x"9a00",
---- 541=>x"9800", 542=>x"9900", 543=>x"9a00", 544=>x"9900",
---- 545=>x"9800", 546=>x"9800", 547=>x"9700", 548=>x"9700",
---- 549=>x"9600", 550=>x"9500", 551=>x"9600", 552=>x"9b00",
---- 553=>x"9800", 554=>x"9700", 555=>x"9500", 556=>x"9900",
---- 557=>x"9700", 558=>x"9700", 559=>x"9400", 560=>x"9700",
---- 561=>x"9500", 562=>x"9500", 563=>x"9400", 564=>x"9600",
---- 565=>x"9300", 566=>x"9200", 567=>x"9200", 568=>x"9300",
---- 569=>x"6d00", 570=>x"9100", 571=>x"9300", 572=>x"9200",
---- 573=>x"9400", 574=>x"9100", 575=>x"8f00", 576=>x"8f00",
---- 577=>x"8f00", 578=>x"8f00", 579=>x"8e00", 580=>x"8f00",
---- 581=>x"8e00", 582=>x"8e00", 583=>x"8c00", 584=>x"8f00",
---- 585=>x"8f00", 586=>x"8b00", 587=>x"8900", 588=>x"6f00",
---- 589=>x"9000", 590=>x"8d00", 591=>x"8a00", 592=>x"8f00",
---- 593=>x"8e00", 594=>x"8b00", 595=>x"8800", 596=>x"8d00",
---- 597=>x"7200", 598=>x"8a00", 599=>x"8800", 600=>x"8b00",
---- 601=>x"8a00", 602=>x"8500", 603=>x"8500", 604=>x"8e00",
---- 605=>x"8800", 606=>x"8500", 607=>x"8300", 608=>x"8a00",
---- 609=>x"8800", 610=>x"8500", 611=>x"8100", 612=>x"8b00",
---- 613=>x"8800", 614=>x"7d00", 615=>x"8200", 616=>x"8800",
---- 617=>x"8500", 618=>x"8100", 619=>x"8900", 620=>x"8700",
---- 621=>x"8500", 622=>x"8200", 623=>x"6c00", 624=>x"8600",
---- 625=>x"8200", 626=>x"8900", 627=>x"a300", 628=>x"8400",
---- 629=>x"8200", 630=>x"9600", 631=>x"af00", 632=>x"8200",
---- 633=>x"8800", 634=>x"a000", 635=>x"b800", 636=>x"8200",
---- 637=>x"9100", 638=>x"aa00", 639=>x"bc00", 640=>x"8500",
---- 641=>x"9e00", 642=>x"4c00", 643=>x"bf00", 644=>x"8800",
---- 645=>x"a400", 646=>x"b600", 647=>x"c000", 648=>x"9100",
---- 649=>x"aa00", 650=>x"bc00", 651=>x"c100", 652=>x"9a00",
---- 653=>x"af00", 654=>x"bf00", 655=>x"c400", 656=>x"a000",
---- 657=>x"b600", 658=>x"c100", 659=>x"c400", 660=>x"a500",
---- 661=>x"b900", 662=>x"c300", 663=>x"c400", 664=>x"a900",
---- 665=>x"bb00", 666=>x"c300", 667=>x"c400", 668=>x"ab00",
---- 669=>x"bd00", 670=>x"c400", 671=>x"c400", 672=>x"b100",
---- 673=>x"bf00", 674=>x"c400", 675=>x"c400", 676=>x"b500",
---- 677=>x"c200", 678=>x"c200", 679=>x"c500", 680=>x"b600",
---- 681=>x"c400", 682=>x"c500", 683=>x"c400", 684=>x"b700",
---- 685=>x"c300", 686=>x"c400", 687=>x"c600", 688=>x"b800",
---- 689=>x"c200", 690=>x"c600", 691=>x"ca00", 692=>x"b900",
---- 693=>x"c300", 694=>x"c700", 695=>x"cb00", 696=>x"ba00",
---- 697=>x"c300", 698=>x"ca00", 699=>x"ce00", 700=>x"bc00",
---- 701=>x"c600", 702=>x"cc00", 703=>x"d100", 704=>x"c000",
---- 705=>x"c900", 706=>x"cf00", 707=>x"d300", 708=>x"c400",
---- 709=>x"cc00", 710=>x"d200", 711=>x"2b00", 712=>x"c700",
---- 713=>x"cf00", 714=>x"d500", 715=>x"d400", 716=>x"ca00",
---- 717=>x"d300", 718=>x"d600", 719=>x"d600", 720=>x"cf00",
---- 721=>x"d400", 722=>x"d700", 723=>x"d700", 724=>x"cf00",
---- 725=>x"d600", 726=>x"d800", 727=>x"d700", 728=>x"d100",
---- 729=>x"d800", 730=>x"d900", 731=>x"d900", 732=>x"d300",
---- 733=>x"db00", 734=>x"dc00", 735=>x"d800", 736=>x"d500",
---- 737=>x"da00", 738=>x"da00", 739=>x"da00", 740=>x"d400",
---- 741=>x"db00", 742=>x"db00", 743=>x"db00", 744=>x"d500",
---- 745=>x"db00", 746=>x"da00", 747=>x"da00", 748=>x"d800",
---- 749=>x"dd00", 750=>x"da00", 751=>x"db00", 752=>x"da00",
---- 753=>x"2100", 754=>x"dc00", 755=>x"db00", 756=>x"dc00",
---- 757=>x"de00", 758=>x"db00", 759=>x"d900", 760=>x"dd00",
---- 761=>x"df00", 762=>x"db00", 763=>x"d700", 764=>x"dc00",
---- 765=>x"dd00", 766=>x"da00", 767=>x"d800", 768=>x"dd00",
---- 769=>x"dc00", 770=>x"d800", 771=>x"d700", 772=>x"db00",
---- 773=>x"da00", 774=>x"d600", 775=>x"d400", 776=>x"db00",
---- 777=>x"d700", 778=>x"d200", 779=>x"d200", 780=>x"d900",
---- 781=>x"d200", 782=>x"d000", 783=>x"d200", 784=>x"d600",
---- 785=>x"cf00", 786=>x"cf00", 787=>x"d000", 788=>x"d400",
---- 789=>x"ce00", 790=>x"cd00", 791=>x"ce00", 792=>x"ce00",
---- 793=>x"cc00", 794=>x"cc00", 795=>x"ce00", 796=>x"cf00",
---- 797=>x"cb00", 798=>x"cc00", 799=>x"cf00", 800=>x"cd00",
---- 801=>x"cc00", 802=>x"cd00", 803=>x"d100", 804=>x"cd00",
---- 805=>x"cc00", 806=>x"d000", 807=>x"d400", 808=>x"d000",
---- 809=>x"cf00", 810=>x"d400", 811=>x"d600", 812=>x"d300",
---- 813=>x"d200", 814=>x"d300", 815=>x"d700", 816=>x"d400",
---- 817=>x"d400", 818=>x"d300", 819=>x"d500", 820=>x"d400",
---- 821=>x"d400", 822=>x"d400", 823=>x"d500", 824=>x"d400",
---- 825=>x"d500", 826=>x"d500", 827=>x"d500", 828=>x"d500",
---- 829=>x"d600", 830=>x"d600", 831=>x"d500", 832=>x"d600",
---- 833=>x"d500", 834=>x"d400", 835=>x"d400", 836=>x"d500",
---- 837=>x"d400", 838=>x"d500", 839=>x"d200", 840=>x"d700",
---- 841=>x"d400", 842=>x"d200", 843=>x"d200", 844=>x"d500",
---- 845=>x"d300", 846=>x"d200", 847=>x"d000", 848=>x"d500",
---- 849=>x"d500", 850=>x"d000", 851=>x"cc00", 852=>x"d600",
---- 853=>x"d100", 854=>x"cf00", 855=>x"3900", 856=>x"d500",
---- 857=>x"cf00", 858=>x"cb00", 859=>x"bd00", 860=>x"d600",
---- 861=>x"d000", 862=>x"c500", 863=>x"ab00", 864=>x"d300",
---- 865=>x"cb00", 866=>x"bb00", 867=>x"9900", 868=>x"cf00",
---- 869=>x"c400", 870=>x"ac00", 871=>x"8600", 872=>x"ce00",
---- 873=>x"bb00", 874=>x"9b00", 875=>x"7700", 876=>x"c800",
---- 877=>x"ad00", 878=>x"8d00", 879=>x"7200", 880=>x"bc00",
---- 881=>x"9e00", 882=>x"8300", 883=>x"7200", 884=>x"ad00",
---- 885=>x"8d00", 886=>x"7800", 887=>x"7800", 888=>x"9d00",
---- 889=>x"8200", 890=>x"7600", 891=>x"7800", 892=>x"9000",
---- 893=>x"7900", 894=>x"7100", 895=>x"8900", 896=>x"8500",
---- 897=>x"7800", 898=>x"7500", 899=>x"7300", 900=>x"7c00",
---- 901=>x"7500", 902=>x"7500", 903=>x"7000", 904=>x"7b00",
---- 905=>x"7100", 906=>x"6f00", 907=>x"7000", 908=>x"7900",
---- 909=>x"6e00", 910=>x"6c00", 911=>x"6a00", 912=>x"7400",
---- 913=>x"7000", 914=>x"6d00", 915=>x"6400", 916=>x"7200",
---- 917=>x"6f00", 918=>x"6a00", 919=>x"6600", 920=>x"7000",
---- 921=>x"6c00", 922=>x"6400", 923=>x"5e00", 924=>x"6b00",
---- 925=>x"6200", 926=>x"5700", 927=>x"4f00", 928=>x"5f00",
---- 929=>x"5900", 930=>x"4f00", 931=>x"4b00", 932=>x"5500",
---- 933=>x"4e00", 934=>x"4a00", 935=>x"4e00", 936=>x"4700",
---- 937=>x"3e00", 938=>x"4400", 939=>x"5000", 940=>x"3a00",
---- 941=>x"3900", 942=>x"4c00", 943=>x"5100", 944=>x"3800",
---- 945=>x"4100", 946=>x"4d00", 947=>x"5200", 948=>x"4200",
---- 949=>x"4d00", 950=>x"4f00", 951=>x"5300", 952=>x"4500",
---- 953=>x"4c00", 954=>x"4f00", 955=>x"4c00", 956=>x"4b00",
---- 957=>x"4a00", 958=>x"4400", 959=>x"4500", 960=>x"4c00",
---- 961=>x"4600", 962=>x"4100", 963=>x"4a00", 964=>x"4100",
---- 965=>x"4000", 966=>x"4900", 967=>x"5600", 968=>x"c000",
---- 969=>x"4500", 970=>x"4f00", 971=>x"5b00", 972=>x"4600",
---- 973=>x"5100", 974=>x"5b00", 975=>x"6700", 976=>x"5100",
---- 977=>x"6000", 978=>x"6b00", 979=>x"6f00", 980=>x"5c00",
---- 981=>x"6800", 982=>x"7200", 983=>x"6c00", 984=>x"6300",
---- 985=>x"6900", 986=>x"6e00", 987=>x"6200", 988=>x"6800",
---- 989=>x"6900", 990=>x"6300", 991=>x"5a00", 992=>x"6900",
---- 993=>x"6400", 994=>x"5700", 995=>x"5400", 996=>x"5900",
---- 997=>x"5400", 998=>x"5000", 999=>x"4700", 1000=>x"5400",
---- 1001=>x"4a00", 1002=>x"4500", 1003=>x"4300", 1004=>x"4f00",
---- 1005=>x"4700", 1006=>x"4500", 1007=>x"4800", 1008=>x"5100",
---- 1009=>x"5200", 1010=>x"4c00", 1011=>x"5000", 1012=>x"5600",
---- 1013=>x"5500", 1014=>x"5200", 1015=>x"4f00", 1016=>x"5800",
---- 1017=>x"5700", 1018=>x"5400", 1019=>x"5300", 1020=>x"5b00",
---- 1021=>x"5a00", 1022=>x"5600", 1023=>x"5300"),
----
---- 58 => (0=>x"7b00", 1=>x"7d00", 2=>x"7a00", 3=>x"7d00", 4=>x"7b00",
---- 5=>x"7c00", 6=>x"7a00", 7=>x"7d00", 8=>x"7c00",
---- 9=>x"7c00", 10=>x"7b00", 11=>x"7c00", 12=>x"7d00",
---- 13=>x"7d00", 14=>x"7d00", 15=>x"7b00", 16=>x"7e00",
---- 17=>x"7b00", 18=>x"7c00", 19=>x"7c00", 20=>x"7900",
---- 21=>x"7b00", 22=>x"7b00", 23=>x"7900", 24=>x"7b00",
---- 25=>x"7900", 26=>x"7a00", 27=>x"7900", 28=>x"7a00",
---- 29=>x"7700", 30=>x"7a00", 31=>x"7b00", 32=>x"7a00",
---- 33=>x"7b00", 34=>x"7c00", 35=>x"7c00", 36=>x"7a00",
---- 37=>x"7e00", 38=>x"7b00", 39=>x"7c00", 40=>x"7800",
---- 41=>x"7a00", 42=>x"7a00", 43=>x"8000", 44=>x"7a00",
---- 45=>x"7900", 46=>x"7e00", 47=>x"8000", 48=>x"7800",
---- 49=>x"7800", 50=>x"7900", 51=>x"7e00", 52=>x"8800",
---- 53=>x"7b00", 54=>x"7b00", 55=>x"7a00", 56=>x"7800",
---- 57=>x"7900", 58=>x"7b00", 59=>x"7d00", 60=>x"7900",
---- 61=>x"7b00", 62=>x"7a00", 63=>x"7e00", 64=>x"7d00",
---- 65=>x"7c00", 66=>x"7c00", 67=>x"7f00", 68=>x"7a00",
---- 69=>x"7f00", 70=>x"7f00", 71=>x"8200", 72=>x"7b00",
---- 73=>x"8100", 74=>x"8400", 75=>x"8600", 76=>x"7e00",
---- 77=>x"8100", 78=>x"7900", 79=>x"8100", 80=>x"7d00",
---- 81=>x"8200", 82=>x"8200", 83=>x"6e00", 84=>x"8200",
---- 85=>x"8100", 86=>x"6e00", 87=>x"4e00", 88=>x"8100",
---- 89=>x"6f00", 90=>x"4c00", 91=>x"3000", 92=>x"6700",
---- 93=>x"4a00", 94=>x"3200", 95=>x"2b00", 96=>x"4900",
---- 97=>x"2a00", 98=>x"2b00", 99=>x"2b00", 100=>x"2e00",
---- 101=>x"2800", 102=>x"2a00", 103=>x"2c00", 104=>x"2800",
---- 105=>x"2700", 106=>x"2b00", 107=>x"2a00", 108=>x"2c00",
---- 109=>x"2a00", 110=>x"2e00", 111=>x"3000", 112=>x"2900",
---- 113=>x"2a00", 114=>x"3100", 115=>x"2d00", 116=>x"2e00",
---- 117=>x"2a00", 118=>x"2e00", 119=>x"2b00", 120=>x"2d00",
---- 121=>x"3000", 122=>x"3000", 123=>x"2d00", 124=>x"2c00",
---- 125=>x"2e00", 126=>x"2f00", 127=>x"3200", 128=>x"2f00",
---- 129=>x"2e00", 130=>x"3100", 131=>x"3500", 132=>x"2e00",
---- 133=>x"3100", 134=>x"3500", 135=>x"3a00", 136=>x"2e00",
---- 137=>x"3400", 138=>x"3400", 139=>x"3300", 140=>x"3100",
---- 141=>x"3200", 142=>x"3100", 143=>x"3200", 144=>x"3200",
---- 145=>x"3100", 146=>x"cd00", 147=>x"3600", 148=>x"3b00",
---- 149=>x"3600", 150=>x"cc00", 151=>x"3100", 152=>x"3500",
---- 153=>x"3800", 154=>x"3600", 155=>x"3200", 156=>x"3500",
---- 157=>x"3200", 158=>x"2c00", 159=>x"2c00", 160=>x"3500",
---- 161=>x"3300", 162=>x"3100", 163=>x"2e00", 164=>x"3500",
---- 165=>x"3200", 166=>x"2d00", 167=>x"2c00", 168=>x"3000",
---- 169=>x"2d00", 170=>x"2a00", 171=>x"2f00", 172=>x"2f00",
---- 173=>x"2700", 174=>x"2c00", 175=>x"3400", 176=>x"2d00",
---- 177=>x"2a00", 178=>x"3500", 179=>x"3c00", 180=>x"2d00",
---- 181=>x"3000", 182=>x"3800", 183=>x"3a00", 184=>x"2e00",
---- 185=>x"3800", 186=>x"3c00", 187=>x"3300", 188=>x"3400",
---- 189=>x"3a00", 190=>x"3e00", 191=>x"2f00", 192=>x"3900",
---- 193=>x"3a00", 194=>x"2e00", 195=>x"2b00", 196=>x"3c00",
---- 197=>x"3200", 198=>x"2d00", 199=>x"2d00", 200=>x"3500",
---- 201=>x"2c00", 202=>x"3100", 203=>x"2f00", 204=>x"3000",
---- 205=>x"2c00", 206=>x"3700", 207=>x"3400", 208=>x"d600",
---- 209=>x"d300", 210=>x"3300", 211=>x"3500", 212=>x"2e00",
---- 213=>x"3300", 214=>x"3600", 215=>x"3100", 216=>x"3400",
---- 217=>x"3700", 218=>x"3b00", 219=>x"3500", 220=>x"3500",
---- 221=>x"3b00", 222=>x"3500", 223=>x"3000", 224=>x"3800",
---- 225=>x"3500", 226=>x"3200", 227=>x"2f00", 228=>x"3700",
---- 229=>x"2f00", 230=>x"2900", 231=>x"2d00", 232=>x"3500",
---- 233=>x"2900", 234=>x"d800", 235=>x"2b00", 236=>x"3700",
---- 237=>x"2d00", 238=>x"2900", 239=>x"3000", 240=>x"3200",
---- 241=>x"2c00", 242=>x"3200", 243=>x"4c00", 244=>x"2f00",
---- 245=>x"3100", 246=>x"4100", 247=>x"6b00", 248=>x"3100",
---- 249=>x"3700", 250=>x"5a00", 251=>x"8300", 252=>x"2f00",
---- 253=>x"4700", 254=>x"7500", 255=>x"9300", 256=>x"3800",
---- 257=>x"6400", 258=>x"8d00", 259=>x"9b00", 260=>x"4c00",
---- 261=>x"8100", 262=>x"9a00", 263=>x"9b00", 264=>x"6e00",
---- 265=>x"9200", 266=>x"9a00", 267=>x"9600", 268=>x"8700",
---- 269=>x"9900", 270=>x"9b00", 271=>x"9600", 272=>x"9200",
---- 273=>x"9c00", 274=>x"9900", 275=>x"9400", 276=>x"9800",
---- 277=>x"9a00", 278=>x"9600", 279=>x"9000", 280=>x"6400",
---- 281=>x"9500", 282=>x"9300", 283=>x"9200", 284=>x"9500",
---- 285=>x"9200", 286=>x"9100", 287=>x"9500", 288=>x"9400",
---- 289=>x"8f00", 290=>x"9300", 291=>x"9800", 292=>x"9100",
---- 293=>x"9200", 294=>x"9700", 295=>x"9c00", 296=>x"9000",
---- 297=>x"9400", 298=>x"9b00", 299=>x"9f00", 300=>x"8f00",
---- 301=>x"9500", 302=>x"9f00", 303=>x"a000", 304=>x"9600",
---- 305=>x"9c00", 306=>x"a000", 307=>x"a000", 308=>x"9c00",
---- 309=>x"a000", 310=>x"a000", 311=>x"a000", 312=>x"9c00",
---- 313=>x"9f00", 314=>x"a000", 315=>x"a200", 316=>x"9e00",
---- 317=>x"9f00", 318=>x"a200", 319=>x"a000", 320=>x"a000",
---- 321=>x"a100", 322=>x"a100", 323=>x"a100", 324=>x"9f00",
---- 325=>x"a200", 326=>x"a000", 327=>x"a200", 328=>x"a000",
---- 329=>x"a100", 330=>x"a000", 331=>x"9e00", 332=>x"a100",
---- 333=>x"a000", 334=>x"9e00", 335=>x"9d00", 336=>x"9f00",
---- 337=>x"9f00", 338=>x"9d00", 339=>x"9d00", 340=>x"9f00",
---- 341=>x"9e00", 342=>x"9e00", 343=>x"9e00", 344=>x"a000",
---- 345=>x"9e00", 346=>x"a000", 347=>x"9c00", 348=>x"9e00",
---- 349=>x"9f00", 350=>x"9e00", 351=>x"9c00", 352=>x"9f00",
---- 353=>x"9f00", 354=>x"9f00", 355=>x"9f00", 356=>x"9f00",
---- 357=>x"9e00", 358=>x"9f00", 359=>x"9e00", 360=>x"9f00",
---- 361=>x"9f00", 362=>x"a000", 363=>x"9d00", 364=>x"9f00",
---- 365=>x"a000", 366=>x"a200", 367=>x"9f00", 368=>x"a200",
---- 369=>x"9f00", 370=>x"a000", 371=>x"9f00", 372=>x"a000",
---- 373=>x"a000", 374=>x"9f00", 375=>x"9f00", 376=>x"a200",
---- 377=>x"a000", 378=>x"a100", 379=>x"9e00", 380=>x"a100",
---- 381=>x"9f00", 382=>x"9f00", 383=>x"9e00", 384=>x"a400",
---- 385=>x"a300", 386=>x"a100", 387=>x"a000", 388=>x"a200",
---- 389=>x"a100", 390=>x"a100", 391=>x"a000", 392=>x"a200",
---- 393=>x"a100", 394=>x"a200", 395=>x"9f00", 396=>x"a200",
---- 397=>x"a300", 398=>x"a200", 399=>x"a000", 400=>x"a200",
---- 401=>x"5c00", 402=>x"a200", 403=>x"a100", 404=>x"a400",
---- 405=>x"a300", 406=>x"a200", 407=>x"a200", 408=>x"a200",
---- 409=>x"a200", 410=>x"a300", 411=>x"a200", 412=>x"a500",
---- 413=>x"a400", 414=>x"a300", 415=>x"5e00", 416=>x"a400",
---- 417=>x"a100", 418=>x"a100", 419=>x"a200", 420=>x"a100",
---- 421=>x"a100", 422=>x"9f00", 423=>x"a300", 424=>x"a400",
---- 425=>x"a200", 426=>x"a100", 427=>x"a400", 428=>x"a400",
---- 429=>x"a500", 430=>x"a300", 431=>x"a000", 432=>x"a300",
---- 433=>x"a200", 434=>x"a300", 435=>x"a400", 436=>x"a400",
---- 437=>x"a100", 438=>x"a300", 439=>x"a400", 440=>x"a100",
---- 441=>x"a200", 442=>x"a000", 443=>x"a300", 444=>x"a000",
---- 445=>x"a100", 446=>x"a100", 447=>x"a200", 448=>x"a100",
---- 449=>x"a100", 450=>x"a000", 451=>x"a200", 452=>x"a100",
---- 453=>x"a000", 454=>x"a200", 455=>x"5e00", 456=>x"9a00",
---- 457=>x"9a00", 458=>x"9d00", 459=>x"9f00", 460=>x"9400",
---- 461=>x"9200", 462=>x"9600", 463=>x"9800", 464=>x"9200",
---- 465=>x"9200", 466=>x"9300", 467=>x"9200", 468=>x"9400",
---- 469=>x"9100", 470=>x"9200", 471=>x"9100", 472=>x"9900",
---- 473=>x"9200", 474=>x"9100", 475=>x"9000", 476=>x"9900",
---- 477=>x"9500", 478=>x"9300", 479=>x"9100", 480=>x"9a00",
---- 481=>x"9700", 482=>x"9400", 483=>x"9400", 484=>x"9c00",
---- 485=>x"9d00", 486=>x"9800", 487=>x"9700", 488=>x"9d00",
---- 489=>x"9e00", 490=>x"9b00", 491=>x"9d00", 492=>x"9900",
---- 493=>x"9900", 494=>x"9b00", 495=>x"9d00", 496=>x"9800",
---- 497=>x"9a00", 498=>x"9c00", 499=>x"9b00", 500=>x"9b00",
---- 501=>x"9b00", 502=>x"9a00", 503=>x"9a00", 504=>x"9c00",
---- 505=>x"9a00", 506=>x"9900", 507=>x"9700", 508=>x"9a00",
---- 509=>x"9c00", 510=>x"9a00", 511=>x"9900", 512=>x"9a00",
---- 513=>x"9900", 514=>x"9800", 515=>x"9800", 516=>x"9900",
---- 517=>x"9800", 518=>x"9a00", 519=>x"9800", 520=>x"9a00",
---- 521=>x"9900", 522=>x"9900", 523=>x"9900", 524=>x"9900",
---- 525=>x"9700", 526=>x"9b00", 527=>x"9c00", 528=>x"9900",
---- 529=>x"9800", 530=>x"9900", 531=>x"9a00", 532=>x"9900",
---- 533=>x"9800", 534=>x"9700", 535=>x"9800", 536=>x"9800",
---- 537=>x"9700", 538=>x"9600", 539=>x"9400", 540=>x"9600",
---- 541=>x"9700", 542=>x"9600", 543=>x"9100", 544=>x"9600",
---- 545=>x"9800", 546=>x"9700", 547=>x"9200", 548=>x"9600",
---- 549=>x"9300", 550=>x"9400", 551=>x"9200", 552=>x"9200",
---- 553=>x"9300", 554=>x"9400", 555=>x"8e00", 556=>x"9000",
---- 557=>x"8e00", 558=>x"9100", 559=>x"8d00", 560=>x"9100",
---- 561=>x"9200", 562=>x"9000", 563=>x"8b00", 564=>x"9000",
---- 565=>x"8e00", 566=>x"8f00", 567=>x"8d00", 568=>x"8e00",
---- 569=>x"8e00", 570=>x"8c00", 571=>x"8d00", 572=>x"8f00",
---- 573=>x"8e00", 574=>x"8f00", 575=>x"8a00", 576=>x"8c00",
---- 577=>x"8c00", 578=>x"8900", 579=>x"8600", 580=>x"8b00",
---- 581=>x"8900", 582=>x"8700", 583=>x"8700", 584=>x"8900",
---- 585=>x"8600", 586=>x"8600", 587=>x"8400", 588=>x"8700",
---- 589=>x"8400", 590=>x"8300", 591=>x"8600", 592=>x"8600",
---- 593=>x"8200", 594=>x"8300", 595=>x"9300", 596=>x"8400",
---- 597=>x"7d00", 598=>x"8a00", 599=>x"a200", 600=>x"8200",
---- 601=>x"8000", 602=>x"9800", 603=>x"af00", 604=>x"8100",
---- 605=>x"9000", 606=>x"a800", 607=>x"bb00", 608=>x"8600",
---- 609=>x"9d00", 610=>x"b300", 611=>x"be00", 612=>x"9200",
---- 613=>x"ac00", 614=>x"bb00", 615=>x"c200", 616=>x"a000",
---- 617=>x"b700", 618=>x"bf00", 619=>x"c300", 620=>x"ad00",
---- 621=>x"bc00", 622=>x"c300", 623=>x"c400", 624=>x"b600",
---- 625=>x"c000", 626=>x"c500", 627=>x"c400", 628=>x"be00",
---- 629=>x"c500", 630=>x"c500", 631=>x"c300", 632=>x"c200",
---- 633=>x"c600", 634=>x"c300", 635=>x"c300", 636=>x"c400",
---- 637=>x"c600", 638=>x"c400", 639=>x"c300", 640=>x"c700",
---- 641=>x"c300", 642=>x"c200", 643=>x"c200", 644=>x"c500",
---- 645=>x"3a00", 646=>x"c100", 647=>x"c200", 648=>x"c500",
---- 649=>x"c300", 650=>x"c500", 651=>x"c400", 652=>x"c400",
---- 653=>x"c400", 654=>x"c400", 655=>x"c300", 656=>x"c400",
---- 657=>x"c500", 658=>x"c400", 659=>x"c500", 660=>x"c400",
---- 661=>x"c400", 662=>x"c500", 663=>x"c800", 664=>x"c300",
---- 665=>x"c400", 666=>x"3a00", 667=>x"c900", 668=>x"c300",
---- 669=>x"c500", 670=>x"c700", 671=>x"cc00", 672=>x"c400",
---- 673=>x"c700", 674=>x"ca00", 675=>x"ce00", 676=>x"c500",
---- 677=>x"c900", 678=>x"cc00", 679=>x"d100", 680=>x"c600",
---- 681=>x"cc00", 682=>x"ce00", 683=>x"2e00", 684=>x"cb00",
---- 685=>x"ce00", 686=>x"d100", 687=>x"cf00", 688=>x"cc00",
---- 689=>x"cf00", 690=>x"d300", 691=>x"d300", 692=>x"cd00",
---- 693=>x"d100", 694=>x"d300", 695=>x"d100", 696=>x"cf00",
---- 697=>x"d400", 698=>x"d100", 699=>x"d200", 700=>x"d300",
---- 701=>x"d400", 702=>x"d400", 703=>x"d200", 704=>x"d500",
---- 705=>x"d400", 706=>x"d300", 707=>x"d300", 708=>x"d400",
---- 709=>x"d400", 710=>x"d200", 711=>x"d200", 712=>x"d400",
---- 713=>x"d400", 714=>x"d300", 715=>x"d200", 716=>x"2b00",
---- 717=>x"d300", 718=>x"d500", 719=>x"d200", 720=>x"d600",
---- 721=>x"d500", 722=>x"d500", 723=>x"d300", 724=>x"d500",
---- 725=>x"d300", 726=>x"d500", 727=>x"d400", 728=>x"d600",
---- 729=>x"2a00", 730=>x"d600", 731=>x"d500", 732=>x"d500",
---- 733=>x"d700", 734=>x"d700", 735=>x"d500", 736=>x"d700",
---- 737=>x"d400", 738=>x"d800", 739=>x"d700", 740=>x"d700",
---- 741=>x"d700", 742=>x"d700", 743=>x"d900", 744=>x"d900",
---- 745=>x"d600", 746=>x"d600", 747=>x"d600", 748=>x"d900",
---- 749=>x"d500", 750=>x"d500", 751=>x"d400", 752=>x"d600",
---- 753=>x"d400", 754=>x"d400", 755=>x"d200", 756=>x"d500",
---- 757=>x"d300", 758=>x"d300", 759=>x"d300", 760=>x"d400",
---- 761=>x"d200", 762=>x"d400", 763=>x"d400", 764=>x"d300",
---- 765=>x"d200", 766=>x"d500", 767=>x"d500", 768=>x"d300",
---- 769=>x"d400", 770=>x"d500", 771=>x"d400", 772=>x"d300",
---- 773=>x"d400", 774=>x"d200", 775=>x"d300", 776=>x"d200",
---- 777=>x"d200", 778=>x"d200", 779=>x"d200", 780=>x"d200",
---- 781=>x"d000", 782=>x"2a00", 783=>x"d100", 784=>x"3000",
---- 785=>x"d200", 786=>x"d200", 787=>x"d000", 788=>x"cf00",
---- 789=>x"d100", 790=>x"d100", 791=>x"d000", 792=>x"d000",
---- 793=>x"d100", 794=>x"d200", 795=>x"d000", 796=>x"cf00",
---- 797=>x"cf00", 798=>x"d100", 799=>x"d000", 800=>x"d100",
---- 801=>x"d000", 802=>x"d000", 803=>x"cf00", 804=>x"d200",
---- 805=>x"cf00", 806=>x"cf00", 807=>x"ce00", 808=>x"d300",
---- 809=>x"d100", 810=>x"d000", 811=>x"ce00", 812=>x"d300",
---- 813=>x"d100", 814=>x"cf00", 815=>x"cd00", 816=>x"d300",
---- 817=>x"ce00", 818=>x"cc00", 819=>x"c500", 820=>x"d100",
---- 821=>x"cb00", 822=>x"c500", 823=>x"ba00", 824=>x"d100",
---- 825=>x"c900", 826=>x"bd00", 827=>x"a900", 828=>x"d000",
---- 829=>x"c500", 830=>x"b400", 831=>x"9700", 832=>x"ce00",
---- 833=>x"c100", 834=>x"a500", 835=>x"8500", 836=>x"cb00",
---- 837=>x"bc00", 838=>x"9700", 839=>x"6b00", 840=>x"c700",
---- 841=>x"b300", 842=>x"8300", 843=>x"5400", 844=>x"c700",
---- 845=>x"a400", 846=>x"6f00", 847=>x"4c00", 848=>x"ba00",
---- 849=>x"9100", 850=>x"6100", 851=>x"5100", 852=>x"ac00",
---- 853=>x"7c00", 854=>x"5700", 855=>x"5a00", 856=>x"9600",
---- 857=>x"6500", 858=>x"5900", 859=>x"5b00", 860=>x"8200",
---- 861=>x"5e00", 862=>x"5900", 863=>x"5d00", 864=>x"7200",
---- 865=>x"5b00", 866=>x"5b00", 867=>x"5f00", 868=>x"6700",
---- 869=>x"5e00", 870=>x"5e00", 871=>x"5b00", 872=>x"6200",
---- 873=>x"6200", 874=>x"5e00", 875=>x"5900", 876=>x"6900",
---- 877=>x"6600", 878=>x"6400", 879=>x"5e00", 880=>x"6b00",
---- 881=>x"6900", 882=>x"6700", 883=>x"6200", 884=>x"7100",
---- 885=>x"6700", 886=>x"6000", 887=>x"5f00", 888=>x"7100",
---- 889=>x"6900", 890=>x"6400", 891=>x"6200", 892=>x"7000",
---- 893=>x"6700", 894=>x"6900", 895=>x"6000", 896=>x"7100",
---- 897=>x"6a00", 898=>x"6600", 899=>x"5d00", 900=>x"6e00",
---- 901=>x"6c00", 902=>x"6500", 903=>x"5d00", 904=>x"6a00",
---- 905=>x"6700", 906=>x"6000", 907=>x"5d00", 908=>x"6600",
---- 909=>x"6000", 910=>x"5a00", 911=>x"5e00", 912=>x"6100",
---- 913=>x"5c00", 914=>x"5900", 915=>x"6000", 916=>x"6000",
---- 917=>x"5900", 918=>x"5c00", 919=>x"6300", 920=>x"5700",
---- 921=>x"a700", 922=>x"6000", 923=>x"6600", 924=>x"5100",
---- 925=>x"5a00", 926=>x"6300", 927=>x"6100", 928=>x"5400",
---- 929=>x"6000", 930=>x"6200", 931=>x"5a00", 932=>x"5a00",
---- 933=>x"6000", 934=>x"5d00", 935=>x"5100", 936=>x"5a00",
---- 937=>x"5700", 938=>x"5200", 939=>x"4c00", 940=>x"5400",
---- 941=>x"4a00", 942=>x"4d00", 943=>x"ad00", 944=>x"4f00",
---- 945=>x"4b00", 946=>x"4e00", 947=>x"5d00", 948=>x"4900",
---- 949=>x"4300", 950=>x"4f00", 951=>x"5e00", 952=>x"4600",
---- 953=>x"4c00", 954=>x"5a00", 955=>x"6600", 956=>x"4a00",
---- 957=>x"5a00", 958=>x"6600", 959=>x"6d00", 960=>x"5200",
---- 961=>x"6100", 962=>x"6c00", 963=>x"6900", 964=>x"6000",
---- 965=>x"6600", 966=>x"6800", 967=>x"5f00", 968=>x"6900",
---- 969=>x"6c00", 970=>x"6600", 971=>x"5d00", 972=>x"6a00",
---- 973=>x"6700", 974=>x"6200", 975=>x"5700", 976=>x"6a00",
---- 977=>x"6000", 978=>x"5700", 979=>x"4f00", 980=>x"6200",
---- 981=>x"5700", 982=>x"4c00", 983=>x"4f00", 984=>x"5700",
---- 985=>x"4d00", 986=>x"4600", 987=>x"4500", 988=>x"4f00",
---- 989=>x"4800", 990=>x"4500", 991=>x"4100", 992=>x"4f00",
---- 993=>x"4f00", 994=>x"4800", 995=>x"4200", 996=>x"4b00",
---- 997=>x"4b00", 998=>x"4800", 999=>x"4700", 1000=>x"4900",
---- 1001=>x"4700", 1002=>x"4b00", 1003=>x"4800", 1004=>x"4800",
---- 1005=>x"4800", 1006=>x"4b00", 1007=>x"4f00", 1008=>x"4d00",
---- 1009=>x"4a00", 1010=>x"5000", 1011=>x"5900", 1012=>x"4b00",
---- 1013=>x"5000", 1014=>x"5b00", 1015=>x"6900", 1016=>x"4f00",
---- 1017=>x"5800", 1018=>x"6600", 1019=>x"7000", 1020=>x"5300",
---- 1021=>x"5e00", 1022=>x"6500", 1023=>x"7600"),
----
---- 59 => (0=>x"7e00", 1=>x"7c00", 2=>x"7c00", 3=>x"7700", 4=>x"7d00",
---- 5=>x"7c00", 6=>x"7d00", 7=>x"7700", 8=>x"7e00",
---- 9=>x"7c00", 10=>x"7e00", 11=>x"7600", 12=>x"7d00",
---- 13=>x"7a00", 14=>x"7c00", 15=>x"7900", 16=>x"7a00",
---- 17=>x"7a00", 18=>x"7b00", 19=>x"7d00", 20=>x"7b00",
---- 21=>x"7c00", 22=>x"7b00", 23=>x"7d00", 24=>x"7b00",
---- 25=>x"7b00", 26=>x"7b00", 27=>x"7900", 28=>x"7b00",
---- 29=>x"7e00", 30=>x"7e00", 31=>x"7b00", 32=>x"7a00",
---- 33=>x"7d00", 34=>x"8100", 35=>x"7d00", 36=>x"7d00",
---- 37=>x"7c00", 38=>x"8000", 39=>x"7e00", 40=>x"8000",
---- 41=>x"7f00", 42=>x"8000", 43=>x"8200", 44=>x"8100",
---- 45=>x"8300", 46=>x"8000", 47=>x"8300", 48=>x"7d00",
---- 49=>x"7e00", 50=>x"8100", 51=>x"8400", 52=>x"7b00",
---- 53=>x"7e00", 54=>x"8300", 55=>x"8500", 56=>x"7e00",
---- 57=>x"8100", 58=>x"8300", 59=>x"8a00", 60=>x"7f00",
---- 61=>x"8300", 62=>x"8600", 63=>x"8100", 64=>x"8100",
---- 65=>x"8300", 66=>x"8500", 67=>x"7300", 68=>x"8700",
---- 69=>x"8400", 70=>x"7000", 71=>x"4900", 72=>x"8200",
---- 73=>x"6d00", 74=>x"4a00", 75=>x"2a00", 76=>x"6c00",
---- 77=>x"4700", 78=>x"2b00", 79=>x"2c00", 80=>x"4a00",
---- 81=>x"3000", 82=>x"2800", 83=>x"2e00", 84=>x"2f00",
---- 85=>x"2b00", 86=>x"2a00", 87=>x"2b00", 88=>x"2c00",
---- 89=>x"2a00", 90=>x"2d00", 91=>x"2b00", 92=>x"2f00",
---- 93=>x"3100", 94=>x"2c00", 95=>x"2d00", 96=>x"2b00",
---- 97=>x"2e00", 98=>x"2b00", 99=>x"3000", 100=>x"d300",
---- 101=>x"2c00", 102=>x"2c00", 103=>x"2e00", 104=>x"2d00",
---- 105=>x"2e00", 106=>x"2c00", 107=>x"2e00", 108=>x"2f00",
---- 109=>x"3200", 110=>x"3100", 111=>x"3600", 112=>x"3400",
---- 113=>x"3500", 114=>x"3600", 115=>x"3500", 116=>x"3300",
---- 117=>x"3700", 118=>x"3500", 119=>x"3400", 120=>x"3200",
---- 121=>x"3700", 122=>x"3400", 123=>x"3100", 124=>x"3600",
---- 125=>x"3700", 126=>x"3500", 127=>x"3600", 128=>x"3700",
---- 129=>x"3200", 130=>x"3400", 131=>x"3900", 132=>x"3600",
---- 133=>x"3700", 134=>x"3800", 135=>x"3800", 136=>x"3300",
---- 137=>x"3700", 138=>x"3800", 139=>x"3400", 140=>x"3600",
---- 141=>x"cb00", 142=>x"3600", 143=>x"2f00", 144=>x"3500",
---- 145=>x"3500", 146=>x"2f00", 147=>x"d700", 148=>x"2e00",
---- 149=>x"2d00", 150=>x"2600", 151=>x"2a00", 152=>x"2c00",
---- 153=>x"2d00", 154=>x"2e00", 155=>x"3200", 156=>x"2c00",
---- 157=>x"2d00", 158=>x"3300", 159=>x"3900", 160=>x"2a00",
---- 161=>x"3000", 162=>x"3700", 163=>x"3b00", 164=>x"2b00",
---- 165=>x"3700", 166=>x"3b00", 167=>x"3700", 168=>x"2f00",
---- 169=>x"3600", 170=>x"3500", 171=>x"2e00", 172=>x"3800",
---- 173=>x"3700", 174=>x"2f00", 175=>x"2d00", 176=>x"3700",
---- 177=>x"3000", 178=>x"2b00", 179=>x"2c00", 180=>x"3300",
---- 181=>x"2e00", 182=>x"2e00", 183=>x"3100", 184=>x"2f00",
---- 185=>x"3100", 186=>x"3300", 187=>x"3400", 188=>x"2d00",
---- 189=>x"3200", 190=>x"3400", 191=>x"3100", 192=>x"3300",
---- 193=>x"3400", 194=>x"3500", 195=>x"3600", 196=>x"3600",
---- 197=>x"3500", 198=>x"3600", 199=>x"3700", 200=>x"3400",
---- 201=>x"3700", 202=>x"3600", 203=>x"3600", 204=>x"3300",
---- 205=>x"3400", 206=>x"3700", 207=>x"3400", 208=>x"3b00",
---- 209=>x"3400", 210=>x"3200", 211=>x"3300", 212=>x"3500",
---- 213=>x"3000", 214=>x"3100", 215=>x"3700", 216=>x"3000",
---- 217=>x"2a00", 218=>x"3000", 219=>x"4600", 220=>x"2800",
---- 221=>x"2600", 222=>x"3600", 223=>x"5b00", 224=>x"2700",
---- 225=>x"2c00", 226=>x"4f00", 227=>x"7a00", 228=>x"3300",
---- 229=>x"4a00", 230=>x"7100", 231=>x"8c00", 232=>x"c000",
---- 233=>x"6a00", 234=>x"8700", 235=>x"9500", 236=>x"5700",
---- 237=>x"8000", 238=>x"9500", 239=>x"9700", 240=>x"7600",
---- 241=>x"9100", 242=>x"9900", 243=>x"9600", 244=>x"8b00",
---- 245=>x"9600", 246=>x"9800", 247=>x"9100", 248=>x"9500",
---- 249=>x"9a00", 250=>x"9300", 251=>x"7100", 252=>x"9c00",
---- 253=>x"9600", 254=>x"9100", 255=>x"8e00", 256=>x"9a00",
---- 257=>x"9400", 258=>x"8f00", 259=>x"9100", 260=>x"9400",
---- 261=>x"9100", 262=>x"8e00", 263=>x"9900", 264=>x"9200",
---- 265=>x"8f00", 266=>x"9300", 267=>x"9d00", 268=>x"8e00",
---- 269=>x"9200", 270=>x"9a00", 271=>x"a000", 272=>x"9000",
---- 273=>x"9600", 274=>x"9f00", 275=>x"a300", 276=>x"9300",
---- 277=>x"9c00", 278=>x"9f00", 279=>x"a200", 280=>x"9600",
---- 281=>x"9e00", 282=>x"a100", 283=>x"a100", 284=>x"9d00",
---- 285=>x"a000", 286=>x"a000", 287=>x"a000", 288=>x"9f00",
---- 289=>x"a200", 290=>x"a000", 291=>x"9f00", 292=>x"9f00",
---- 293=>x"a100", 294=>x"a100", 295=>x"a000", 296=>x"a100",
---- 297=>x"a200", 298=>x"a200", 299=>x"a000", 300=>x"a100",
---- 301=>x"a000", 302=>x"9f00", 303=>x"a100", 304=>x"a100",
---- 305=>x"a200", 306=>x"a000", 307=>x"a100", 308=>x"a300",
---- 309=>x"a200", 310=>x"a100", 311=>x"9f00", 312=>x"a300",
---- 313=>x"a000", 314=>x"a000", 315=>x"a000", 316=>x"a100",
---- 317=>x"9c00", 318=>x"9e00", 319=>x"a100", 320=>x"a000",
---- 321=>x"9e00", 322=>x"a000", 323=>x"9f00", 324=>x"a300",
---- 325=>x"9e00", 326=>x"9e00", 327=>x"9e00", 328=>x"9e00",
---- 329=>x"6300", 330=>x"6400", 331=>x"9b00", 332=>x"9c00",
---- 333=>x"9b00", 334=>x"9e00", 335=>x"9d00", 336=>x"9d00",
---- 337=>x"9c00", 338=>x"9c00", 339=>x"9d00", 340=>x"9b00",
---- 341=>x"9c00", 342=>x"9c00", 343=>x"9b00", 344=>x"9c00",
---- 345=>x"9b00", 346=>x"9c00", 347=>x"9c00", 348=>x"9e00",
---- 349=>x"9d00", 350=>x"9e00", 351=>x"9c00", 352=>x"9c00",
---- 353=>x"9b00", 354=>x"9d00", 355=>x"9e00", 356=>x"9d00",
---- 357=>x"9a00", 358=>x"9b00", 359=>x"9c00", 360=>x"a000",
---- 361=>x"9e00", 362=>x"9d00", 363=>x"9c00", 364=>x"9d00",
---- 365=>x"9f00", 366=>x"9e00", 367=>x"9d00", 368=>x"9e00",
---- 369=>x"9e00", 370=>x"6100", 371=>x"9b00", 372=>x"9e00",
---- 373=>x"9e00", 374=>x"9d00", 375=>x"9d00", 376=>x"9f00",
---- 377=>x"9f00", 378=>x"9d00", 379=>x"9e00", 380=>x"a000",
---- 381=>x"a000", 382=>x"9e00", 383=>x"9e00", 384=>x"9f00",
---- 385=>x"9f00", 386=>x"9c00", 387=>x"9f00", 388=>x"9f00",
---- 389=>x"9f00", 390=>x"9e00", 391=>x"a000", 392=>x"9d00",
---- 393=>x"6100", 394=>x"9d00", 395=>x"9f00", 396=>x"9f00",
---- 397=>x"9f00", 398=>x"a000", 399=>x"6000", 400=>x"a000",
---- 401=>x"a100", 402=>x"9c00", 403=>x"9e00", 404=>x"a100",
---- 405=>x"a100", 406=>x"9d00", 407=>x"9f00", 408=>x"a100",
---- 409=>x"a000", 410=>x"a100", 411=>x"a100", 412=>x"a200",
---- 413=>x"9f00", 414=>x"a100", 415=>x"a000", 416=>x"a200",
---- 417=>x"9f00", 418=>x"9f00", 419=>x"9f00", 420=>x"a100",
---- 421=>x"a200", 422=>x"a200", 423=>x"9f00", 424=>x"a300",
---- 425=>x"a200", 426=>x"a100", 427=>x"a100", 428=>x"a200",
---- 429=>x"a300", 430=>x"9e00", 431=>x"a000", 432=>x"a200",
---- 433=>x"a200", 434=>x"a100", 435=>x"a200", 436=>x"a200",
---- 437=>x"a300", 438=>x"a200", 439=>x"a200", 440=>x"a400",
---- 441=>x"a400", 442=>x"a100", 443=>x"a100", 444=>x"a100",
---- 445=>x"a400", 446=>x"a400", 447=>x"a100", 448=>x"a300",
---- 449=>x"a300", 450=>x"a500", 451=>x"a100", 452=>x"a000",
---- 453=>x"a000", 454=>x"a100", 455=>x"a200", 456=>x"9f00",
---- 457=>x"a200", 458=>x"a400", 459=>x"a000", 460=>x"9a00",
---- 461=>x"9e00", 462=>x"a100", 463=>x"a100", 464=>x"9000",
---- 465=>x"6900", 466=>x"9a00", 467=>x"9b00", 468=>x"9100",
---- 469=>x"9100", 470=>x"9300", 471=>x"9000", 472=>x"9300",
---- 473=>x"9500", 474=>x"9200", 475=>x"9100", 476=>x"9200",
---- 477=>x"9600", 478=>x"9200", 479=>x"9100", 480=>x"9500",
---- 481=>x"9400", 482=>x"9200", 483=>x"9000", 484=>x"9500",
---- 485=>x"9300", 486=>x"9400", 487=>x"9000", 488=>x"9900",
---- 489=>x"9700", 490=>x"9600", 491=>x"9300", 492=>x"9c00",
---- 493=>x"9a00", 494=>x"9900", 495=>x"9800", 496=>x"9b00",
---- 497=>x"9a00", 498=>x"9a00", 499=>x"9b00", 500=>x"9c00",
---- 501=>x"9a00", 502=>x"9a00", 503=>x"9a00", 504=>x"9b00",
---- 505=>x"9a00", 506=>x"9c00", 507=>x"9d00", 508=>x"9900",
---- 509=>x"9b00", 510=>x"9900", 511=>x"9a00", 512=>x"9a00",
---- 513=>x"9a00", 514=>x"9900", 515=>x"9a00", 516=>x"9c00",
---- 517=>x"9a00", 518=>x"9800", 519=>x"9900", 520=>x"9900",
---- 521=>x"9800", 522=>x"9800", 523=>x"9800", 524=>x"9900",
---- 525=>x"6700", 526=>x"9800", 527=>x"9500", 528=>x"9a00",
---- 529=>x"9800", 530=>x"9800", 531=>x"9500", 532=>x"9700",
---- 533=>x"9500", 534=>x"9200", 535=>x"9200", 536=>x"9400",
---- 537=>x"9700", 538=>x"9400", 539=>x"9000", 540=>x"9200",
---- 541=>x"9500", 542=>x"9100", 543=>x"9500", 544=>x"9500",
---- 545=>x"9300", 546=>x"9000", 547=>x"8f00", 548=>x"9100",
---- 549=>x"9200", 550=>x"8f00", 551=>x"8e00", 552=>x"8b00",
---- 553=>x"8f00", 554=>x"8e00", 555=>x"8b00", 556=>x"8b00",
---- 557=>x"8b00", 558=>x"8800", 559=>x"8700", 560=>x"8d00",
---- 561=>x"8a00", 562=>x"8600", 563=>x"8800", 564=>x"8c00",
---- 565=>x"8900", 566=>x"8900", 567=>x"8500", 568=>x"8900",
---- 569=>x"8500", 570=>x"8300", 571=>x"8100", 572=>x"8600",
---- 573=>x"8300", 574=>x"8100", 575=>x"9000", 576=>x"8500",
---- 577=>x"8200", 578=>x"9000", 579=>x"a500", 580=>x"8300",
---- 581=>x"8e00", 582=>x"a400", 583=>x"b400", 584=>x"8b00",
---- 585=>x"a200", 586=>x"4c00", 587=>x"bd00", 588=>x"9a00",
---- 589=>x"b000", 590=>x"ba00", 591=>x"c000", 592=>x"ab00",
---- 593=>x"b800", 594=>x"c000", 595=>x"c300", 596=>x"b700",
---- 597=>x"bf00", 598=>x"c400", 599=>x"c400", 600=>x"bc00",
---- 601=>x"c200", 602=>x"c400", 603=>x"c400", 604=>x"c100",
---- 605=>x"c400", 606=>x"c400", 607=>x"c100", 608=>x"c300",
---- 609=>x"c200", 610=>x"c300", 611=>x"c000", 612=>x"c500",
---- 613=>x"c300", 614=>x"c300", 615=>x"c000", 616=>x"c400",
---- 617=>x"3c00", 618=>x"c000", 619=>x"c000", 620=>x"c300",
---- 621=>x"c200", 622=>x"c100", 623=>x"c200", 624=>x"c200",
---- 625=>x"c200", 626=>x"c100", 627=>x"c300", 628=>x"c300",
---- 629=>x"c100", 630=>x"c200", 631=>x"c200", 632=>x"c200",
---- 633=>x"c300", 634=>x"c200", 635=>x"c400", 636=>x"c200",
---- 637=>x"c200", 638=>x"c000", 639=>x"c500", 640=>x"c200",
---- 641=>x"c200", 642=>x"c500", 643=>x"ca00", 644=>x"c200",
---- 645=>x"c500", 646=>x"c800", 647=>x"cc00", 648=>x"c500",
---- 649=>x"c700", 650=>x"cb00", 651=>x"ce00", 652=>x"c700",
---- 653=>x"c900", 654=>x"ce00", 655=>x"cf00", 656=>x"ca00",
---- 657=>x"cc00", 658=>x"d000", 659=>x"d100", 660=>x"cc00",
---- 661=>x"cc00", 662=>x"cf00", 663=>x"d000", 664=>x"cd00",
---- 665=>x"d000", 666=>x"d100", 667=>x"d000", 668=>x"cf00",
---- 669=>x"d100", 670=>x"d100", 671=>x"d000", 672=>x"d100",
---- 673=>x"d200", 674=>x"d100", 675=>x"cf00", 676=>x"d100",
---- 677=>x"d100", 678=>x"d100", 679=>x"ce00", 680=>x"d100",
---- 681=>x"d100", 682=>x"d000", 683=>x"cf00", 684=>x"d100",
---- 685=>x"d000", 686=>x"d000", 687=>x"cf00", 688=>x"d100",
---- 689=>x"cf00", 690=>x"cf00", 691=>x"d000", 692=>x"d100",
---- 693=>x"d100", 694=>x"d000", 695=>x"d100", 696=>x"d100",
---- 697=>x"d100", 698=>x"d300", 699=>x"d100", 700=>x"d200",
---- 701=>x"d300", 702=>x"d100", 703=>x"d100", 704=>x"d300",
---- 705=>x"d100", 706=>x"d100", 707=>x"d100", 708=>x"d300",
---- 709=>x"d200", 710=>x"d300", 711=>x"d100", 712=>x"d200",
---- 713=>x"d300", 714=>x"2c00", 715=>x"d100", 716=>x"d300",
---- 717=>x"d300", 718=>x"d300", 719=>x"d500", 720=>x"d200",
---- 721=>x"d500", 722=>x"d600", 723=>x"d600", 724=>x"d600",
---- 725=>x"d400", 726=>x"d600", 727=>x"d800", 728=>x"d400",
---- 729=>x"d600", 730=>x"d700", 731=>x"d900", 732=>x"d600",
---- 733=>x"d700", 734=>x"d800", 735=>x"d900", 736=>x"d800",
---- 737=>x"d700", 738=>x"d700", 739=>x"d900", 740=>x"d800",
---- 741=>x"d600", 742=>x"d600", 743=>x"d700", 744=>x"d600",
---- 745=>x"d500", 746=>x"d500", 747=>x"d400", 748=>x"d400",
---- 749=>x"d400", 750=>x"2c00", 751=>x"d500", 752=>x"d500",
---- 753=>x"d400", 754=>x"d500", 755=>x"d800", 756=>x"d500",
---- 757=>x"d600", 758=>x"d600", 759=>x"d700", 760=>x"d600",
---- 761=>x"d700", 762=>x"d600", 763=>x"d800", 764=>x"d400",
---- 765=>x"d600", 766=>x"d600", 767=>x"d600", 768=>x"d500",
---- 769=>x"d500", 770=>x"d500", 771=>x"d300", 772=>x"d300",
---- 773=>x"d400", 774=>x"d200", 775=>x"d200", 776=>x"d200",
---- 777=>x"d200", 778=>x"d100", 779=>x"d000", 780=>x"d000",
---- 781=>x"d000", 782=>x"cf00", 783=>x"ce00", 784=>x"d100",
---- 785=>x"d100", 786=>x"cd00", 787=>x"cc00", 788=>x"d100",
---- 789=>x"d100", 790=>x"cb00", 791=>x"c700", 792=>x"d000",
---- 793=>x"d200", 794=>x"cc00", 795=>x"c200", 796=>x"d000",
---- 797=>x"d100", 798=>x"cb00", 799=>x"bf00", 800=>x"ce00",
---- 801=>x"ca00", 802=>x"c400", 803=>x"b600", 804=>x"c800",
---- 805=>x"bd00", 806=>x"b300", 807=>x"9a00", 808=>x"c100",
---- 809=>x"a800", 810=>x"8a00", 811=>x"5b00", 812=>x"b900",
---- 813=>x"8b00", 814=>x"5400", 815=>x"3300", 816=>x"a900",
---- 817=>x"7300", 818=>x"3700", 819=>x"2a00", 820=>x"9800",
---- 821=>x"5a00", 822=>x"2c00", 823=>x"2b00", 824=>x"8500",
---- 825=>x"4900", 826=>x"3000", 827=>x"3a00", 828=>x"7000",
---- 829=>x"4200", 830=>x"3a00", 831=>x"4e00", 832=>x"5a00",
---- 833=>x"4200", 834=>x"4800", 835=>x"5900", 836=>x"4c00",
---- 837=>x"4700", 838=>x"5200", 839=>x"6100", 840=>x"4b00",
---- 841=>x"5200", 842=>x"5700", 843=>x"5f00", 844=>x"4f00",
---- 845=>x"5700", 846=>x"5d00", 847=>x"5a00", 848=>x"5800",
---- 849=>x"a200", 850=>x"5e00", 851=>x"5800", 852=>x"5b00",
---- 853=>x"6200", 854=>x"5e00", 855=>x"5b00", 856=>x"5d00",
---- 857=>x"5f00", 858=>x"5b00", 859=>x"6200", 860=>x"5c00",
---- 861=>x"5b00", 862=>x"5e00", 863=>x"6800", 864=>x"5c00",
---- 865=>x"5b00", 866=>x"6300", 867=>x"6600", 868=>x"5a00",
---- 869=>x"5d00", 870=>x"6200", 871=>x"6800", 872=>x"5700",
---- 873=>x"5e00", 874=>x"6100", 875=>x"6b00", 876=>x"5e00",
---- 877=>x"5e00", 878=>x"6400", 879=>x"6e00", 880=>x"6200",
---- 881=>x"6100", 882=>x"6500", 883=>x"7100", 884=>x"6200",
---- 885=>x"6500", 886=>x"6500", 887=>x"6c00", 888=>x"6100",
---- 889=>x"9b00", 890=>x"6a00", 891=>x"6d00", 892=>x"6000",
---- 893=>x"6700", 894=>x"6a00", 895=>x"6c00", 896=>x"5c00",
---- 897=>x"6500", 898=>x"6600", 899=>x"6800", 900=>x"5d00",
---- 901=>x"6100", 902=>x"6700", 903=>x"6200", 904=>x"5c00",
---- 905=>x"6600", 906=>x"6600", 907=>x"5b00", 908=>x"6300",
---- 909=>x"6400", 910=>x"6000", 911=>x"5600", 912=>x"6300",
---- 913=>x"6000", 914=>x"5700", 915=>x"4a00", 916=>x"6300",
---- 917=>x"5800", 918=>x"5000", 919=>x"4d00", 920=>x"5d00",
---- 921=>x"4d00", 922=>x"4a00", 923=>x"5100", 924=>x"5200",
---- 925=>x"4700", 926=>x"4900", 927=>x"5200", 928=>x"4800",
---- 929=>x"4700", 930=>x"5400", 931=>x"5f00", 932=>x"4700",
---- 933=>x"4f00", 934=>x"6000", 935=>x"6600", 936=>x"4e00",
---- 937=>x"5a00", 938=>x"6800", 939=>x"6a00", 940=>x"5a00",
---- 941=>x"6700", 942=>x"6d00", 943=>x"6600", 944=>x"6300",
---- 945=>x"6b00", 946=>x"6c00", 947=>x"6200", 948=>x"6700",
---- 949=>x"6b00", 950=>x"6500", 951=>x"5d00", 952=>x"7300",
---- 953=>x"6900", 954=>x"5700", 955=>x"5500", 956=>x"6900",
---- 957=>x"5d00", 958=>x"5500", 959=>x"5000", 960=>x"6100",
---- 961=>x"5200", 962=>x"4b00", 963=>x"4d00", 964=>x"5b00",
---- 965=>x"5100", 966=>x"4900", 967=>x"4d00", 968=>x"5000",
---- 969=>x"4e00", 970=>x"4b00", 971=>x"4c00", 972=>x"4900",
---- 973=>x"4700", 974=>x"4700", 975=>x"4d00", 976=>x"4500",
---- 977=>x"4200", 978=>x"4100", 979=>x"4c00", 980=>x"4700",
---- 981=>x"3f00", 982=>x"4200", 983=>x"4f00", 984=>x"4000",
---- 985=>x"3f00", 986=>x"4800", 987=>x"5c00", 988=>x"3c00",
---- 989=>x"4200", 990=>x"5400", 991=>x"6700", 992=>x"4000",
---- 993=>x"4b00", 994=>x"5f00", 995=>x"6c00", 996=>x"4800",
---- 997=>x"5400", 998=>x"6300", 999=>x"7200", 1000=>x"5000",
---- 1001=>x"6100", 1002=>x"6f00", 1003=>x"7400", 1004=>x"5f00",
---- 1005=>x"6b00", 1006=>x"7600", 1007=>x"7b00", 1008=>x"6b00",
---- 1009=>x"7700", 1010=>x"7c00", 1011=>x"7d00", 1012=>x"7500",
---- 1013=>x"8000", 1014=>x"7e00", 1015=>x"7e00", 1016=>x"7d00",
---- 1017=>x"8100", 1018=>x"7f00", 1019=>x"7e00", 1020=>x"7f00",
---- 1021=>x"8000", 1022=>x"7f00", 1023=>x"7b00"),
----
---- 60 => (0=>x"7c00", 1=>x"7d00", 2=>x"7f00", 3=>x"7e00", 4=>x"7c00",
---- 5=>x"7d00", 6=>x"7f00", 7=>x"7e00", 8=>x"7c00",
---- 9=>x"7d00", 10=>x"7f00", 11=>x"7e00", 12=>x"7a00",
---- 13=>x"7b00", 14=>x"7e00", 15=>x"7d00", 16=>x"7a00",
---- 17=>x"7d00", 18=>x"7f00", 19=>x"7e00", 20=>x"7b00",
---- 21=>x"7d00", 22=>x"7d00", 23=>x"7e00", 24=>x"7e00",
---- 25=>x"7e00", 26=>x"7b00", 27=>x"7b00", 28=>x"7d00",
---- 29=>x"7d00", 30=>x"7d00", 31=>x"8000", 32=>x"8000",
---- 33=>x"8000", 34=>x"8000", 35=>x"8300", 36=>x"8100",
---- 37=>x"8300", 38=>x"8300", 39=>x"8500", 40=>x"8400",
---- 41=>x"8600", 42=>x"8800", 43=>x"8b00", 44=>x"8400",
---- 45=>x"8600", 46=>x"8a00", 47=>x"8800", 48=>x"8800",
---- 49=>x"8700", 50=>x"8700", 51=>x"7100", 52=>x"8800",
---- 53=>x"8700", 54=>x"8f00", 55=>x"4a00", 56=>x"8600",
---- 57=>x"6c00", 58=>x"4800", 59=>x"2b00", 60=>x"7000",
---- 61=>x"4600", 62=>x"2a00", 63=>x"2c00", 64=>x"5000",
---- 65=>x"3000", 66=>x"2c00", 67=>x"2800", 68=>x"3000",
---- 69=>x"2800", 70=>x"d400", 71=>x"2b00", 72=>x"2a00",
---- 73=>x"2900", 74=>x"2b00", 75=>x"2d00", 76=>x"2d00",
---- 77=>x"2b00", 78=>x"2a00", 79=>x"2e00", 80=>x"2b00",
---- 81=>x"2e00", 82=>x"d300", 83=>x"2d00", 84=>x"2c00",
---- 85=>x"2d00", 86=>x"3200", 87=>x"3500", 88=>x"3000",
---- 89=>x"3100", 90=>x"3400", 91=>x"3500", 92=>x"cf00",
---- 93=>x"3000", 94=>x"3500", 95=>x"3700", 96=>x"3300",
---- 97=>x"3800", 98=>x"3600", 99=>x"3800", 100=>x"3400",
---- 101=>x"3600", 102=>x"3500", 103=>x"3700", 104=>x"3500",
---- 105=>x"3600", 106=>x"3300", 107=>x"3200", 108=>x"3700",
---- 109=>x"3700", 110=>x"3500", 111=>x"3100", 112=>x"3700",
---- 113=>x"3600", 114=>x"3300", 115=>x"3300", 116=>x"3800",
---- 117=>x"3300", 118=>x"3600", 119=>x"3600", 120=>x"3400",
---- 121=>x"3700", 122=>x"3300", 123=>x"2e00", 124=>x"3600",
---- 125=>x"3500", 126=>x"2d00", 127=>x"2d00", 128=>x"3400",
---- 129=>x"2f00", 130=>x"2c00", 131=>x"2c00", 132=>x"3400",
---- 133=>x"2c00", 134=>x"2a00", 135=>x"2d00", 136=>x"3000",
---- 137=>x"2d00", 138=>x"2c00", 139=>x"3300", 140=>x"2e00",
---- 141=>x"3400", 142=>x"3500", 143=>x"3600", 144=>x"2f00",
---- 145=>x"3a00", 146=>x"3800", 147=>x"3100", 148=>x"3300",
---- 149=>x"3900", 150=>x"3800", 151=>x"3400", 152=>x"3700",
---- 153=>x"3900", 154=>x"3300", 155=>x"3000", 156=>x"3700",
---- 157=>x"3600", 158=>x"3000", 159=>x"2f00", 160=>x"3100",
---- 161=>x"2d00", 162=>x"3200", 163=>x"2d00", 164=>x"2e00",
---- 165=>x"3000", 166=>x"3000", 167=>x"2d00", 168=>x"2c00",
---- 169=>x"2f00", 170=>x"cf00", 171=>x"3100", 172=>x"2f00",
---- 173=>x"2f00", 174=>x"3f00", 175=>x"4400", 176=>x"2e00",
---- 177=>x"3600", 178=>x"3f00", 179=>x"4200", 180=>x"3000",
---- 181=>x"3c00", 182=>x"3a00", 183=>x"4000", 184=>x"3000",
---- 185=>x"3700", 186=>x"4000", 187=>x"4500", 188=>x"3300",
---- 189=>x"3600", 190=>x"3e00", 191=>x"4a00", 192=>x"3e00",
---- 193=>x"3f00", 194=>x"3900", 195=>x"4600", 196=>x"3b00",
---- 197=>x"3e00", 198=>x"3d00", 199=>x"4900", 200=>x"3a00",
---- 201=>x"3e00", 202=>x"4600", 203=>x"5c00", 204=>x"3500",
---- 205=>x"3e00", 206=>x"5b00", 207=>x"7b00", 208=>x"c500",
---- 209=>x"5600", 210=>x"7800", 211=>x"8c00", 212=>x"4600",
---- 213=>x"6e00", 214=>x"7400", 215=>x"9700", 216=>x"6800",
---- 217=>x"8700", 218=>x"9500", 219=>x"9800", 220=>x"8300",
---- 221=>x"9500", 222=>x"9800", 223=>x"9200", 224=>x"9200",
---- 225=>x"9800", 226=>x"9100", 227=>x"8c00", 228=>x"9700",
---- 229=>x"9500", 230=>x"9000", 231=>x"8900", 232=>x"9600",
---- 233=>x"8f00", 234=>x"8e00", 235=>x"8900", 236=>x"9300",
---- 237=>x"8f00", 238=>x"8b00", 239=>x"8f00", 240=>x"9000",
---- 241=>x"8b00", 242=>x"8e00", 243=>x"9900", 244=>x"8b00",
---- 245=>x"8c00", 246=>x"9800", 247=>x"9e00", 248=>x"8d00",
---- 249=>x"9400", 250=>x"9e00", 251=>x"9f00", 252=>x"9100",
---- 253=>x"9a00", 254=>x"9f00", 255=>x"5f00", 256=>x"9900",
---- 257=>x"9f00", 258=>x"a000", 259=>x"a000", 260=>x"9f00",
---- 261=>x"a100", 262=>x"a300", 263=>x"9f00", 264=>x"a000",
---- 265=>x"a200", 266=>x"a300", 267=>x"9f00", 268=>x"a100",
---- 269=>x"a000", 270=>x"9f00", 271=>x"9e00", 272=>x"9f00",
---- 273=>x"a000", 274=>x"a000", 275=>x"9c00", 276=>x"a100",
---- 277=>x"9f00", 278=>x"a000", 279=>x"9d00", 280=>x"a100",
---- 281=>x"a000", 282=>x"9d00", 283=>x"9e00", 284=>x"a100",
---- 285=>x"9f00", 286=>x"a100", 287=>x"9e00", 288=>x"9f00",
---- 289=>x"9e00", 290=>x"9f00", 291=>x"9c00", 292=>x"a000",
---- 293=>x"9f00", 294=>x"9f00", 295=>x"9d00", 296=>x"9f00",
---- 297=>x"9f00", 298=>x"9d00", 299=>x"a000", 300=>x"9e00",
---- 301=>x"a000", 302=>x"a000", 303=>x"9d00", 304=>x"a000",
---- 305=>x"a000", 306=>x"a100", 307=>x"9f00", 308=>x"a000",
---- 309=>x"a100", 310=>x"a000", 311=>x"9f00", 312=>x"9e00",
---- 313=>x"a200", 314=>x"a000", 315=>x"9b00", 316=>x"9f00",
---- 317=>x"9f00", 318=>x"9f00", 319=>x"9e00", 320=>x"9f00",
---- 321=>x"9e00", 322=>x"9d00", 323=>x"9f00", 324=>x"9f00",
---- 325=>x"9d00", 326=>x"9f00", 327=>x"9e00", 328=>x"9d00",
---- 329=>x"9d00", 330=>x"9d00", 331=>x"9f00", 332=>x"9d00",
---- 333=>x"5f00", 334=>x"9f00", 335=>x"9d00", 336=>x"9b00",
---- 337=>x"9e00", 338=>x"a000", 339=>x"9e00", 340=>x"9c00",
---- 341=>x"9d00", 342=>x"9c00", 343=>x"9c00", 344=>x"9b00",
---- 345=>x"9e00", 346=>x"9c00", 347=>x"9b00", 348=>x"9c00",
---- 349=>x"9d00", 350=>x"9d00", 351=>x"9b00", 352=>x"9c00",
---- 353=>x"9b00", 354=>x"9b00", 355=>x"9b00", 356=>x"9d00",
---- 357=>x"9b00", 358=>x"9b00", 359=>x"9c00", 360=>x"9e00",
---- 361=>x"9a00", 362=>x"9800", 363=>x"9a00", 364=>x"9d00",
---- 365=>x"9a00", 366=>x"6600", 367=>x"9900", 368=>x"9b00",
---- 369=>x"9b00", 370=>x"9c00", 371=>x"9b00", 372=>x"9c00",
---- 373=>x"9d00", 374=>x"9c00", 375=>x"9c00", 376=>x"9e00",
---- 377=>x"9f00", 378=>x"9b00", 379=>x"9d00", 380=>x"9f00",
---- 381=>x"9e00", 382=>x"9c00", 383=>x"9c00", 384=>x"9f00",
---- 385=>x"9c00", 386=>x"9a00", 387=>x"9b00", 388=>x"9d00",
---- 389=>x"9d00", 390=>x"9b00", 391=>x"9a00", 392=>x"9e00",
---- 393=>x"9e00", 394=>x"9e00", 395=>x"9c00", 396=>x"a000",
---- 397=>x"9c00", 398=>x"9b00", 399=>x"9c00", 400=>x"9e00",
---- 401=>x"9c00", 402=>x"9c00", 403=>x"9e00", 404=>x"9e00",
---- 405=>x"9d00", 406=>x"9e00", 407=>x"9d00", 408=>x"9f00",
---- 409=>x"9f00", 410=>x"a000", 411=>x"9e00", 412=>x"9e00",
---- 413=>x"9e00", 414=>x"9f00", 415=>x"9f00", 416=>x"9d00",
---- 417=>x"9f00", 418=>x"a000", 419=>x"a000", 420=>x"a100",
---- 421=>x"5f00", 422=>x"a100", 423=>x"6000", 424=>x"a300",
---- 425=>x"a300", 426=>x"a200", 427=>x"9f00", 428=>x"a100",
---- 429=>x"a100", 430=>x"a200", 431=>x"9f00", 432=>x"a200",
---- 433=>x"a100", 434=>x"9f00", 435=>x"a000", 436=>x"a000",
---- 437=>x"a000", 438=>x"a100", 439=>x"a000", 440=>x"a100",
---- 441=>x"9e00", 442=>x"a000", 443=>x"9e00", 444=>x"a000",
---- 445=>x"9e00", 446=>x"9f00", 447=>x"9e00", 448=>x"9f00",
---- 449=>x"9f00", 450=>x"a100", 451=>x"a100", 452=>x"a200",
---- 453=>x"9f00", 454=>x"9f00", 455=>x"9e00", 456=>x"a100",
---- 457=>x"a100", 458=>x"a100", 459=>x"9d00", 460=>x"a000",
---- 461=>x"9f00", 462=>x"9e00", 463=>x"9c00", 464=>x"9b00",
---- 465=>x"6300", 466=>x"9d00", 467=>x"9d00", 468=>x"9200",
---- 469=>x"9600", 470=>x"6700", 471=>x"9900", 472=>x"9100",
---- 473=>x"8f00", 474=>x"9200", 475=>x"8e00", 476=>x"9000",
---- 477=>x"9000", 478=>x"9000", 479=>x"8e00", 480=>x"9100",
---- 481=>x"8e00", 482=>x"8f00", 483=>x"8e00", 484=>x"9000",
---- 485=>x"8f00", 486=>x"9000", 487=>x"9000", 488=>x"9300",
---- 489=>x"9200", 490=>x"9300", 491=>x"9200", 492=>x"9500",
---- 493=>x"9500", 494=>x"9600", 495=>x"9400", 496=>x"9800",
---- 497=>x"9b00", 498=>x"9900", 499=>x"9800", 500=>x"9b00",
---- 501=>x"9c00", 502=>x"9c00", 503=>x"9d00", 504=>x"9900",
---- 505=>x"9b00", 506=>x"9c00", 507=>x"9b00", 508=>x"9a00",
---- 509=>x"9d00", 510=>x"9d00", 511=>x"9c00", 512=>x"9c00",
---- 513=>x"9b00", 514=>x"6200", 515=>x"9c00", 516=>x"9a00",
---- 517=>x"9a00", 518=>x"9b00", 519=>x"9a00", 520=>x"9900",
---- 521=>x"9900", 522=>x"9800", 523=>x"9900", 524=>x"6800",
---- 525=>x"9700", 526=>x"9800", 527=>x"9700", 528=>x"9500",
---- 529=>x"9700", 530=>x"9800", 531=>x"9200", 532=>x"9500",
---- 533=>x"9300", 534=>x"9300", 535=>x"8f00", 536=>x"9200",
---- 537=>x"9100", 538=>x"8f00", 539=>x"9000", 540=>x"9100",
---- 541=>x"9100", 542=>x"8e00", 543=>x"8a00", 544=>x"8d00",
---- 545=>x"8d00", 546=>x"8e00", 547=>x"8b00", 548=>x"8900",
---- 549=>x"8a00", 550=>x"8d00", 551=>x"8a00", 552=>x"8800",
---- 553=>x"8800", 554=>x"8a00", 555=>x"7700", 556=>x"8800",
---- 557=>x"8600", 558=>x"8700", 559=>x"8800", 560=>x"8800",
---- 561=>x"8300", 562=>x"8900", 563=>x"9700", 564=>x"8400",
---- 565=>x"8a00", 566=>x"9d00", 567=>x"a900", 568=>x"8e00",
---- 569=>x"a600", 570=>x"b200", 571=>x"bd00", 572=>x"a700",
---- 573=>x"b200", 574=>x"bc00", 575=>x"c300", 576=>x"b500",
---- 577=>x"bd00", 578=>x"c200", 579=>x"c400", 580=>x"bd00",
---- 581=>x"c300", 582=>x"c600", 583=>x"c500", 584=>x"c100",
---- 585=>x"c600", 586=>x"c600", 587=>x"c400", 588=>x"c300",
---- 589=>x"c400", 590=>x"c400", 591=>x"c300", 592=>x"c200",
---- 593=>x"c200", 594=>x"c200", 595=>x"c300", 596=>x"c200",
---- 597=>x"c100", 598=>x"c100", 599=>x"c100", 600=>x"c200",
---- 601=>x"c200", 602=>x"c200", 603=>x"c300", 604=>x"c300",
---- 605=>x"c100", 606=>x"c000", 607=>x"c200", 608=>x"c100",
---- 609=>x"c000", 610=>x"c100", 611=>x"c200", 612=>x"c000",
---- 613=>x"c100", 614=>x"c100", 615=>x"c100", 616=>x"c000",
---- 617=>x"c100", 618=>x"c200", 619=>x"c500", 620=>x"c100",
---- 621=>x"c200", 622=>x"c300", 623=>x"ca00", 624=>x"c100",
---- 625=>x"c400", 626=>x"c800", 627=>x"cc00", 628=>x"c300",
---- 629=>x"c900", 630=>x"cd00", 631=>x"d100", 632=>x"c700",
---- 633=>x"cb00", 634=>x"ce00", 635=>x"d100", 636=>x"c800",
---- 637=>x"cd00", 638=>x"d000", 639=>x"cf00", 640=>x"ca00",
---- 641=>x"cd00", 642=>x"ce00", 643=>x"cd00", 644=>x"cd00",
---- 645=>x"ce00", 646=>x"cd00", 647=>x"cd00", 648=>x"cd00",
---- 649=>x"ce00", 650=>x"cc00", 651=>x"cc00", 652=>x"cf00",
---- 653=>x"d000", 654=>x"d000", 655=>x"cf00", 656=>x"cf00",
---- 657=>x"cf00", 658=>x"2f00", 659=>x"cf00", 660=>x"ce00",
---- 661=>x"ce00", 662=>x"d000", 663=>x"cc00", 664=>x"cf00",
---- 665=>x"d000", 666=>x"ce00", 667=>x"ce00", 668=>x"cf00",
---- 669=>x"ce00", 670=>x"cd00", 671=>x"ce00", 672=>x"ce00",
---- 673=>x"ce00", 674=>x"cd00", 675=>x"ce00", 676=>x"cf00",
---- 677=>x"d000", 678=>x"d000", 679=>x"ce00", 680=>x"cf00",
---- 681=>x"d300", 682=>x"d000", 683=>x"d000", 684=>x"d100",
---- 685=>x"d200", 686=>x"d000", 687=>x"cf00", 688=>x"d100",
---- 689=>x"d100", 690=>x"d200", 691=>x"d000", 692=>x"d100",
---- 693=>x"d200", 694=>x"d200", 695=>x"d000", 696=>x"ce00",
---- 697=>x"d100", 698=>x"d200", 699=>x"d000", 700=>x"cf00",
---- 701=>x"d100", 702=>x"d100", 703=>x"2e00", 704=>x"d000",
---- 705=>x"d300", 706=>x"d300", 707=>x"d100", 708=>x"d300",
---- 709=>x"d400", 710=>x"d300", 711=>x"d400", 712=>x"d300",
---- 713=>x"d500", 714=>x"2b00", 715=>x"d500", 716=>x"d400",
---- 717=>x"d500", 718=>x"d400", 719=>x"d500", 720=>x"d600",
---- 721=>x"d600", 722=>x"d600", 723=>x"2800", 724=>x"d900",
---- 725=>x"d700", 726=>x"d700", 727=>x"d600", 728=>x"d900",
---- 729=>x"d800", 730=>x"d600", 731=>x"d400", 732=>x"d900",
---- 733=>x"d800", 734=>x"d500", 735=>x"2d00", 736=>x"d500",
---- 737=>x"d500", 738=>x"d300", 739=>x"d100", 740=>x"d500",
---- 741=>x"d400", 742=>x"d200", 743=>x"d200", 744=>x"d500",
---- 745=>x"d400", 746=>x"d400", 747=>x"d400", 748=>x"d600",
---- 749=>x"d600", 750=>x"d600", 751=>x"d500", 752=>x"d700",
---- 753=>x"d700", 754=>x"d700", 755=>x"d400", 756=>x"d700",
---- 757=>x"d700", 758=>x"d500", 759=>x"d300", 760=>x"d600",
---- 761=>x"d500", 762=>x"d400", 763=>x"d100", 764=>x"d500",
---- 765=>x"d400", 766=>x"d200", 767=>x"d000", 768=>x"d300",
---- 769=>x"d200", 770=>x"d000", 771=>x"cf00", 772=>x"d200",
---- 773=>x"d100", 774=>x"ce00", 775=>x"ca00", 776=>x"d200",
---- 777=>x"cd00", 778=>x"c700", 779=>x"bf00", 780=>x"cd00",
---- 781=>x"c800", 782=>x"be00", 783=>x"b200", 784=>x"c900",
---- 785=>x"3a00", 786=>x"ba00", 787=>x"ab00", 788=>x"be00",
---- 789=>x"bb00", 790=>x"b200", 791=>x"a100", 792=>x"b900",
---- 793=>x"af00", 794=>x"9600", 795=>x"7200", 796=>x"b100",
---- 797=>x"9700", 798=>x"5f00", 799=>x"3600", 800=>x"9e00",
---- 801=>x"6b00", 802=>x"3100", 803=>x"2900", 804=>x"6f00",
---- 805=>x"3f00", 806=>x"d300", 807=>x"3500", 808=>x"3200",
---- 809=>x"2a00", 810=>x"3600", 811=>x"4600", 812=>x"2800",
---- 813=>x"3100", 814=>x"4d00", 815=>x"5700", 816=>x"3500",
---- 817=>x"4b00", 818=>x"5c00", 819=>x"5b00", 820=>x"4300",
---- 821=>x"5600", 822=>x"5b00", 823=>x"5a00", 824=>x"5400",
---- 825=>x"5c00", 826=>x"5900", 827=>x"5d00", 828=>x"6100",
---- 829=>x"5f00", 830=>x"5800", 831=>x"5b00", 832=>x"6200",
---- 833=>x"5800", 834=>x"5a00", 835=>x"5c00", 836=>x"5e00",
---- 837=>x"5900", 838=>x"6100", 839=>x"5f00", 840=>x"5800",
---- 841=>x"5e00", 842=>x"6400", 843=>x"6100", 844=>x"5800",
---- 845=>x"6200", 846=>x"6800", 847=>x"6900", 848=>x"5e00",
---- 849=>x"6700", 850=>x"6800", 851=>x"6e00", 852=>x"6400",
---- 853=>x"6600", 854=>x"6a00", 855=>x"7000", 856=>x"6800",
---- 857=>x"6900", 858=>x"6e00", 859=>x"7200", 860=>x"6b00",
---- 861=>x"6f00", 862=>x"7100", 863=>x"8c00", 864=>x"9100",
---- 865=>x"7300", 866=>x"7200", 867=>x"7400", 868=>x"7000",
---- 869=>x"7200", 870=>x"7300", 871=>x"6f00", 872=>x"6f00",
---- 873=>x"7300", 874=>x"6f00", 875=>x"6400", 876=>x"7500",
---- 877=>x"7000", 878=>x"6900", 879=>x"6300", 880=>x"7400",
---- 881=>x"7000", 882=>x"6a00", 883=>x"6500", 884=>x"7000",
---- 885=>x"6f00", 886=>x"6800", 887=>x"5c00", 888=>x"6f00",
---- 889=>x"6800", 890=>x"5f00", 891=>x"5c00", 892=>x"6800",
---- 893=>x"6300", 894=>x"5a00", 895=>x"5600", 896=>x"6400",
---- 897=>x"5a00", 898=>x"5700", 899=>x"5500", 900=>x"5900",
---- 901=>x"4d00", 902=>x"5600", 903=>x"6000", 904=>x"b700",
---- 905=>x"4900", 906=>x"5900", 907=>x"6600", 908=>x"4b00",
---- 909=>x"5000", 910=>x"6000", 911=>x"6c00", 912=>x"4d00",
---- 913=>x"5900", 914=>x"6600", 915=>x"6c00", 916=>x"5300",
---- 917=>x"5d00", 918=>x"6800", 919=>x"6900", 920=>x"5e00",
---- 921=>x"6500", 922=>x"6700", 923=>x"6300", 924=>x"6400",
---- 925=>x"6a00", 926=>x"6300", 927=>x"5f00", 928=>x"6b00",
---- 929=>x"6300", 930=>x"5e00", 931=>x"5f00", 932=>x"6a00",
---- 933=>x"6000", 934=>x"5c00", 935=>x"5f00", 936=>x"5b00",
---- 937=>x"5c00", 938=>x"5d00", 939=>x"6000", 940=>x"5a00",
---- 941=>x"5900", 942=>x"5a00", 943=>x"5a00", 944=>x"5b00",
---- 945=>x"5900", 946=>x"5600", 947=>x"5500", 948=>x"5600",
---- 949=>x"5500", 950=>x"5500", 951=>x"5400", 952=>x"5200",
---- 953=>x"5400", 954=>x"5400", 955=>x"5200", 956=>x"4e00",
---- 957=>x"5100", 958=>x"5100", 959=>x"5600", 960=>x"4d00",
---- 961=>x"4c00", 962=>x"5100", 963=>x"5c00", 964=>x"4e00",
---- 965=>x"5000", 966=>x"5300", 967=>x"5f00", 968=>x"4e00",
---- 969=>x"5300", 970=>x"6100", 971=>x"6b00", 972=>x"5100",
---- 973=>x"5a00", 974=>x"6300", 975=>x"7000", 976=>x"5800",
---- 977=>x"5e00", 978=>x"6900", 979=>x"7100", 980=>x"6000",
---- 981=>x"6700", 982=>x"7000", 983=>x"7200", 984=>x"6a00",
---- 985=>x"6f00", 986=>x"7400", 987=>x"7500", 988=>x"6c00",
---- 989=>x"6d00", 990=>x"7300", 991=>x"7600", 992=>x"6f00",
---- 993=>x"7400", 994=>x"7900", 995=>x"7300", 996=>x"7300",
---- 997=>x"7900", 998=>x"7900", 999=>x"6d00", 1000=>x"7e00",
---- 1001=>x"7d00", 1002=>x"7100", 1003=>x"6b00", 1004=>x"7a00",
---- 1005=>x"7500", 1006=>x"6d00", 1007=>x"6700", 1008=>x"8400",
---- 1009=>x"6f00", 1010=>x"6b00", 1011=>x"6200", 1012=>x"7500",
---- 1013=>x"6d00", 1014=>x"6300", 1015=>x"5800", 1016=>x"7800",
---- 1017=>x"6600", 1018=>x"5600", 1019=>x"4d00", 1020=>x"7100",
---- 1021=>x"5e00", 1022=>x"4a00", 1023=>x"3d00"),
----
---- 61 => (0=>x"8300", 1=>x"7d00", 2=>x"7e00", 3=>x"7900", 4=>x"7b00",
---- 5=>x"7d00", 6=>x"7e00", 7=>x"7a00", 8=>x"7d00",
---- 9=>x"7d00", 10=>x"7d00", 11=>x"7a00", 12=>x"7c00",
---- 13=>x"7f00", 14=>x"7e00", 15=>x"7d00", 16=>x"7d00",
---- 17=>x"7e00", 18=>x"7f00", 19=>x"8100", 20=>x"7e00",
---- 21=>x"7c00", 22=>x"7f00", 23=>x"8300", 24=>x"7d00",
---- 25=>x"7d00", 26=>x"8300", 27=>x"8500", 28=>x"8100",
---- 29=>x"8000", 30=>x"8700", 31=>x"8400", 32=>x"8500",
---- 33=>x"8700", 34=>x"8300", 35=>x"7000", 36=>x"8800",
---- 37=>x"8300", 38=>x"6e00", 39=>x"4e00", 40=>x"8400",
---- 41=>x"7100", 42=>x"4d00", 43=>x"3400", 44=>x"7200",
---- 45=>x"4600", 46=>x"3400", 47=>x"2f00", 48=>x"4900",
---- 49=>x"4000", 50=>x"3600", 51=>x"2f00", 52=>x"2f00",
---- 53=>x"3700", 54=>x"3500", 55=>x"2800", 56=>x"2700",
---- 57=>x"2c00", 58=>x"2f00", 59=>x"2d00", 60=>x"2e00",
---- 61=>x"d100", 62=>x"2e00", 63=>x"2e00", 64=>x"3300",
---- 65=>x"2f00", 66=>x"3000", 67=>x"2b00", 68=>x"2f00",
---- 69=>x"c700", 70=>x"3700", 71=>x"3400", 72=>x"3000",
---- 73=>x"3200", 74=>x"3500", 75=>x"3800", 76=>x"3700",
---- 77=>x"3800", 78=>x"3800", 79=>x"3a00", 80=>x"3800",
---- 81=>x"3b00", 82=>x"3800", 83=>x"3700", 84=>x"3700",
---- 85=>x"3900", 86=>x"3700", 87=>x"3400", 88=>x"3900",
---- 89=>x"3c00", 90=>x"3900", 91=>x"3700", 92=>x"3800",
---- 93=>x"3c00", 94=>x"3800", 95=>x"3600", 96=>x"c300",
---- 97=>x"3c00", 98=>x"3a00", 99=>x"3800", 100=>x"3900",
---- 101=>x"3700", 102=>x"3700", 103=>x"3800", 104=>x"3400",
---- 105=>x"3200", 106=>x"3400", 107=>x"3200", 108=>x"3600",
---- 109=>x"3300", 110=>x"2e00", 111=>x"2c00", 112=>x"3400",
---- 113=>x"2e00", 114=>x"2b00", 115=>x"3200", 116=>x"3300",
---- 117=>x"3300", 118=>x"2f00", 119=>x"3100", 120=>x"2c00",
---- 121=>x"2e00", 122=>x"3000", 123=>x"3900", 124=>x"2b00",
---- 125=>x"2e00", 126=>x"3700", 127=>x"3400", 128=>x"2c00",
---- 129=>x"3100", 130=>x"3500", 131=>x"3400", 132=>x"3000",
---- 133=>x"3400", 134=>x"3200", 135=>x"2c00", 136=>x"3500",
---- 137=>x"3300", 138=>x"d100", 139=>x"2b00", 140=>x"3700",
---- 141=>x"3400", 142=>x"2d00", 143=>x"2f00", 144=>x"3100",
---- 145=>x"2e00", 146=>x"d300", 147=>x"3300", 148=>x"3200",
---- 149=>x"3000", 150=>x"3200", 151=>x"3600", 152=>x"2e00",
---- 153=>x"3100", 154=>x"3200", 155=>x"3700", 156=>x"3200",
---- 157=>x"3100", 158=>x"3700", 159=>x"3d00", 160=>x"2f00",
---- 161=>x"3300", 162=>x"3e00", 163=>x"4f00", 164=>x"3200",
---- 165=>x"3b00", 166=>x"4200", 167=>x"4d00", 168=>x"3600",
---- 169=>x"4400", 170=>x"4b00", 171=>x"4300", 172=>x"3e00",
---- 173=>x"4700", 174=>x"5100", 175=>x"4100", 176=>x"4400",
---- 177=>x"4800", 178=>x"4c00", 179=>x"4500", 180=>x"4900",
---- 181=>x"4a00", 182=>x"4d00", 183=>x"5800", 184=>x"4d00",
---- 185=>x"4c00", 186=>x"5800", 187=>x"6f00", 188=>x"4e00",
---- 189=>x"5b00", 190=>x"7000", 191=>x"8500", 192=>x"5900",
---- 193=>x"7100", 194=>x"8200", 195=>x"9200", 196=>x"6900",
---- 197=>x"8300", 198=>x"8e00", 199=>x"9100", 200=>x"7e00",
---- 201=>x"8d00", 202=>x"9200", 203=>x"8f00", 204=>x"8e00",
---- 205=>x"9000", 206=>x"8c00", 207=>x"8f00", 208=>x"9400",
---- 209=>x"8f00", 210=>x"8f00", 211=>x"8d00", 212=>x"9400",
---- 213=>x"8d00", 214=>x"8900", 215=>x"8700", 216=>x"9100",
---- 217=>x"8d00", 218=>x"8200", 219=>x"8b00", 220=>x"8e00",
---- 221=>x"8500", 222=>x"8900", 223=>x"9a00", 224=>x"8600",
---- 225=>x"8700", 226=>x"9400", 227=>x"9e00", 228=>x"8900",
---- 229=>x"9400", 230=>x"9c00", 231=>x"a200", 232=>x"9300",
---- 233=>x"9c00", 234=>x"a100", 235=>x"a700", 236=>x"9900",
---- 237=>x"a300", 238=>x"a300", 239=>x"a600", 240=>x"9f00",
---- 241=>x"a200", 242=>x"a200", 243=>x"a200", 244=>x"a000",
---- 245=>x"a100", 246=>x"a000", 247=>x"a100", 248=>x"9e00",
---- 249=>x"a100", 250=>x"9d00", 251=>x"a000", 252=>x"9b00",
---- 253=>x"9e00", 254=>x"9e00", 255=>x"9d00", 256=>x"a000",
---- 257=>x"9e00", 258=>x"9e00", 259=>x"9e00", 260=>x"9f00",
---- 261=>x"9e00", 262=>x"9d00", 263=>x"9f00", 264=>x"9e00",
---- 265=>x"9d00", 266=>x"9e00", 267=>x"9d00", 268=>x"9d00",
---- 269=>x"9d00", 270=>x"9b00", 271=>x"9d00", 272=>x"9f00",
---- 273=>x"9c00", 274=>x"9c00", 275=>x"9a00", 276=>x"9d00",
---- 277=>x"9e00", 278=>x"9c00", 279=>x"9b00", 280=>x"9d00",
---- 281=>x"9f00", 282=>x"9c00", 283=>x"9e00", 284=>x"9d00",
---- 285=>x"9d00", 286=>x"9d00", 287=>x"a000", 288=>x"9b00",
---- 289=>x"9c00", 290=>x"9c00", 291=>x"6200", 292=>x"9c00",
---- 293=>x"9d00", 294=>x"9c00", 295=>x"9e00", 296=>x"9c00",
---- 297=>x"9c00", 298=>x"9c00", 299=>x"9e00", 300=>x"9c00",
---- 301=>x"9f00", 302=>x"9f00", 303=>x"9e00", 304=>x"9d00",
---- 305=>x"9d00", 306=>x"9e00", 307=>x"a000", 308=>x"9d00",
---- 309=>x"9d00", 310=>x"9c00", 311=>x"9f00", 312=>x"9e00",
---- 313=>x"9d00", 314=>x"9f00", 315=>x"9d00", 316=>x"9d00",
---- 317=>x"9d00", 318=>x"9e00", 319=>x"6200", 320=>x"a000",
---- 321=>x"9c00", 322=>x"9b00", 323=>x"9c00", 324=>x"a000",
---- 325=>x"9c00", 326=>x"9d00", 327=>x"9d00", 328=>x"9b00",
---- 329=>x"9d00", 330=>x"9d00", 331=>x"9b00", 332=>x"9b00",
---- 333=>x"9d00", 334=>x"9d00", 335=>x"9c00", 336=>x"9d00",
---- 337=>x"9c00", 338=>x"9d00", 339=>x"6400", 340=>x"9c00",
---- 341=>x"9b00", 342=>x"9c00", 343=>x"9c00", 344=>x"9c00",
---- 345=>x"9c00", 346=>x"9b00", 347=>x"9c00", 348=>x"9b00",
---- 349=>x"9b00", 350=>x"9b00", 351=>x"9c00", 352=>x"9b00",
---- 353=>x"9900", 354=>x"9900", 355=>x"9900", 356=>x"9c00",
---- 357=>x"9b00", 358=>x"9a00", 359=>x"9b00", 360=>x"9a00",
---- 361=>x"9c00", 362=>x"9c00", 363=>x"9a00", 364=>x"9900",
---- 365=>x"9a00", 366=>x"9d00", 367=>x"9b00", 368=>x"9c00",
---- 369=>x"9a00", 370=>x"9800", 371=>x"9c00", 372=>x"9b00",
---- 373=>x"9a00", 374=>x"9900", 375=>x"9a00", 376=>x"9c00",
---- 377=>x"9c00", 378=>x"9c00", 379=>x"9b00", 380=>x"9c00",
---- 381=>x"9c00", 382=>x"9b00", 383=>x"9b00", 384=>x"9c00",
---- 385=>x"9c00", 386=>x"9a00", 387=>x"9d00", 388=>x"9b00",
---- 389=>x"9a00", 390=>x"9900", 391=>x"9b00", 392=>x"9d00",
---- 393=>x"9c00", 394=>x"9b00", 395=>x"9d00", 396=>x"9d00",
---- 397=>x"9c00", 398=>x"9b00", 399=>x"9c00", 400=>x"9e00",
---- 401=>x"9d00", 402=>x"9e00", 403=>x"9e00", 404=>x"9d00",
---- 405=>x"9e00", 406=>x"9c00", 407=>x"9c00", 408=>x"9e00",
---- 409=>x"9f00", 410=>x"9d00", 411=>x"9d00", 412=>x"a000",
---- 413=>x"9f00", 414=>x"6200", 415=>x"9d00", 416=>x"9f00",
---- 417=>x"9e00", 418=>x"9e00", 419=>x"9c00", 420=>x"9e00",
---- 421=>x"9d00", 422=>x"9e00", 423=>x"9e00", 424=>x"9d00",
---- 425=>x"9b00", 426=>x"9e00", 427=>x"9e00", 428=>x"a000",
---- 429=>x"9d00", 430=>x"9d00", 431=>x"9d00", 432=>x"a000",
---- 433=>x"9e00", 434=>x"a000", 435=>x"a000", 436=>x"9d00",
---- 437=>x"9d00", 438=>x"9d00", 439=>x"9e00", 440=>x"9e00",
---- 441=>x"9e00", 442=>x"9f00", 443=>x"9e00", 444=>x"9d00",
---- 445=>x"9d00", 446=>x"9f00", 447=>x"9e00", 448=>x"9c00",
---- 449=>x"9e00", 450=>x"9d00", 451=>x"9c00", 452=>x"9f00",
---- 453=>x"9d00", 454=>x"9d00", 455=>x"9c00", 456=>x"9f00",
---- 457=>x"9d00", 458=>x"9b00", 459=>x"9d00", 460=>x"9c00",
---- 461=>x"9d00", 462=>x"9c00", 463=>x"9a00", 464=>x"9a00",
---- 465=>x"9c00", 466=>x"9900", 467=>x"9900", 468=>x"9900",
---- 469=>x"9900", 470=>x"9900", 471=>x"9700", 472=>x"9300",
---- 473=>x"9500", 474=>x"9700", 475=>x"6600", 476=>x"8e00",
---- 477=>x"8f00", 478=>x"9000", 479=>x"9300", 480=>x"8e00",
---- 481=>x"9100", 482=>x"8d00", 483=>x"8d00", 484=>x"8e00",
---- 485=>x"9000", 486=>x"8e00", 487=>x"9000", 488=>x"6e00",
---- 489=>x"9000", 490=>x"9000", 491=>x"8d00", 492=>x"9600",
---- 493=>x"9100", 494=>x"8e00", 495=>x"8e00", 496=>x"9500",
---- 497=>x"9600", 498=>x"9100", 499=>x"8f00", 500=>x"9900",
---- 501=>x"9900", 502=>x"9200", 503=>x"9200", 504=>x"9a00",
---- 505=>x"9900", 506=>x"6700", 507=>x"9700", 508=>x"9e00",
---- 509=>x"9a00", 510=>x"9600", 511=>x"9600", 512=>x"9a00",
---- 513=>x"9600", 514=>x"9400", 515=>x"9100", 516=>x"9a00",
---- 517=>x"9800", 518=>x"9200", 519=>x"9300", 520=>x"9600",
---- 521=>x"9300", 522=>x"9300", 523=>x"9100", 524=>x"9300",
---- 525=>x"9100", 526=>x"9000", 527=>x"8f00", 528=>x"8f00",
---- 529=>x"8e00", 530=>x"8e00", 531=>x"8c00", 532=>x"8f00",
---- 533=>x"8e00", 534=>x"8d00", 535=>x"8b00", 536=>x"8c00",
---- 537=>x"8c00", 538=>x"8b00", 539=>x"8700", 540=>x"8900",
---- 541=>x"7600", 542=>x"8800", 543=>x"8400", 544=>x"8800",
---- 545=>x"8600", 546=>x"8500", 547=>x"8100", 548=>x"8600",
---- 549=>x"8400", 550=>x"8300", 551=>x"8600", 552=>x"8500",
---- 553=>x"7900", 554=>x"8f00", 555=>x"9d00", 556=>x"9000",
---- 557=>x"9b00", 558=>x"a500", 559=>x"ad00", 560=>x"a300",
---- 561=>x"ab00", 562=>x"b400", 563=>x"b900", 564=>x"b400",
---- 565=>x"b900", 566=>x"be00", 567=>x"c000", 568=>x"bf00",
---- 569=>x"c100", 570=>x"c100", 571=>x"c100", 572=>x"c500",
---- 573=>x"c600", 574=>x"c300", 575=>x"c000", 576=>x"c600",
---- 577=>x"c500", 578=>x"c300", 579=>x"c000", 580=>x"c600",
---- 581=>x"c400", 582=>x"c200", 583=>x"c000", 584=>x"c500",
---- 585=>x"c300", 586=>x"c200", 587=>x"c100", 588=>x"c500",
---- 589=>x"c300", 590=>x"c300", 591=>x"c200", 592=>x"c400",
---- 593=>x"c200", 594=>x"c100", 595=>x"c100", 596=>x"c400",
---- 597=>x"c300", 598=>x"c200", 599=>x"c300", 600=>x"c300",
---- 601=>x"c300", 602=>x"c200", 603=>x"c300", 604=>x"c200",
---- 605=>x"c200", 606=>x"c400", 607=>x"c700", 608=>x"c300",
---- 609=>x"c300", 610=>x"c600", 611=>x"ca00", 612=>x"c500",
---- 613=>x"c700", 614=>x"cc00", 615=>x"cd00", 616=>x"c900",
---- 617=>x"cc00", 618=>x"ce00", 619=>x"d000", 620=>x"cd00",
---- 621=>x"3000", 622=>x"ce00", 623=>x"cf00", 624=>x"2f00",
---- 625=>x"d200", 626=>x"d000", 627=>x"ce00", 628=>x"d100",
---- 629=>x"d100", 630=>x"d000", 631=>x"ce00", 632=>x"d000",
---- 633=>x"cf00", 634=>x"ce00", 635=>x"cd00", 636=>x"cf00",
---- 637=>x"ce00", 638=>x"cd00", 639=>x"cc00", 640=>x"cf00",
---- 641=>x"cd00", 642=>x"ce00", 643=>x"ce00", 644=>x"ce00",
---- 645=>x"ce00", 646=>x"d000", 647=>x"d000", 648=>x"cf00",
---- 649=>x"d000", 650=>x"d000", 651=>x"d300", 652=>x"cf00",
---- 653=>x"cf00", 654=>x"cf00", 655=>x"d400", 656=>x"ce00",
---- 657=>x"cf00", 658=>x"2d00", 659=>x"d400", 660=>x"cf00",
---- 661=>x"ce00", 662=>x"d200", 663=>x"d100", 664=>x"2e00",
---- 665=>x"d100", 666=>x"d100", 667=>x"d300", 668=>x"d000",
---- 669=>x"cf00", 670=>x"d000", 671=>x"d200", 672=>x"cf00",
---- 673=>x"d000", 674=>x"d100", 675=>x"d200", 676=>x"d000",
---- 677=>x"cf00", 678=>x"cf00", 679=>x"d100", 680=>x"d100",
---- 681=>x"cf00", 682=>x"cf00", 683=>x"d200", 684=>x"cf00",
---- 685=>x"cf00", 686=>x"d100", 687=>x"d300", 688=>x"d000",
---- 689=>x"2f00", 690=>x"d200", 691=>x"d200", 692=>x"d100",
---- 693=>x"d100", 694=>x"d200", 695=>x"d300", 696=>x"d300",
---- 697=>x"d300", 698=>x"2a00", 699=>x"d500", 700=>x"d300",
---- 701=>x"d300", 702=>x"d300", 703=>x"d300", 704=>x"d300",
---- 705=>x"d200", 706=>x"d300", 707=>x"d500", 708=>x"d400",
---- 709=>x"d500", 710=>x"d600", 711=>x"d500", 712=>x"d500",
---- 713=>x"d500", 714=>x"d400", 715=>x"d600", 716=>x"d600",
---- 717=>x"d600", 718=>x"d500", 719=>x"d500", 720=>x"d800",
---- 721=>x"d700", 722=>x"d500", 723=>x"d200", 724=>x"d700",
---- 725=>x"d500", 726=>x"d100", 727=>x"cf00", 728=>x"d300",
---- 729=>x"d000", 730=>x"ce00", 731=>x"cd00", 732=>x"d100",
---- 733=>x"ce00", 734=>x"cd00", 735=>x"cf00", 736=>x"d000",
---- 737=>x"d000", 738=>x"d100", 739=>x"d200", 740=>x"d200",
---- 741=>x"d300", 742=>x"d400", 743=>x"d400", 744=>x"d600",
---- 745=>x"d500", 746=>x"d500", 747=>x"d400", 748=>x"d400",
---- 749=>x"d400", 750=>x"d200", 751=>x"d200", 752=>x"d200",
---- 753=>x"d200", 754=>x"d000", 755=>x"cf00", 756=>x"d200",
---- 757=>x"cf00", 758=>x"cd00", 759=>x"cf00", 760=>x"cf00",
---- 761=>x"cd00", 762=>x"ce00", 763=>x"cc00", 764=>x"cd00",
---- 765=>x"ce00", 766=>x"cd00", 767=>x"cc00", 768=>x"cd00",
---- 769=>x"ca00", 770=>x"c500", 771=>x"c100", 772=>x"3800",
---- 773=>x"bf00", 774=>x"b100", 775=>x"a200", 776=>x"b700",
---- 777=>x"a700", 778=>x"8b00", 779=>x"6400", 780=>x"a500",
---- 781=>x"8b00", 782=>x"6200", 783=>x"3a00", 784=>x"9600",
---- 785=>x"7400", 786=>x"4700", 787=>x"3100", 788=>x"7e00",
---- 789=>x"4d00", 790=>x"2f00", 791=>x"2a00", 792=>x"4a00",
---- 793=>x"2c00", 794=>x"2700", 795=>x"2d00", 796=>x"d200",
---- 797=>x"2e00", 798=>x"3200", 799=>x"3c00", 800=>x"3300",
---- 801=>x"3f00", 802=>x"4300", 803=>x"4600", 804=>x"4400",
---- 805=>x"5000", 806=>x"4f00", 807=>x"4b00", 808=>x"5000",
---- 809=>x"4f00", 810=>x"4f00", 811=>x"5000", 812=>x"5500",
---- 813=>x"4f00", 814=>x"4d00", 815=>x"4d00", 816=>x"5600",
---- 817=>x"5400", 818=>x"5000", 819=>x"5200", 820=>x"5600",
---- 821=>x"5600", 822=>x"5500", 823=>x"5a00", 824=>x"6000",
---- 825=>x"5800", 826=>x"5500", 827=>x"6300", 828=>x"5c00",
---- 829=>x"5b00", 830=>x"6100", 831=>x"6e00", 832=>x"5c00",
---- 833=>x"6000", 834=>x"6900", 835=>x"6e00", 836=>x"6200",
---- 837=>x"6800", 838=>x"6f00", 839=>x"7400", 840=>x"6500",
---- 841=>x"6f00", 842=>x"7500", 843=>x"6f00", 844=>x"6b00",
---- 845=>x"7200", 846=>x"6b00", 847=>x"6200", 848=>x"7100",
---- 849=>x"7100", 850=>x"6600", 851=>x"5d00", 852=>x"7000",
---- 853=>x"6b00", 854=>x"6100", 855=>x"5a00", 856=>x"6f00",
---- 857=>x"6500", 858=>x"5b00", 859=>x"5800", 860=>x"6c00",
---- 861=>x"5f00", 862=>x"5d00", 863=>x"5b00", 864=>x"6800",
---- 865=>x"5c00", 866=>x"5900", 867=>x"5b00", 868=>x"6300",
---- 869=>x"5c00", 870=>x"5700", 871=>x"5b00", 872=>x"5f00",
---- 873=>x"5c00", 874=>x"5a00", 875=>x"6000", 876=>x"5c00",
---- 877=>x"5b00", 878=>x"5e00", 879=>x"6400", 880=>x"5c00",
---- 881=>x"5b00", 882=>x"a100", 883=>x"6400", 884=>x"5a00",
---- 885=>x"5c00", 886=>x"6000", 887=>x"6a00", 888=>x"5a00",
---- 889=>x"5a00", 890=>x"6200", 891=>x"6b00", 892=>x"5500",
---- 893=>x"6000", 894=>x"6700", 895=>x"6900", 896=>x"5c00",
---- 897=>x"6400", 898=>x"6a00", 899=>x"6800", 900=>x"6600",
---- 901=>x"6900", 902=>x"6500", 903=>x"9a00", 904=>x"6900",
---- 905=>x"6600", 906=>x"6500", 907=>x"6100", 908=>x"6c00",
---- 909=>x"6300", 910=>x"6600", 911=>x"5c00", 912=>x"6900",
---- 913=>x"6100", 914=>x"5d00", 915=>x"5a00", 916=>x"6500",
---- 917=>x"6000", 918=>x"5d00", 919=>x"5600", 920=>x"6100",
---- 921=>x"6100", 922=>x"5800", 923=>x"5900", 924=>x"6000",
---- 925=>x"5f00", 926=>x"5900", 927=>x"5a00", 928=>x"5e00",
---- 929=>x"5d00", 930=>x"5d00", 931=>x"5c00", 932=>x"5d00",
---- 933=>x"5b00", 934=>x"5d00", 935=>x"6300", 936=>x"5c00",
---- 937=>x"5900", 938=>x"5e00", 939=>x"6500", 940=>x"5d00",
---- 941=>x"5a00", 942=>x"5e00", 943=>x"6600", 944=>x"5a00",
---- 945=>x"5d00", 946=>x"6200", 947=>x"6700", 948=>x"5700",
---- 949=>x"5e00", 950=>x"6800", 951=>x"6a00", 952=>x"5600",
---- 953=>x"6300", 954=>x"6c00", 955=>x"7100", 956=>x"5b00",
---- 957=>x"6900", 958=>x"7300", 959=>x"6d00", 960=>x"6300",
---- 961=>x"6c00", 962=>x"7400", 963=>x"6900", 964=>x"6a00",
---- 965=>x"7200", 966=>x"6d00", 967=>x"6300", 968=>x"7200",
---- 969=>x"7000", 970=>x"6700", 971=>x"5c00", 972=>x"7300",
---- 973=>x"6a00", 974=>x"6700", 975=>x"6000", 976=>x"6f00",
---- 977=>x"9400", 978=>x"6500", 979=>x"6100", 980=>x"7000",
---- 981=>x"6a00", 982=>x"6600", 983=>x"6200", 984=>x"7400",
---- 985=>x"6800", 986=>x"6500", 987=>x"5d00", 988=>x"7100",
---- 989=>x"6b00", 990=>x"6500", 991=>x"5700", 992=>x"6a00",
---- 993=>x"6800", 994=>x"5f00", 995=>x"4e00", 996=>x"6b00",
---- 997=>x"6200", 998=>x"5500", 999=>x"4700", 1000=>x"6100",
---- 1001=>x"5a00", 1002=>x"5000", 1003=>x"4300", 1004=>x"5b00",
---- 1005=>x"5300", 1006=>x"4700", 1007=>x"3f00", 1008=>x"5600",
---- 1009=>x"4a00", 1010=>x"3d00", 1011=>x"3600", 1012=>x"4b00",
---- 1013=>x"3d00", 1014=>x"3a00", 1015=>x"2f00", 1016=>x"3d00",
---- 1017=>x"3300", 1018=>x"3200", 1019=>x"3100", 1020=>x"3a00",
---- 1021=>x"3400", 1022=>x"2c00", 1023=>x"2b00"),
----
---- 62 => (0=>x"7600", 1=>x"7700", 2=>x"7500", 3=>x"7500", 4=>x"7500",
---- 5=>x"7600", 6=>x"7500", 7=>x"7500", 8=>x"7600",
---- 9=>x"7500", 10=>x"7700", 11=>x"7700", 12=>x"7800",
---- 13=>x"7700", 14=>x"7e00", 15=>x"7f00", 16=>x"7e00",
---- 17=>x"7e00", 18=>x"8000", 19=>x"7a00", 20=>x"8400",
---- 21=>x"8100", 22=>x"7400", 23=>x"5a00", 24=>x"8500",
---- 25=>x"7a00", 26=>x"5c00", 27=>x"3c00", 28=>x"7100",
---- 29=>x"5700", 30=>x"3600", 31=>x"3600", 32=>x"4f00",
---- 33=>x"3200", 34=>x"2d00", 35=>x"2a00", 36=>x"3000",
---- 37=>x"2c00", 38=>x"3000", 39=>x"2e00", 40=>x"2a00",
---- 41=>x"3200", 42=>x"3400", 43=>x"2f00", 44=>x"2f00",
---- 45=>x"d200", 46=>x"3600", 47=>x"3300", 48=>x"3200",
---- 49=>x"2e00", 50=>x"2c00", 51=>x"d100", 52=>x"2800",
---- 53=>x"2d00", 54=>x"2a00", 55=>x"2e00", 56=>x"2b00",
---- 57=>x"2e00", 58=>x"2f00", 59=>x"3000", 60=>x"3100",
---- 61=>x"2e00", 62=>x"3200", 63=>x"3300", 64=>x"3100",
---- 65=>x"3300", 66=>x"3500", 67=>x"3200", 68=>x"3600",
---- 69=>x"3200", 70=>x"3500", 71=>x"3300", 72=>x"3200",
---- 73=>x"3200", 74=>x"3500", 75=>x"3100", 76=>x"3900",
---- 77=>x"3600", 78=>x"3500", 79=>x"3400", 80=>x"3400",
---- 81=>x"3400", 82=>x"3200", 83=>x"2f00", 84=>x"3300",
---- 85=>x"3500", 86=>x"3200", 87=>x"3000", 88=>x"3500",
---- 89=>x"3300", 90=>x"3600", 91=>x"2e00", 92=>x"ca00",
---- 93=>x"3200", 94=>x"3400", 95=>x"2f00", 96=>x"3400",
---- 97=>x"2d00", 98=>x"2a00", 99=>x"2b00", 100=>x"cd00",
---- 101=>x"2b00", 102=>x"2a00", 103=>x"2b00", 104=>x"2f00",
---- 105=>x"2c00", 106=>x"2f00", 107=>x"3000", 108=>x"3100",
---- 109=>x"3500", 110=>x"3500", 111=>x"3100", 112=>x"c900",
---- 113=>x"3700", 114=>x"3000", 115=>x"2d00", 116=>x"3600",
---- 117=>x"3100", 118=>x"2e00", 119=>x"3200", 120=>x"3300",
---- 121=>x"3100", 122=>x"2d00", 123=>x"3300", 124=>x"3000",
---- 125=>x"2f00", 126=>x"2a00", 127=>x"2e00", 128=>x"3000",
---- 129=>x"2b00", 130=>x"2c00", 131=>x"2c00", 132=>x"2e00",
---- 133=>x"2d00", 134=>x"2f00", 135=>x"3100", 136=>x"2c00",
---- 137=>x"2d00", 138=>x"3300", 139=>x"3900", 140=>x"3000",
---- 141=>x"3000", 142=>x"3a00", 143=>x"4300", 144=>x"3300",
---- 145=>x"3b00", 146=>x"4800", 147=>x"4300", 148=>x"3800",
---- 149=>x"4300", 150=>x"4200", 151=>x"3100", 152=>x"4500",
---- 153=>x"4300", 154=>x"3200", 155=>x"2700", 156=>x"4f00",
---- 157=>x"4100", 158=>x"2900", 159=>x"2500", 160=>x"5300",
---- 161=>x"3e00", 162=>x"2900", 163=>x"3000", 164=>x"4b00",
---- 165=>x"3600", 166=>x"2f00", 167=>x"5400", 168=>x"3e00",
---- 169=>x"3c00", 170=>x"5400", 171=>x"7900", 172=>x"3e00",
---- 173=>x"5600", 174=>x"7800", 175=>x"8b00", 176=>x"5b00",
---- 177=>x"7600", 178=>x"8b00", 179=>x"9600", 180=>x"7100",
---- 181=>x"8800", 182=>x"9300", 183=>x"9600", 184=>x"8300",
---- 185=>x"8f00", 186=>x"9300", 187=>x"9600", 188=>x"6e00",
---- 189=>x"9400", 190=>x"9300", 191=>x"9700", 192=>x"9500",
---- 193=>x"9700", 194=>x"9100", 195=>x"8b00", 196=>x"9500",
---- 197=>x"9700", 198=>x"8f00", 199=>x"8a00", 200=>x"9600",
---- 201=>x"9700", 202=>x"8b00", 203=>x"9600", 204=>x"9300",
---- 205=>x"8d00", 206=>x"9400", 207=>x"9f00", 208=>x"8800",
---- 209=>x"8d00", 210=>x"9c00", 211=>x"a400", 212=>x"8e00",
---- 213=>x"9b00", 214=>x"a000", 215=>x"a500", 216=>x"9900",
---- 217=>x"9e00", 218=>x"a200", 219=>x"a100", 220=>x"9e00",
---- 221=>x"9e00", 222=>x"a300", 223=>x"a300", 224=>x"a000",
---- 225=>x"a200", 226=>x"a300", 227=>x"a100", 228=>x"a200",
---- 229=>x"a200", 230=>x"a000", 231=>x"a000", 232=>x"a100",
---- 233=>x"a100", 234=>x"a000", 235=>x"a000", 236=>x"a100",
---- 237=>x"a000", 238=>x"9e00", 239=>x"9f00", 240=>x"9f00",
---- 241=>x"a000", 242=>x"a000", 243=>x"a000", 244=>x"a100",
---- 245=>x"a000", 246=>x"9e00", 247=>x"9f00", 248=>x"a000",
---- 249=>x"a000", 250=>x"9e00", 251=>x"9f00", 252=>x"9f00",
---- 253=>x"9f00", 254=>x"9f00", 255=>x"9b00", 256=>x"9e00",
---- 257=>x"6300", 258=>x"9d00", 259=>x"9d00", 260=>x"9e00",
---- 261=>x"9f00", 262=>x"9e00", 263=>x"9b00", 264=>x"9e00",
---- 265=>x"9d00", 266=>x"9c00", 267=>x"9d00", 268=>x"9c00",
---- 269=>x"9b00", 270=>x"9c00", 271=>x"9a00", 272=>x"9d00",
---- 273=>x"9d00", 274=>x"9b00", 275=>x"9c00", 276=>x"9e00",
---- 277=>x"9d00", 278=>x"9c00", 279=>x"9b00", 280=>x"9c00",
---- 281=>x"9a00", 282=>x"9c00", 283=>x"9b00", 284=>x"9e00",
---- 285=>x"9a00", 286=>x"9a00", 287=>x"9800", 288=>x"9b00",
---- 289=>x"9900", 290=>x"9c00", 291=>x"9b00", 292=>x"9c00",
---- 293=>x"6500", 294=>x"9c00", 295=>x"9c00", 296=>x"9c00",
---- 297=>x"9b00", 298=>x"9b00", 299=>x"9b00", 300=>x"9d00",
---- 301=>x"9d00", 302=>x"9f00", 303=>x"9a00", 304=>x"9e00",
---- 305=>x"9e00", 306=>x"9e00", 307=>x"9f00", 308=>x"9d00",
---- 309=>x"9d00", 310=>x"9c00", 311=>x"a000", 312=>x"9c00",
---- 313=>x"9e00", 314=>x"9f00", 315=>x"9f00", 316=>x"9e00",
---- 317=>x"9d00", 318=>x"9f00", 319=>x"9f00", 320=>x"9e00",
---- 321=>x"9c00", 322=>x"9e00", 323=>x"9d00", 324=>x"9c00",
---- 325=>x"9a00", 326=>x"9d00", 327=>x"9e00", 328=>x"9e00",
---- 329=>x"9c00", 330=>x"9f00", 331=>x"9c00", 332=>x"9d00",
---- 333=>x"9d00", 334=>x"9c00", 335=>x"9c00", 336=>x"9c00",
---- 337=>x"9c00", 338=>x"9e00", 339=>x"9d00", 340=>x"9c00",
---- 341=>x"6100", 342=>x"9b00", 343=>x"9c00", 344=>x"9a00",
---- 345=>x"9d00", 346=>x"9d00", 347=>x"9c00", 348=>x"9b00",
---- 349=>x"9c00", 350=>x"9b00", 351=>x"9c00", 352=>x"9a00",
---- 353=>x"9b00", 354=>x"9900", 355=>x"9a00", 356=>x"9a00",
---- 357=>x"9a00", 358=>x"9b00", 359=>x"9a00", 360=>x"9b00",
---- 361=>x"9800", 362=>x"9a00", 363=>x"9900", 364=>x"9a00",
---- 365=>x"9b00", 366=>x"9b00", 367=>x"9a00", 368=>x"9c00",
---- 369=>x"9b00", 370=>x"9a00", 371=>x"9a00", 372=>x"9900",
---- 373=>x"9800", 374=>x"9900", 375=>x"9900", 376=>x"9a00",
---- 377=>x"9900", 378=>x"9c00", 379=>x"9b00", 380=>x"9a00",
---- 381=>x"9a00", 382=>x"9b00", 383=>x"9a00", 384=>x"9b00",
---- 385=>x"9c00", 386=>x"9b00", 387=>x"9b00", 388=>x"9d00",
---- 389=>x"9c00", 390=>x"9c00", 391=>x"9a00", 392=>x"9b00",
---- 393=>x"9900", 394=>x"9b00", 395=>x"9900", 396=>x"9b00",
---- 397=>x"9a00", 398=>x"9a00", 399=>x"9800", 400=>x"9c00",
---- 401=>x"9b00", 402=>x"9c00", 403=>x"9900", 404=>x"9c00",
---- 405=>x"9c00", 406=>x"9a00", 407=>x"9800", 408=>x"9d00",
---- 409=>x"9a00", 410=>x"9b00", 411=>x"9a00", 412=>x"9d00",
---- 413=>x"9d00", 414=>x"9b00", 415=>x"9a00", 416=>x"9b00",
---- 417=>x"9c00", 418=>x"9c00", 419=>x"9900", 420=>x"9d00",
---- 421=>x"9c00", 422=>x"9d00", 423=>x"9900", 424=>x"9c00",
---- 425=>x"9c00", 426=>x"9d00", 427=>x"9a00", 428=>x"9e00",
---- 429=>x"9d00", 430=>x"9c00", 431=>x"9a00", 432=>x"9e00",
---- 433=>x"9e00", 434=>x"9d00", 435=>x"9e00", 436=>x"9c00",
---- 437=>x"9f00", 438=>x"9e00", 439=>x"9b00", 440=>x"9d00",
---- 441=>x"9e00", 442=>x"9b00", 443=>x"9a00", 444=>x"9d00",
---- 445=>x"6000", 446=>x"9d00", 447=>x"9b00", 448=>x"9d00",
---- 449=>x"9d00", 450=>x"9c00", 451=>x"9c00", 452=>x"9c00",
---- 453=>x"9c00", 454=>x"9c00", 455=>x"9a00", 456=>x"9d00",
---- 457=>x"9b00", 458=>x"9b00", 459=>x"9b00", 460=>x"9b00",
---- 461=>x"9a00", 462=>x"9c00", 463=>x"9a00", 464=>x"9a00",
---- 465=>x"9900", 466=>x"9a00", 467=>x"9b00", 468=>x"9700",
---- 469=>x"9800", 470=>x"9800", 471=>x"9b00", 472=>x"9800",
---- 473=>x"9500", 474=>x"9a00", 475=>x"9b00", 476=>x"9400",
---- 477=>x"9900", 478=>x"9a00", 479=>x"9800", 480=>x"9000",
---- 481=>x"9300", 482=>x"9600", 483=>x"9600", 484=>x"8c00",
---- 485=>x"8d00", 486=>x"8f00", 487=>x"9000", 488=>x"8c00",
---- 489=>x"8f00", 490=>x"8f00", 491=>x"8c00", 492=>x"8d00",
---- 493=>x"8e00", 494=>x"8d00", 495=>x"8c00", 496=>x"8e00",
---- 497=>x"8e00", 498=>x"8f00", 499=>x"7300", 500=>x"9000",
---- 501=>x"8f00", 502=>x"9000", 503=>x"8b00", 504=>x"9400",
---- 505=>x"9100", 506=>x"8f00", 507=>x"8d00", 508=>x"9900",
---- 509=>x"9800", 510=>x"9300", 511=>x"8e00", 512=>x"9400",
---- 513=>x"9500", 514=>x"9300", 515=>x"9100", 516=>x"9100",
---- 517=>x"9100", 518=>x"9200", 519=>x"8e00", 520=>x"9100",
---- 521=>x"9000", 522=>x"9000", 523=>x"8f00", 524=>x"8f00",
---- 525=>x"8a00", 526=>x"8900", 527=>x"8a00", 528=>x"8a00",
---- 529=>x"8900", 530=>x"8600", 531=>x"8700", 532=>x"8800",
---- 533=>x"8400", 534=>x"8700", 535=>x"8400", 536=>x"7b00",
---- 537=>x"8400", 538=>x"8100", 539=>x"8000", 540=>x"8200",
---- 541=>x"8000", 542=>x"8100", 543=>x"7c00", 544=>x"8200",
---- 545=>x"8700", 546=>x"9100", 547=>x"9900", 548=>x"9300",
---- 549=>x"9e00", 550=>x"a300", 551=>x"ac00", 552=>x"a500",
---- 553=>x"ae00", 554=>x"b200", 555=>x"b500", 556=>x"b300",
---- 557=>x"b700", 558=>x"bd00", 559=>x"bc00", 560=>x"bd00",
---- 561=>x"bd00", 562=>x"be00", 563=>x"be00", 564=>x"c000",
---- 565=>x"c000", 566=>x"be00", 567=>x"bd00", 568=>x"c100",
---- 569=>x"c000", 570=>x"c000", 571=>x"bd00", 572=>x"bf00",
---- 573=>x"bf00", 574=>x"bf00", 575=>x"bd00", 576=>x"c000",
---- 577=>x"bf00", 578=>x"bc00", 579=>x"bc00", 580=>x"c000",
---- 581=>x"be00", 582=>x"bd00", 583=>x"bc00", 584=>x"be00",
---- 585=>x"bf00", 586=>x"be00", 587=>x"be00", 588=>x"c000",
---- 589=>x"bf00", 590=>x"bd00", 591=>x"c000", 592=>x"c300",
---- 593=>x"c000", 594=>x"c100", 595=>x"c300", 596=>x"c300",
---- 597=>x"c100", 598=>x"c500", 599=>x"c600", 600=>x"c500",
---- 601=>x"c800", 602=>x"ca00", 603=>x"ca00", 604=>x"ca00",
---- 605=>x"cb00", 606=>x"cd00", 607=>x"ce00", 608=>x"cc00",
---- 609=>x"d000", 610=>x"d000", 611=>x"ce00", 612=>x"d000",
---- 613=>x"d300", 614=>x"d100", 615=>x"cf00", 616=>x"d100",
---- 617=>x"d100", 618=>x"d100", 619=>x"cf00", 620=>x"d100",
---- 621=>x"cf00", 622=>x"d000", 623=>x"d000", 624=>x"cf00",
---- 625=>x"ce00", 626=>x"d100", 627=>x"cf00", 628=>x"cc00",
---- 629=>x"ce00", 630=>x"ce00", 631=>x"cf00", 632=>x"cc00",
---- 633=>x"ce00", 634=>x"ce00", 635=>x"ce00", 636=>x"cd00",
---- 637=>x"cd00", 638=>x"cf00", 639=>x"cf00", 640=>x"cd00",
---- 641=>x"ce00", 642=>x"cf00", 643=>x"d100", 644=>x"cf00",
---- 645=>x"d200", 646=>x"d100", 647=>x"d100", 648=>x"d200",
---- 649=>x"d100", 650=>x"d200", 651=>x"d100", 652=>x"d200",
---- 653=>x"d100", 654=>x"d200", 655=>x"2c00", 656=>x"d300",
---- 657=>x"d100", 658=>x"d200", 659=>x"d200", 660=>x"d200",
---- 661=>x"d200", 662=>x"d300", 663=>x"d100", 664=>x"d100",
---- 665=>x"d100", 666=>x"d400", 667=>x"d100", 668=>x"d200",
---- 669=>x"d200", 670=>x"d300", 671=>x"d200", 672=>x"d000",
---- 673=>x"d300", 674=>x"d300", 675=>x"d300", 676=>x"d200",
---- 677=>x"d500", 678=>x"d300", 679=>x"d000", 680=>x"d200",
---- 681=>x"d500", 682=>x"d400", 683=>x"d100", 684=>x"d400",
---- 685=>x"d300", 686=>x"d400", 687=>x"d400", 688=>x"d500",
---- 689=>x"d500", 690=>x"d500", 691=>x"d300", 692=>x"d500",
---- 693=>x"d500", 694=>x"d700", 695=>x"d400", 696=>x"d500",
---- 697=>x"d500", 698=>x"d500", 699=>x"d500", 700=>x"2b00",
---- 701=>x"d600", 702=>x"d700", 703=>x"d500", 704=>x"d500",
---- 705=>x"d600", 706=>x"d700", 707=>x"d600", 708=>x"d600",
---- 709=>x"d400", 710=>x"d500", 711=>x"d500", 712=>x"d600",
---- 713=>x"d600", 714=>x"d400", 715=>x"d300", 716=>x"d600",
---- 717=>x"d300", 718=>x"d200", 719=>x"d200", 720=>x"d200",
---- 721=>x"d000", 722=>x"cf00", 723=>x"cf00", 724=>x"cf00",
---- 725=>x"cd00", 726=>x"cd00", 727=>x"cc00", 728=>x"3100",
---- 729=>x"cd00", 730=>x"cd00", 731=>x"cd00", 732=>x"d000",
---- 733=>x"d000", 734=>x"d100", 735=>x"d100", 736=>x"2e00",
---- 737=>x"d000", 738=>x"d300", 739=>x"d200", 740=>x"d300",
---- 741=>x"d300", 742=>x"d200", 743=>x"d200", 744=>x"d200",
---- 745=>x"d100", 746=>x"d100", 747=>x"cf00", 748=>x"d100",
---- 749=>x"d000", 750=>x"cf00", 751=>x"cf00", 752=>x"cf00",
---- 753=>x"cf00", 754=>x"cf00", 755=>x"cf00", 756=>x"cd00",
---- 757=>x"cb00", 758=>x"cc00", 759=>x"cc00", 760=>x"cb00",
---- 761=>x"c900", 762=>x"c700", 763=>x"3900", 764=>x"c800",
---- 765=>x"c400", 766=>x"b800", 767=>x"af00", 768=>x"ba00",
---- 769=>x"aa00", 770=>x"8e00", 771=>x"6700", 772=>x"8700",
---- 773=>x"6100", 774=>x"4000", 775=>x"2d00", 776=>x"3f00",
---- 777=>x"2e00", 778=>x"2900", 779=>x"2a00", 780=>x"2a00",
---- 781=>x"2b00", 782=>x"2a00", 783=>x"2c00", 784=>x"2a00",
---- 785=>x"2700", 786=>x"2a00", 787=>x"3400", 788=>x"2e00",
---- 789=>x"3300", 790=>x"3800", 791=>x"4000", 792=>x"3600",
---- 793=>x"3c00", 794=>x"4100", 795=>x"4b00", 796=>x"3f00",
---- 797=>x"4000", 798=>x"4600", 799=>x"5100", 800=>x"4600",
---- 801=>x"4a00", 802=>x"4f00", 803=>x"5300", 804=>x"4c00",
---- 805=>x"4d00", 806=>x"5400", 807=>x"5600", 808=>x"5200",
---- 809=>x"5600", 810=>x"5900", 811=>x"5b00", 812=>x"5500",
---- 813=>x"5c00", 814=>x"5d00", 815=>x"6100", 816=>x"5e00",
---- 817=>x"6000", 818=>x"6500", 819=>x"6200", 820=>x"6400",
---- 821=>x"6600", 822=>x"6800", 823=>x"5f00", 824=>x"6a00",
---- 825=>x"7100", 826=>x"6800", 827=>x"6200", 828=>x"8d00",
---- 829=>x"7100", 830=>x"6700", 831=>x"6000", 832=>x"6f00",
---- 833=>x"6b00", 834=>x"6500", 835=>x"5e00", 836=>x"6f00",
---- 837=>x"6200", 838=>x"5e00", 839=>x"5d00", 840=>x"6300",
---- 841=>x"5900", 842=>x"5c00", 843=>x"5d00", 844=>x"5a00",
---- 845=>x"5800", 846=>x"5b00", 847=>x"6300", 848=>x"5700",
---- 849=>x"5800", 850=>x"5b00", 851=>x"6500", 852=>x"5800",
---- 853=>x"5b00", 854=>x"6000", 855=>x"6800", 856=>x"5b00",
---- 857=>x"5e00", 858=>x"6500", 859=>x"6a00", 860=>x"5b00",
---- 861=>x"6300", 862=>x"6600", 863=>x"6800", 864=>x"5e00",
---- 865=>x"6800", 866=>x"6800", 867=>x"6900", 868=>x"6500",
---- 869=>x"6800", 870=>x"6a00", 871=>x"6600", 872=>x"6800",
---- 873=>x"6900", 874=>x"6800", 875=>x"6700", 876=>x"6a00",
---- 877=>x"6a00", 878=>x"6800", 879=>x"6500", 880=>x"6800",
---- 881=>x"6800", 882=>x"6700", 883=>x"6100", 884=>x"6500",
---- 885=>x"6a00", 886=>x"6400", 887=>x"5e00", 888=>x"6600",
---- 889=>x"6500", 890=>x"6200", 891=>x"6200", 892=>x"6900",
---- 893=>x"5d00", 894=>x"5c00", 895=>x"6000", 896=>x"6700",
---- 897=>x"5f00", 898=>x"5e00", 899=>x"6000", 900=>x"6200",
---- 901=>x"5c00", 902=>x"6200", 903=>x"5e00", 904=>x"5a00",
---- 905=>x"5a00", 906=>x"5f00", 907=>x"a300", 908=>x"5800",
---- 909=>x"5b00", 910=>x"5d00", 911=>x"6000", 912=>x"5800",
---- 913=>x"5800", 914=>x"5d00", 915=>x"6200", 916=>x"5900",
---- 917=>x"5a00", 918=>x"6000", 919=>x"5e00", 920=>x"5e00",
---- 921=>x"6300", 922=>x"6500", 923=>x"5d00", 924=>x"6300",
---- 925=>x"6a00", 926=>x"6300", 927=>x"5c00", 928=>x"6500",
---- 929=>x"6b00", 930=>x"6100", 931=>x"5e00", 932=>x"6800",
---- 933=>x"6500", 934=>x"6100", 935=>x"5e00", 936=>x"6900",
---- 937=>x"5e00", 938=>x"6000", 939=>x"5a00", 940=>x"6500",
---- 941=>x"6200", 942=>x"5e00", 943=>x"a700", 944=>x"6400",
---- 945=>x"6200", 946=>x"5a00", 947=>x"b100", 948=>x"6700",
---- 949=>x"5f00", 950=>x"5500", 951=>x"4600", 952=>x"6600",
---- 953=>x"5a00", 954=>x"5400", 955=>x"4800", 956=>x"6300",
---- 957=>x"5d00", 958=>x"5200", 959=>x"4d00", 960=>x"6000",
---- 961=>x"5700", 962=>x"5200", 963=>x"5500", 964=>x"5f00",
---- 965=>x"a800", 966=>x"5000", 967=>x"4b00", 968=>x"5e00",
---- 969=>x"5900", 970=>x"4f00", 971=>x"4700", 972=>x"5d00",
---- 973=>x"5600", 974=>x"4c00", 975=>x"3e00", 976=>x"5c00",
---- 977=>x"4b00", 978=>x"3f00", 979=>x"3b00", 980=>x"5500",
---- 981=>x"4400", 982=>x"3d00", 983=>x"4400", 984=>x"4b00",
---- 985=>x"4300", 986=>x"4100", 987=>x"3e00", 988=>x"4b00",
---- 989=>x"4400", 990=>x"3f00", 991=>x"3d00", 992=>x"b700",
---- 993=>x"4100", 994=>x"3a00", 995=>x"3b00", 996=>x"3e00",
---- 997=>x"3a00", 998=>x"3b00", 999=>x"3900", 1000=>x"3d00",
---- 1001=>x"3900", 1002=>x"3800", 1003=>x"3b00", 1004=>x"3800",
---- 1005=>x"3700", 1006=>x"3d00", 1007=>x"3700", 1008=>x"3200",
---- 1009=>x"3300", 1010=>x"3a00", 1011=>x"c200", 1012=>x"2f00",
---- 1013=>x"3600", 1014=>x"3400", 1015=>x"3d00", 1016=>x"3300",
---- 1017=>x"3200", 1018=>x"3700", 1019=>x"3c00", 1020=>x"3000",
---- 1021=>x"3300", 1022=>x"3f00", 1023=>x"4b00"),
----
---- 63 => (0=>x"8c00", 1=>x"a900", 2=>x"ac00", 3=>x"9500", 4=>x"8d00",
---- 5=>x"a900", 6=>x"ae00", 7=>x"9900", 8=>x"8c00",
---- 9=>x"a700", 10=>x"a800", 11=>x"8c00", 12=>x"7f00",
---- 13=>x"7700", 14=>x"6000", 15=>x"4300", 16=>x"5f00",
---- 17=>x"3c00", 18=>x"2f00", 19=>x"2d00", 20=>x"3c00",
---- 21=>x"2f00", 22=>x"2f00", 23=>x"3000", 24=>x"3100",
---- 25=>x"2900", 26=>x"2e00", 27=>x"3000", 28=>x"3600",
---- 29=>x"2c00", 30=>x"3300", 31=>x"3200", 32=>x"2e00",
---- 33=>x"3000", 34=>x"2d00", 35=>x"2f00", 36=>x"3200",
---- 37=>x"3100", 38=>x"2c00", 39=>x"2f00", 40=>x"3300",
---- 41=>x"3000", 42=>x"2e00", 43=>x"3100", 44=>x"2e00",
---- 45=>x"2e00", 46=>x"3100", 47=>x"3400", 48=>x"2e00",
---- 49=>x"3200", 50=>x"3300", 51=>x"3500", 52=>x"2d00",
---- 53=>x"3200", 54=>x"3800", 55=>x"3300", 56=>x"2f00",
---- 57=>x"3400", 58=>x"3200", 59=>x"3900", 60=>x"3300",
---- 61=>x"3100", 62=>x"3200", 63=>x"3800", 64=>x"3200",
---- 65=>x"2f00", 66=>x"3500", 67=>x"3900", 68=>x"3100",
---- 69=>x"3300", 70=>x"3600", 71=>x"3600", 72=>x"cf00",
---- 73=>x"3600", 74=>x"3400", 75=>x"2d00", 76=>x"3200",
---- 77=>x"2f00", 78=>x"2f00", 79=>x"3000", 80=>x"3000",
---- 81=>x"2d00", 82=>x"2c00", 83=>x"2f00", 84=>x"2f00",
---- 85=>x"2d00", 86=>x"2e00", 87=>x"2b00", 88=>x"2b00",
---- 89=>x"2f00", 90=>x"3100", 91=>x"2c00", 92=>x"2c00",
---- 93=>x"2f00", 94=>x"2e00", 95=>x"2e00", 96=>x"3000",
---- 97=>x"2e00", 98=>x"2f00", 99=>x"3100", 100=>x"d200",
---- 101=>x"2e00", 102=>x"2f00", 103=>x"2d00", 104=>x"3000",
---- 105=>x"2a00", 106=>x"2b00", 107=>x"2c00", 108=>x"3000",
---- 109=>x"2f00", 110=>x"2c00", 111=>x"2e00", 112=>x"2d00",
---- 113=>x"2a00", 114=>x"3000", 115=>x"3000", 116=>x"2d00",
---- 117=>x"2d00", 118=>x"2d00", 119=>x"3000", 120=>x"3600",
---- 121=>x"2d00", 122=>x"3000", 123=>x"3300", 124=>x"2f00",
---- 125=>x"2c00", 126=>x"3600", 127=>x"3700", 128=>x"2f00",
---- 129=>x"3600", 130=>x"3600", 131=>x"3200", 132=>x"3600",
---- 133=>x"3700", 134=>x"2d00", 135=>x"2200", 136=>x"3b00",
---- 137=>x"3400", 138=>x"2200", 139=>x"1d00", 140=>x"3c00",
---- 141=>x"2600", 142=>x"1a00", 143=>x"2000", 144=>x"3100",
---- 145=>x"2300", 146=>x"1a00", 147=>x"3e00", 148=>x"2100",
---- 149=>x"1d00", 150=>x"3500", 151=>x"7a00", 152=>x"2200",
---- 153=>x"3100", 154=>x"6a00", 155=>x"9a00", 156=>x"2f00",
---- 157=>x"5900", 158=>x"8c00", 159=>x"a300", 160=>x"5800",
---- 161=>x"8300", 162=>x"9800", 163=>x"a600", 164=>x"8000",
---- 165=>x"9400", 166=>x"9b00", 167=>x"a300", 168=>x"9000",
---- 169=>x"9600", 170=>x"6700", 171=>x"9c00", 172=>x"9700",
---- 173=>x"9300", 174=>x"9200", 175=>x"9700", 176=>x"9800",
---- 177=>x"9100", 178=>x"8e00", 179=>x"8e00", 180=>x"9c00",
---- 181=>x"8f00", 182=>x"8300", 183=>x"9100", 184=>x"9900",
---- 185=>x"8900", 186=>x"8a00", 187=>x"9c00", 188=>x"8f00",
---- 189=>x"8900", 190=>x"9b00", 191=>x"a400", 192=>x"8d00",
---- 193=>x"9800", 194=>x"a000", 195=>x"a300", 196=>x"9b00",
---- 197=>x"a200", 198=>x"a100", 199=>x"a500", 200=>x"a300",
---- 201=>x"a500", 202=>x"a400", 203=>x"a400", 204=>x"a600",
---- 205=>x"a500", 206=>x"a500", 207=>x"a200", 208=>x"a700",
---- 209=>x"a500", 210=>x"a400", 211=>x"a300", 212=>x"a500",
---- 213=>x"a500", 214=>x"a400", 215=>x"a300", 216=>x"a300",
---- 217=>x"a000", 218=>x"a400", 219=>x"a600", 220=>x"a100",
---- 221=>x"a200", 222=>x"a200", 223=>x"5e00", 224=>x"a000",
---- 225=>x"9e00", 226=>x"9f00", 227=>x"9f00", 228=>x"a000",
---- 229=>x"9f00", 230=>x"9e00", 231=>x"9f00", 232=>x"a000",
---- 233=>x"9e00", 234=>x"9e00", 235=>x"9e00", 236=>x"9e00",
---- 237=>x"9d00", 238=>x"9e00", 239=>x"9e00", 240=>x"9f00",
---- 241=>x"9e00", 242=>x"9d00", 243=>x"9d00", 244=>x"9e00",
---- 245=>x"9d00", 246=>x"9d00", 247=>x"9d00", 248=>x"9e00",
---- 249=>x"9e00", 250=>x"9e00", 251=>x"9d00", 252=>x"9d00",
---- 253=>x"9d00", 254=>x"9d00", 255=>x"9f00", 256=>x"9c00",
---- 257=>x"9e00", 258=>x"9d00", 259=>x"a000", 260=>x"9c00",
---- 261=>x"9900", 262=>x"6100", 263=>x"9f00", 264=>x"9c00",
---- 265=>x"9900", 266=>x"9b00", 267=>x"9c00", 268=>x"9c00",
---- 269=>x"9c00", 270=>x"9a00", 271=>x"9a00", 272=>x"9b00",
---- 273=>x"9a00", 274=>x"9a00", 275=>x"9900", 276=>x"9c00",
---- 277=>x"9900", 278=>x"9a00", 279=>x"9a00", 280=>x"9c00",
---- 281=>x"9a00", 282=>x"9a00", 283=>x"9900", 284=>x"9b00",
---- 285=>x"9800", 286=>x"9800", 287=>x"9a00", 288=>x"6300",
---- 289=>x"9a00", 290=>x"9a00", 291=>x"9a00", 292=>x"9b00",
---- 293=>x"9900", 294=>x"9b00", 295=>x"9c00", 296=>x"9d00",
---- 297=>x"9b00", 298=>x"9c00", 299=>x"9b00", 300=>x"9b00",
---- 301=>x"9c00", 302=>x"9d00", 303=>x"9c00", 304=>x"9c00",
---- 305=>x"9d00", 306=>x"a000", 307=>x"9e00", 308=>x"9e00",
---- 309=>x"9d00", 310=>x"9d00", 311=>x"9d00", 312=>x"9d00",
---- 313=>x"9b00", 314=>x"9c00", 315=>x"9d00", 316=>x"9e00",
---- 317=>x"9c00", 318=>x"9e00", 319=>x"9d00", 320=>x"9f00",
---- 321=>x"9b00", 322=>x"9900", 323=>x"9e00", 324=>x"9c00",
---- 325=>x"9c00", 326=>x"9f00", 327=>x"9e00", 328=>x"9c00",
---- 329=>x"9b00", 330=>x"9c00", 331=>x"9c00", 332=>x"9d00",
---- 333=>x"9c00", 334=>x"9d00", 335=>x"9d00", 336=>x"9e00",
---- 337=>x"9b00", 338=>x"9c00", 339=>x"9b00", 340=>x"9b00",
---- 341=>x"9b00", 342=>x"9b00", 343=>x"9a00", 344=>x"9a00",
---- 345=>x"9a00", 346=>x"9a00", 347=>x"9a00", 348=>x"6400",
---- 349=>x"9800", 350=>x"9b00", 351=>x"9a00", 352=>x"9a00",
---- 353=>x"9700", 354=>x"9a00", 355=>x"9900", 356=>x"9b00",
---- 357=>x"9800", 358=>x"9c00", 359=>x"9a00", 360=>x"9b00",
---- 361=>x"9c00", 362=>x"9b00", 363=>x"9900", 364=>x"9700",
---- 365=>x"9900", 366=>x"9a00", 367=>x"9a00", 368=>x"9a00",
---- 369=>x"9700", 370=>x"9700", 371=>x"9900", 372=>x"9900",
---- 373=>x"9b00", 374=>x"9a00", 375=>x"9900", 376=>x"9c00",
---- 377=>x"9900", 378=>x"6500", 379=>x"9800", 380=>x"9b00",
---- 381=>x"9800", 382=>x"9800", 383=>x"9600", 384=>x"9c00",
---- 385=>x"9700", 386=>x"9800", 387=>x"9600", 388=>x"9a00",
---- 389=>x"9800", 390=>x"9800", 391=>x"9700", 392=>x"9b00",
---- 393=>x"9900", 394=>x"9800", 395=>x"9800", 396=>x"9a00",
---- 397=>x"9a00", 398=>x"9a00", 399=>x"9700", 400=>x"9b00",
---- 401=>x"9900", 402=>x"9800", 403=>x"9700", 404=>x"9900",
---- 405=>x"9800", 406=>x"9600", 407=>x"9a00", 408=>x"9a00",
---- 409=>x"9800", 410=>x"9600", 411=>x"9600", 412=>x"9c00",
---- 413=>x"9800", 414=>x"9900", 415=>x"9900", 416=>x"9b00",
---- 417=>x"9900", 418=>x"9900", 419=>x"9800", 420=>x"9800",
---- 421=>x"9800", 422=>x"9600", 423=>x"9700", 424=>x"9b00",
---- 425=>x"9900", 426=>x"9700", 427=>x"9900", 428=>x"9b00",
---- 429=>x"9900", 430=>x"9a00", 431=>x"9800", 432=>x"9b00",
---- 433=>x"9900", 434=>x"9600", 435=>x"9700", 436=>x"9c00",
---- 437=>x"9a00", 438=>x"9900", 439=>x"9600", 440=>x"9c00",
---- 441=>x"9a00", 442=>x"9900", 443=>x"9700", 444=>x"9b00",
---- 445=>x"9800", 446=>x"9900", 447=>x"9700", 448=>x"9b00",
---- 449=>x"9900", 450=>x"9600", 451=>x"9700", 452=>x"9d00",
---- 453=>x"6400", 454=>x"9900", 455=>x"9700", 456=>x"9b00",
---- 457=>x"9900", 458=>x"9900", 459=>x"9600", 460=>x"9700",
---- 461=>x"9400", 462=>x"9700", 463=>x"9400", 464=>x"9900",
---- 465=>x"9900", 466=>x"9800", 467=>x"9600", 468=>x"9a00",
---- 469=>x"9800", 470=>x"9700", 471=>x"9600", 472=>x"9a00",
---- 473=>x"9800", 474=>x"9700", 475=>x"9700", 476=>x"9700",
---- 477=>x"6700", 478=>x"9600", 479=>x"9500", 480=>x"9600",
---- 481=>x"9800", 482=>x"9800", 483=>x"9800", 484=>x"9000",
---- 485=>x"9300", 486=>x"9500", 487=>x"9600", 488=>x"8c00",
---- 489=>x"8d00", 490=>x"8c00", 491=>x"8e00", 492=>x"8b00",
---- 493=>x"8c00", 494=>x"8800", 495=>x"8800", 496=>x"8c00",
---- 497=>x"8a00", 498=>x"8500", 499=>x"8600", 500=>x"8d00",
---- 501=>x"8600", 502=>x"8600", 503=>x"8500", 504=>x"8b00",
---- 505=>x"8700", 506=>x"8500", 507=>x"8400", 508=>x"8900",
---- 509=>x"8700", 510=>x"8700", 511=>x"8400", 512=>x"9000",
---- 513=>x"8b00", 514=>x"8b00", 515=>x"8800", 516=>x"8e00",
---- 517=>x"8e00", 518=>x"8a00", 519=>x"8700", 520=>x"8b00",
---- 521=>x"8b00", 522=>x"8900", 523=>x"8700", 524=>x"8900",
---- 525=>x"8900", 526=>x"8800", 527=>x"8600", 528=>x"8700",
---- 529=>x"8500", 530=>x"8700", 531=>x"8400", 532=>x"8300",
---- 533=>x"7e00", 534=>x"7f00", 535=>x"8300", 536=>x"8000",
---- 537=>x"8500", 538=>x"8b00", 539=>x"9700", 540=>x"8d00",
---- 541=>x"9600", 542=>x"9f00", 543=>x"5700", 544=>x"a100",
---- 545=>x"a600", 546=>x"ac00", 547=>x"b400", 548=>x"b100",
---- 549=>x"b300", 550=>x"b700", 551=>x"bb00", 552=>x"b900",
---- 553=>x"ba00", 554=>x"bb00", 555=>x"be00", 556=>x"bd00",
---- 557=>x"bc00", 558=>x"bb00", 559=>x"bd00", 560=>x"bf00",
---- 561=>x"be00", 562=>x"bc00", 563=>x"bc00", 564=>x"be00",
---- 565=>x"be00", 566=>x"bc00", 567=>x"bd00", 568=>x"bc00",
---- 569=>x"bd00", 570=>x"bd00", 571=>x"be00", 572=>x"bd00",
---- 573=>x"be00", 574=>x"bd00", 575=>x"be00", 576=>x"be00",
---- 577=>x"be00", 578=>x"be00", 579=>x"bf00", 580=>x"bf00",
---- 581=>x"c000", 582=>x"bf00", 583=>x"3d00", 584=>x"c100",
---- 585=>x"c100", 586=>x"c100", 587=>x"c300", 588=>x"c200",
---- 589=>x"c500", 590=>x"c700", 591=>x"c700", 592=>x"c500",
---- 593=>x"c800", 594=>x"c900", 595=>x"ca00", 596=>x"cb00",
---- 597=>x"cb00", 598=>x"cc00", 599=>x"cb00", 600=>x"cc00",
---- 601=>x"ce00", 602=>x"cc00", 603=>x"cc00", 604=>x"cc00",
---- 605=>x"cd00", 606=>x"cc00", 607=>x"cb00", 608=>x"cc00",
---- 609=>x"cb00", 610=>x"cb00", 611=>x"ca00", 612=>x"cd00",
---- 613=>x"ca00", 614=>x"c900", 615=>x"c900", 616=>x"cd00",
---- 617=>x"cc00", 618=>x"ca00", 619=>x"cb00", 620=>x"cd00",
---- 621=>x"cd00", 622=>x"cc00", 623=>x"cd00", 624=>x"cf00",
---- 625=>x"d000", 626=>x"ce00", 627=>x"ce00", 628=>x"d000",
---- 629=>x"d000", 630=>x"ce00", 631=>x"cf00", 632=>x"d100",
---- 633=>x"d000", 634=>x"ce00", 635=>x"cf00", 636=>x"d000",
---- 637=>x"2d00", 638=>x"d100", 639=>x"ce00", 640=>x"d000",
---- 641=>x"d000", 642=>x"d000", 643=>x"cf00", 644=>x"d200",
---- 645=>x"d000", 646=>x"d000", 647=>x"cf00", 648=>x"d200",
---- 649=>x"d200", 650=>x"cf00", 651=>x"cf00", 652=>x"2d00",
---- 653=>x"cf00", 654=>x"ce00", 655=>x"cf00", 656=>x"d000",
---- 657=>x"3000", 658=>x"cf00", 659=>x"d000", 660=>x"d000",
---- 661=>x"cf00", 662=>x"cf00", 663=>x"d200", 664=>x"d100",
---- 665=>x"d200", 666=>x"d200", 667=>x"d300", 668=>x"d200",
---- 669=>x"d300", 670=>x"d300", 671=>x"d300", 672=>x"d200",
---- 673=>x"d500", 674=>x"d400", 675=>x"d400", 676=>x"d200",
---- 677=>x"d300", 678=>x"d200", 679=>x"d400", 680=>x"d200",
---- 681=>x"d300", 682=>x"d200", 683=>x"2c00", 684=>x"d200",
---- 685=>x"d400", 686=>x"d400", 687=>x"d400", 688=>x"d400",
---- 689=>x"d500", 690=>x"d500", 691=>x"d300", 692=>x"d400",
---- 693=>x"d600", 694=>x"d300", 695=>x"d300", 696=>x"d500",
---- 697=>x"d400", 698=>x"d400", 699=>x"d600", 700=>x"d400",
---- 701=>x"d600", 702=>x"d500", 703=>x"d500", 704=>x"d600",
---- 705=>x"d600", 706=>x"d500", 707=>x"d400", 708=>x"d300",
---- 709=>x"d400", 710=>x"d500", 711=>x"d500", 712=>x"d300",
---- 713=>x"d300", 714=>x"d400", 715=>x"d200", 716=>x"d100",
---- 717=>x"d000", 718=>x"cf00", 719=>x"cf00", 720=>x"cf00",
---- 721=>x"cd00", 722=>x"cd00", 723=>x"cd00", 724=>x"cc00",
---- 725=>x"cd00", 726=>x"cc00", 727=>x"cb00", 728=>x"ce00",
---- 729=>x"d100", 730=>x"d000", 731=>x"cf00", 732=>x"d100",
---- 733=>x"d100", 734=>x"d300", 735=>x"d100", 736=>x"d200",
---- 737=>x"d400", 738=>x"2c00", 739=>x"d500", 740=>x"d200",
---- 741=>x"d200", 742=>x"d200", 743=>x"d100", 744=>x"d000",
---- 745=>x"d000", 746=>x"ce00", 747=>x"cf00", 748=>x"cf00",
---- 749=>x"cf00", 750=>x"cf00", 751=>x"cd00", 752=>x"d000",
---- 753=>x"cf00", 754=>x"cd00", 755=>x"cb00", 756=>x"cc00",
---- 757=>x"c900", 758=>x"c800", 759=>x"c300", 760=>x"c300",
---- 761=>x"bc00", 762=>x"b200", 763=>x"9900", 764=>x"9a00",
---- 765=>x"7f00", 766=>x"6200", 767=>x"4400", 768=>x"4600",
---- 769=>x"3300", 770=>x"2d00", 771=>x"2a00", 772=>x"2600",
---- 773=>x"2800", 774=>x"2b00", 775=>x"2d00", 776=>x"2700",
---- 777=>x"2b00", 778=>x"3300", 779=>x"3500", 780=>x"2b00",
---- 781=>x"3500", 782=>x"4400", 783=>x"4500", 784=>x"3d00",
---- 785=>x"4900", 786=>x"5000", 787=>x"4d00", 788=>x"4b00",
---- 789=>x"5500", 790=>x"5200", 791=>x"4c00", 792=>x"5300",
---- 793=>x"5700", 794=>x"5300", 795=>x"5600", 796=>x"5400",
---- 797=>x"5100", 798=>x"5300", 799=>x"5700", 800=>x"5100",
---- 801=>x"5400", 802=>x"5700", 803=>x"5500", 804=>x"a900",
---- 805=>x"5800", 806=>x"5a00", 807=>x"5700", 808=>x"5e00",
---- 809=>x"5400", 810=>x"5300", 811=>x"5500", 812=>x"5b00",
---- 813=>x"5600", 814=>x"5000", 815=>x"5500", 816=>x"5e00",
---- 817=>x"5700", 818=>x"5100", 819=>x"5900", 820=>x"5a00",
---- 821=>x"5b00", 822=>x"5600", 823=>x"6200", 824=>x"5c00",
---- 825=>x"5500", 826=>x"5800", 827=>x"6000", 828=>x"5c00",
---- 829=>x"5700", 830=>x"6100", 831=>x"6500", 832=>x"5b00",
---- 833=>x"5d00", 834=>x"6400", 835=>x"6800", 836=>x"5d00",
---- 837=>x"6500", 838=>x"6600", 839=>x"6600", 840=>x"6200",
---- 841=>x"6600", 842=>x"6b00", 843=>x"6700", 844=>x"6700",
---- 845=>x"6800", 846=>x"6700", 847=>x"6600", 848=>x"6800",
---- 849=>x"6800", 850=>x"6400", 851=>x"6500", 852=>x"6700",
---- 853=>x"6500", 854=>x"6400", 855=>x"6900", 856=>x"6500",
---- 857=>x"5e00", 858=>x"6500", 859=>x"6700", 860=>x"6300",
---- 861=>x"6200", 862=>x"9500", 863=>x"6a00", 864=>x"6500",
---- 865=>x"6200", 866=>x"6700", 867=>x"6500", 868=>x"6600",
---- 869=>x"6500", 870=>x"6800", 871=>x"5f00", 872=>x"6700",
---- 873=>x"6600", 874=>x"6800", 875=>x"5a00", 876=>x"5f00",
---- 877=>x"6200", 878=>x"5800", 879=>x"5600", 880=>x"5f00",
---- 881=>x"5b00", 882=>x"5400", 883=>x"5100", 884=>x"9f00",
---- 885=>x"5700", 886=>x"5700", 887=>x"5100", 888=>x"5d00",
---- 889=>x"5200", 890=>x"5c00", 891=>x"5800", 892=>x"5800",
---- 893=>x"5900", 894=>x"5d00", 895=>x"5b00", 896=>x"5a00",
---- 897=>x"5900", 898=>x"5e00", 899=>x"5f00", 900=>x"5e00",
---- 901=>x"5c00", 902=>x"5c00", 903=>x"6100", 904=>x"5f00",
---- 905=>x"5f00", 906=>x"5f00", 907=>x"6100", 908=>x"5f00",
---- 909=>x"5f00", 910=>x"6100", 911=>x"5800", 912=>x"5f00",
---- 913=>x"6300", 914=>x"5e00", 915=>x"4d00", 916=>x"5c00",
---- 917=>x"6000", 918=>x"5900", 919=>x"4700", 920=>x"5d00",
---- 921=>x"5900", 922=>x"4a00", 923=>x"3d00", 924=>x"5900",
---- 925=>x"5300", 926=>x"4400", 927=>x"3b00", 928=>x"5600",
---- 929=>x"4c00", 930=>x"3c00", 931=>x"3800", 932=>x"4f00",
---- 933=>x"4500", 934=>x"3500", 935=>x"3400", 936=>x"4f00",
---- 937=>x"4200", 938=>x"3800", 939=>x"3400", 940=>x"4500",
---- 941=>x"3a00", 942=>x"3800", 943=>x"3600", 944=>x"3d00",
---- 945=>x"3b00", 946=>x"3300", 947=>x"3200", 948=>x"3d00",
---- 949=>x"3c00", 950=>x"3400", 951=>x"3500", 952=>x"4700",
---- 953=>x"3f00", 954=>x"3600", 955=>x"3a00", 956=>x"4a00",
---- 957=>x"3f00", 958=>x"3b00", 959=>x"3d00", 960=>x"4800",
---- 961=>x"3c00", 962=>x"3a00", 963=>x"4100", 964=>x"4100",
---- 965=>x"3900", 966=>x"4400", 967=>x"4600", 968=>x"3e00",
---- 969=>x"4100", 970=>x"4400", 971=>x"3d00", 972=>x"3d00",
---- 973=>x"4700", 974=>x"4900", 975=>x"3e00", 976=>x"4500",
---- 977=>x"4500", 978=>x"4900", 979=>x"3e00", 980=>x"4900",
---- 981=>x"4200", 982=>x"4100", 983=>x"3900", 984=>x"3f00",
---- 985=>x"4000", 986=>x"3a00", 987=>x"cf00", 988=>x"3c00",
---- 989=>x"3c00", 990=>x"3500", 991=>x"3400", 992=>x"3e00",
---- 993=>x"3900", 994=>x"3600", 995=>x"3700", 996=>x"3500",
---- 997=>x"3400", 998=>x"3300", 999=>x"3000", 1000=>x"3500",
---- 1001=>x"3700", 1002=>x"3200", 1003=>x"3500", 1004=>x"3400",
---- 1005=>x"3700", 1006=>x"3800", 1007=>x"4600", 1008=>x"3900",
---- 1009=>x"3a00", 1010=>x"4700", 1011=>x"5100", 1012=>x"4100",
---- 1013=>x"4b00", 1014=>x"5900", 1015=>x"5b00", 1016=>x"4900",
---- 1017=>x"5700", 1018=>x"6100", 1019=>x"6100", 1020=>x"5700",
---- 1021=>x"6000", 1022=>x"6500", 1023=>x"6800")
---- );
--
end content_package;

package body content_package is
end content_package;
